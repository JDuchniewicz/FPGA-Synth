module triangle_lut(input[8:0] i_phase,
								output reg signed[15:0] o_val);
        initial o_val = 16'b0;

		always @(i_phase) begin
			case(i_phase)
            9'h000 	:	o_val <= 16'b0000000000000000;
            9'h001 	:	o_val <= 16'b0000000001000000;
            9'h002 	:	o_val <= 16'b0000000010000000;
            9'h003 	:	o_val <= 16'b0000000011000000;
            9'h004 	:	o_val <= 16'b0000000100000000;
            9'h005 	:	o_val <= 16'b0000000101000000;
            9'h006 	:	o_val <= 16'b0000000110000000;
            9'h007 	:	o_val <= 16'b0000000111000000;
            9'h008 	:	o_val <= 16'b0000001000000000;
            9'h009 	:	o_val <= 16'b0000001001000000;
            9'h00a 	:	o_val <= 16'b0000001010000000;
            9'h00b 	:	o_val <= 16'b0000001011000000;
            9'h00c 	:	o_val <= 16'b0000001100000000;
            9'h00d 	:	o_val <= 16'b0000001101000000;
            9'h00e 	:	o_val <= 16'b0000001110000000;
            9'h00f 	:	o_val <= 16'b0000001111000000;
            9'h010 	:	o_val <= 16'b0000010000000000;
            9'h011 	:	o_val <= 16'b0000010001000000;
            9'h012 	:	o_val <= 16'b0000010010000000;
            9'h013 	:	o_val <= 16'b0000010011000000;
            9'h014 	:	o_val <= 16'b0000010100000000;
            9'h015 	:	o_val <= 16'b0000010101000000;
            9'h016 	:	o_val <= 16'b0000010110000000;
            9'h017 	:	o_val <= 16'b0000010111000000;
            9'h018 	:	o_val <= 16'b0000011000000000;
            9'h019 	:	o_val <= 16'b0000011001000000;
            9'h01a 	:	o_val <= 16'b0000011010000000;
            9'h01b 	:	o_val <= 16'b0000011011000000;
            9'h01c 	:	o_val <= 16'b0000011100000000;
            9'h01d 	:	o_val <= 16'b0000011101000000;
            9'h01e 	:	o_val <= 16'b0000011110000000;
            9'h01f 	:	o_val <= 16'b0000011111000000;
            9'h020 	:	o_val <= 16'b0000100000000000;
            9'h021 	:	o_val <= 16'b0000100001000000;
            9'h022 	:	o_val <= 16'b0000100010000000;
            9'h023 	:	o_val <= 16'b0000100011000000;
            9'h024 	:	o_val <= 16'b0000100100000000;
            9'h025 	:	o_val <= 16'b0000100101000000;
            9'h026 	:	o_val <= 16'b0000100110000000;
            9'h027 	:	o_val <= 16'b0000100111000000;
            9'h028 	:	o_val <= 16'b0000101000000000;
            9'h029 	:	o_val <= 16'b0000101001000000;
            9'h02a 	:	o_val <= 16'b0000101010000000;
            9'h02b 	:	o_val <= 16'b0000101011000000;
            9'h02c 	:	o_val <= 16'b0000101100000000;
            9'h02d 	:	o_val <= 16'b0000101101000000;
            9'h02e 	:	o_val <= 16'b0000101110000000;
            9'h02f 	:	o_val <= 16'b0000101111000000;
            9'h030 	:	o_val <= 16'b0000110000000000;
            9'h031 	:	o_val <= 16'b0000110001000000;
            9'h032 	:	o_val <= 16'b0000110010000000;
            9'h033 	:	o_val <= 16'b0000110011000000;
            9'h034 	:	o_val <= 16'b0000110100000000;
            9'h035 	:	o_val <= 16'b0000110101000000;
            9'h036 	:	o_val <= 16'b0000110110000000;
            9'h037 	:	o_val <= 16'b0000110111000000;
            9'h038 	:	o_val <= 16'b0000111000000000;
            9'h039 	:	o_val <= 16'b0000111001000000;
            9'h03a 	:	o_val <= 16'b0000111010000000;
            9'h03b 	:	o_val <= 16'b0000111011000000;
            9'h03c 	:	o_val <= 16'b0000111100000000;
            9'h03d 	:	o_val <= 16'b0000111101000000;
            9'h03e 	:	o_val <= 16'b0000111110000000;
            9'h03f 	:	o_val <= 16'b0000111111000000;
            9'h040 	:	o_val <= 16'b0001000000000000;
            9'h041 	:	o_val <= 16'b0001000001000000;
            9'h042 	:	o_val <= 16'b0001000010000000;
            9'h043 	:	o_val <= 16'b0001000011000000;
            9'h044 	:	o_val <= 16'b0001000100000000;
            9'h045 	:	o_val <= 16'b0001000101000000;
            9'h046 	:	o_val <= 16'b0001000110000000;
            9'h047 	:	o_val <= 16'b0001000111000000;
            9'h048 	:	o_val <= 16'b0001001000000000;
            9'h049 	:	o_val <= 16'b0001001001000000;
            9'h04a 	:	o_val <= 16'b0001001010000000;
            9'h04b 	:	o_val <= 16'b0001001011000000;
            9'h04c 	:	o_val <= 16'b0001001100000000;
            9'h04d 	:	o_val <= 16'b0001001101000000;
            9'h04e 	:	o_val <= 16'b0001001110000000;
            9'h04f 	:	o_val <= 16'b0001001111000000;
            9'h050 	:	o_val <= 16'b0001010000000000;
            9'h051 	:	o_val <= 16'b0001010001000000;
            9'h052 	:	o_val <= 16'b0001010010000000;
            9'h053 	:	o_val <= 16'b0001010011000000;
            9'h054 	:	o_val <= 16'b0001010100000000;
            9'h055 	:	o_val <= 16'b0001010101000000;
            9'h056 	:	o_val <= 16'b0001010110000000;
            9'h057 	:	o_val <= 16'b0001010111000000;
            9'h058 	:	o_val <= 16'b0001011000000000;
            9'h059 	:	o_val <= 16'b0001011001000000;
            9'h05a 	:	o_val <= 16'b0001011010000000;
            9'h05b 	:	o_val <= 16'b0001011011000000;
            9'h05c 	:	o_val <= 16'b0001011100000000;
            9'h05d 	:	o_val <= 16'b0001011101000000;
            9'h05e 	:	o_val <= 16'b0001011110000000;
            9'h05f 	:	o_val <= 16'b0001011111000000;
            9'h060 	:	o_val <= 16'b0001100000000000;
            9'h061 	:	o_val <= 16'b0001100001000000;
            9'h062 	:	o_val <= 16'b0001100010000000;
            9'h063 	:	o_val <= 16'b0001100011000000;
            9'h064 	:	o_val <= 16'b0001100100000000;
            9'h065 	:	o_val <= 16'b0001100101000000;
            9'h066 	:	o_val <= 16'b0001100110000000;
            9'h067 	:	o_val <= 16'b0001100111000000;
            9'h068 	:	o_val <= 16'b0001101000000000;
            9'h069 	:	o_val <= 16'b0001101001000000;
            9'h06a 	:	o_val <= 16'b0001101010000000;
            9'h06b 	:	o_val <= 16'b0001101011000000;
            9'h06c 	:	o_val <= 16'b0001101100000000;
            9'h06d 	:	o_val <= 16'b0001101101000000;
            9'h06e 	:	o_val <= 16'b0001101110000000;
            9'h06f 	:	o_val <= 16'b0001101111000000;
            9'h070 	:	o_val <= 16'b0001110000000000;
            9'h071 	:	o_val <= 16'b0001110001000000;
            9'h072 	:	o_val <= 16'b0001110010000000;
            9'h073 	:	o_val <= 16'b0001110011000000;
            9'h074 	:	o_val <= 16'b0001110100000000;
            9'h075 	:	o_val <= 16'b0001110101000000;
            9'h076 	:	o_val <= 16'b0001110110000000;
            9'h077 	:	o_val <= 16'b0001110111000000;
            9'h078 	:	o_val <= 16'b0001111000000000;
            9'h079 	:	o_val <= 16'b0001111001000000;
            9'h07a 	:	o_val <= 16'b0001111010000000;
            9'h07b 	:	o_val <= 16'b0001111011000000;
            9'h07c 	:	o_val <= 16'b0001111100000000;
            9'h07d 	:	o_val <= 16'b0001111101000000;
            9'h07e 	:	o_val <= 16'b0001111110000000;
            9'h07f 	:	o_val <= 16'b0001111111000000;
            9'h080 	:	o_val <= 16'b0010000000000000;
            9'h081 	:	o_val <= 16'b0010000001000000;
            9'h082 	:	o_val <= 16'b0010000010000000;
            9'h083 	:	o_val <= 16'b0010000011000000;
            9'h084 	:	o_val <= 16'b0010000100000000;
            9'h085 	:	o_val <= 16'b0010000101000000;
            9'h086 	:	o_val <= 16'b0010000110000000;
            9'h087 	:	o_val <= 16'b0010000111000000;
            9'h088 	:	o_val <= 16'b0010001000000000;
            9'h089 	:	o_val <= 16'b0010001001000000;
            9'h08a 	:	o_val <= 16'b0010001010000000;
            9'h08b 	:	o_val <= 16'b0010001011000000;
            9'h08c 	:	o_val <= 16'b0010001100000000;
            9'h08d 	:	o_val <= 16'b0010001101000000;
            9'h08e 	:	o_val <= 16'b0010001110000000;
            9'h08f 	:	o_val <= 16'b0010001111000000;
            9'h090 	:	o_val <= 16'b0010010000000000;
            9'h091 	:	o_val <= 16'b0010010001000000;
            9'h092 	:	o_val <= 16'b0010010010000000;
            9'h093 	:	o_val <= 16'b0010010011000000;
            9'h094 	:	o_val <= 16'b0010010100000000;
            9'h095 	:	o_val <= 16'b0010010101000000;
            9'h096 	:	o_val <= 16'b0010010110000000;
            9'h097 	:	o_val <= 16'b0010010111000000;
            9'h098 	:	o_val <= 16'b0010011000000000;
            9'h099 	:	o_val <= 16'b0010011001000000;
            9'h09a 	:	o_val <= 16'b0010011010000000;
            9'h09b 	:	o_val <= 16'b0010011011000000;
            9'h09c 	:	o_val <= 16'b0010011100000000;
            9'h09d 	:	o_val <= 16'b0010011101000000;
            9'h09e 	:	o_val <= 16'b0010011110000000;
            9'h09f 	:	o_val <= 16'b0010011111000000;
            9'h0a0 	:	o_val <= 16'b0010100000000000;
            9'h0a1 	:	o_val <= 16'b0010100001000000;
            9'h0a2 	:	o_val <= 16'b0010100010000000;
            9'h0a3 	:	o_val <= 16'b0010100011000000;
            9'h0a4 	:	o_val <= 16'b0010100100000000;
            9'h0a5 	:	o_val <= 16'b0010100101000000;
            9'h0a6 	:	o_val <= 16'b0010100110000000;
            9'h0a7 	:	o_val <= 16'b0010100111000000;
            9'h0a8 	:	o_val <= 16'b0010101000000000;
            9'h0a9 	:	o_val <= 16'b0010101001000000;
            9'h0aa 	:	o_val <= 16'b0010101010000000;
            9'h0ab 	:	o_val <= 16'b0010101011000000;
            9'h0ac 	:	o_val <= 16'b0010101100000000;
            9'h0ad 	:	o_val <= 16'b0010101101000000;
            9'h0ae 	:	o_val <= 16'b0010101110000000;
            9'h0af 	:	o_val <= 16'b0010101111000000;
            9'h0b0 	:	o_val <= 16'b0010110000000000;
            9'h0b1 	:	o_val <= 16'b0010110001000000;
            9'h0b2 	:	o_val <= 16'b0010110010000000;
            9'h0b3 	:	o_val <= 16'b0010110011000000;
            9'h0b4 	:	o_val <= 16'b0010110100000000;
            9'h0b5 	:	o_val <= 16'b0010110101000000;
            9'h0b6 	:	o_val <= 16'b0010110110000000;
            9'h0b7 	:	o_val <= 16'b0010110111000000;
            9'h0b8 	:	o_val <= 16'b0010111000000000;
            9'h0b9 	:	o_val <= 16'b0010111001000000;
            9'h0ba 	:	o_val <= 16'b0010111010000000;
            9'h0bb 	:	o_val <= 16'b0010111011000000;
            9'h0bc 	:	o_val <= 16'b0010111100000000;
            9'h0bd 	:	o_val <= 16'b0010111101000000;
            9'h0be 	:	o_val <= 16'b0010111110000000;
            9'h0bf 	:	o_val <= 16'b0010111111000000;
            9'h0c0 	:	o_val <= 16'b0011000000000000;
            9'h0c1 	:	o_val <= 16'b0011000001000000;
            9'h0c2 	:	o_val <= 16'b0011000010000000;
            9'h0c3 	:	o_val <= 16'b0011000011000000;
            9'h0c4 	:	o_val <= 16'b0011000100000000;
            9'h0c5 	:	o_val <= 16'b0011000101000000;
            9'h0c6 	:	o_val <= 16'b0011000110000000;
            9'h0c7 	:	o_val <= 16'b0011000111000000;
            9'h0c8 	:	o_val <= 16'b0011001000000000;
            9'h0c9 	:	o_val <= 16'b0011001001000000;
            9'h0ca 	:	o_val <= 16'b0011001010000000;
            9'h0cb 	:	o_val <= 16'b0011001011000000;
            9'h0cc 	:	o_val <= 16'b0011001100000000;
            9'h0cd 	:	o_val <= 16'b0011001101000000;
            9'h0ce 	:	o_val <= 16'b0011001110000000;
            9'h0cf 	:	o_val <= 16'b0011001111000000;
            9'h0d0 	:	o_val <= 16'b0011010000000000;
            9'h0d1 	:	o_val <= 16'b0011010001000000;
            9'h0d2 	:	o_val <= 16'b0011010010000000;
            9'h0d3 	:	o_val <= 16'b0011010011000000;
            9'h0d4 	:	o_val <= 16'b0011010100000000;
            9'h0d5 	:	o_val <= 16'b0011010101000000;
            9'h0d6 	:	o_val <= 16'b0011010110000000;
            9'h0d7 	:	o_val <= 16'b0011010111000000;
            9'h0d8 	:	o_val <= 16'b0011011000000000;
            9'h0d9 	:	o_val <= 16'b0011011001000000;
            9'h0da 	:	o_val <= 16'b0011011010000000;
            9'h0db 	:	o_val <= 16'b0011011011000000;
            9'h0dc 	:	o_val <= 16'b0011011100000000;
            9'h0dd 	:	o_val <= 16'b0011011101000000;
            9'h0de 	:	o_val <= 16'b0011011110000000;
            9'h0df 	:	o_val <= 16'b0011011111000000;
            9'h0e0 	:	o_val <= 16'b0011100000000000;
            9'h0e1 	:	o_val <= 16'b0011100001000000;
            9'h0e2 	:	o_val <= 16'b0011100010000000;
            9'h0e3 	:	o_val <= 16'b0011100011000000;
            9'h0e4 	:	o_val <= 16'b0011100100000000;
            9'h0e5 	:	o_val <= 16'b0011100101000000;
            9'h0e6 	:	o_val <= 16'b0011100110000000;
            9'h0e7 	:	o_val <= 16'b0011100111000000;
            9'h0e8 	:	o_val <= 16'b0011101000000000;
            9'h0e9 	:	o_val <= 16'b0011101001000000;
            9'h0ea 	:	o_val <= 16'b0011101010000000;
            9'h0eb 	:	o_val <= 16'b0011101011000000;
            9'h0ec 	:	o_val <= 16'b0011101100000000;
            9'h0ed 	:	o_val <= 16'b0011101101000000;
            9'h0ee 	:	o_val <= 16'b0011101110000000;
            9'h0ef 	:	o_val <= 16'b0011101111000000;
            9'h0f0 	:	o_val <= 16'b0011110000000000;
            9'h0f1 	:	o_val <= 16'b0011110001000000;
            9'h0f2 	:	o_val <= 16'b0011110010000000;
            9'h0f3 	:	o_val <= 16'b0011110011000000;
            9'h0f4 	:	o_val <= 16'b0011110100000000;
            9'h0f5 	:	o_val <= 16'b0011110101000000;
            9'h0f6 	:	o_val <= 16'b0011110110000000;
            9'h0f7 	:	o_val <= 16'b0011110111000000;
            9'h0f8 	:	o_val <= 16'b0011111000000000;
            9'h0f9 	:	o_val <= 16'b0011111001000000;
            9'h0fa 	:	o_val <= 16'b0011111010000000;
            9'h0fb 	:	o_val <= 16'b0011111011000000;
            9'h0fc 	:	o_val <= 16'b0011111100000000;
            9'h0fd 	:	o_val <= 16'b0011111101000000;
            9'h0fe 	:	o_val <= 16'b0011111110000000;
            9'h0ff 	:	o_val <= 16'b0011111111000000;
            9'h100 	:	o_val <= 16'b0100000000000000;
            9'h101 	:	o_val <= 16'b0100000001000000;
            9'h102 	:	o_val <= 16'b0100000010000000;
            9'h103 	:	o_val <= 16'b0100000011000000;
            9'h104 	:	o_val <= 16'b0100000100000000;
            9'h105 	:	o_val <= 16'b0100000101000000;
            9'h106 	:	o_val <= 16'b0100000110000000;
            9'h107 	:	o_val <= 16'b0100000111000000;
            9'h108 	:	o_val <= 16'b0100001000000000;
            9'h109 	:	o_val <= 16'b0100001001000000;
            9'h10a 	:	o_val <= 16'b0100001010000000;
            9'h10b 	:	o_val <= 16'b0100001011000000;
            9'h10c 	:	o_val <= 16'b0100001100000000;
            9'h10d 	:	o_val <= 16'b0100001101000000;
            9'h10e 	:	o_val <= 16'b0100001110000000;
            9'h10f 	:	o_val <= 16'b0100001111000000;
            9'h110 	:	o_val <= 16'b0100010000000000;
            9'h111 	:	o_val <= 16'b0100010001000000;
            9'h112 	:	o_val <= 16'b0100010010000000;
            9'h113 	:	o_val <= 16'b0100010011000000;
            9'h114 	:	o_val <= 16'b0100010100000000;
            9'h115 	:	o_val <= 16'b0100010101000000;
            9'h116 	:	o_val <= 16'b0100010110000000;
            9'h117 	:	o_val <= 16'b0100010111000000;
            9'h118 	:	o_val <= 16'b0100011000000000;
            9'h119 	:	o_val <= 16'b0100011001000000;
            9'h11a 	:	o_val <= 16'b0100011010000000;
            9'h11b 	:	o_val <= 16'b0100011011000000;
            9'h11c 	:	o_val <= 16'b0100011100000000;
            9'h11d 	:	o_val <= 16'b0100011101000000;
            9'h11e 	:	o_val <= 16'b0100011110000000;
            9'h11f 	:	o_val <= 16'b0100011111000000;
            9'h120 	:	o_val <= 16'b0100100000000000;
            9'h121 	:	o_val <= 16'b0100100001000000;
            9'h122 	:	o_val <= 16'b0100100010000000;
            9'h123 	:	o_val <= 16'b0100100011000000;
            9'h124 	:	o_val <= 16'b0100100100000000;
            9'h125 	:	o_val <= 16'b0100100101000000;
            9'h126 	:	o_val <= 16'b0100100110000000;
            9'h127 	:	o_val <= 16'b0100100111000000;
            9'h128 	:	o_val <= 16'b0100101000000000;
            9'h129 	:	o_val <= 16'b0100101001000000;
            9'h12a 	:	o_val <= 16'b0100101010000000;
            9'h12b 	:	o_val <= 16'b0100101011000000;
            9'h12c 	:	o_val <= 16'b0100101100000000;
            9'h12d 	:	o_val <= 16'b0100101101000000;
            9'h12e 	:	o_val <= 16'b0100101110000000;
            9'h12f 	:	o_val <= 16'b0100101111000000;
            9'h130 	:	o_val <= 16'b0100110000000000;
            9'h131 	:	o_val <= 16'b0100110001000000;
            9'h132 	:	o_val <= 16'b0100110010000000;
            9'h133 	:	o_val <= 16'b0100110011000000;
            9'h134 	:	o_val <= 16'b0100110100000000;
            9'h135 	:	o_val <= 16'b0100110101000000;
            9'h136 	:	o_val <= 16'b0100110110000000;
            9'h137 	:	o_val <= 16'b0100110111000000;
            9'h138 	:	o_val <= 16'b0100111000000000;
            9'h139 	:	o_val <= 16'b0100111001000000;
            9'h13a 	:	o_val <= 16'b0100111010000000;
            9'h13b 	:	o_val <= 16'b0100111011000000;
            9'h13c 	:	o_val <= 16'b0100111100000000;
            9'h13d 	:	o_val <= 16'b0100111101000000;
            9'h13e 	:	o_val <= 16'b0100111110000000;
            9'h13f 	:	o_val <= 16'b0100111111000000;
            9'h140 	:	o_val <= 16'b0101000000000000;
            9'h141 	:	o_val <= 16'b0101000001000000;
            9'h142 	:	o_val <= 16'b0101000010000000;
            9'h143 	:	o_val <= 16'b0101000011000000;
            9'h144 	:	o_val <= 16'b0101000100000000;
            9'h145 	:	o_val <= 16'b0101000101000000;
            9'h146 	:	o_val <= 16'b0101000110000000;
            9'h147 	:	o_val <= 16'b0101000111000000;
            9'h148 	:	o_val <= 16'b0101001000000000;
            9'h149 	:	o_val <= 16'b0101001001000000;
            9'h14a 	:	o_val <= 16'b0101001010000000;
            9'h14b 	:	o_val <= 16'b0101001011000000;
            9'h14c 	:	o_val <= 16'b0101001100000000;
            9'h14d 	:	o_val <= 16'b0101001101000000;
            9'h14e 	:	o_val <= 16'b0101001110000000;
            9'h14f 	:	o_val <= 16'b0101001111000000;
            9'h150 	:	o_val <= 16'b0101010000000000;
            9'h151 	:	o_val <= 16'b0101010001000000;
            9'h152 	:	o_val <= 16'b0101010010000000;
            9'h153 	:	o_val <= 16'b0101010011000000;
            9'h154 	:	o_val <= 16'b0101010100000000;
            9'h155 	:	o_val <= 16'b0101010101000000;
            9'h156 	:	o_val <= 16'b0101010110000000;
            9'h157 	:	o_val <= 16'b0101010111000000;
            9'h158 	:	o_val <= 16'b0101011000000000;
            9'h159 	:	o_val <= 16'b0101011001000000;
            9'h15a 	:	o_val <= 16'b0101011010000000;
            9'h15b 	:	o_val <= 16'b0101011011000000;
            9'h15c 	:	o_val <= 16'b0101011100000000;
            9'h15d 	:	o_val <= 16'b0101011101000000;
            9'h15e 	:	o_val <= 16'b0101011110000000;
            9'h15f 	:	o_val <= 16'b0101011111000000;
            9'h160 	:	o_val <= 16'b0101100000000000;
            9'h161 	:	o_val <= 16'b0101100001000000;
            9'h162 	:	o_val <= 16'b0101100010000000;
            9'h163 	:	o_val <= 16'b0101100011000000;
            9'h164 	:	o_val <= 16'b0101100100000000;
            9'h165 	:	o_val <= 16'b0101100101000000;
            9'h166 	:	o_val <= 16'b0101100110000000;
            9'h167 	:	o_val <= 16'b0101100111000000;
            9'h168 	:	o_val <= 16'b0101101000000000;
            9'h169 	:	o_val <= 16'b0101101001000000;
            9'h16a 	:	o_val <= 16'b0101101010000000;
            9'h16b 	:	o_val <= 16'b0101101011000000;
            9'h16c 	:	o_val <= 16'b0101101100000000;
            9'h16d 	:	o_val <= 16'b0101101101000000;
            9'h16e 	:	o_val <= 16'b0101101110000000;
            9'h16f 	:	o_val <= 16'b0101101111000000;
            9'h170 	:	o_val <= 16'b0101110000000000;
            9'h171 	:	o_val <= 16'b0101110001000000;
            9'h172 	:	o_val <= 16'b0101110010000000;
            9'h173 	:	o_val <= 16'b0101110011000000;
            9'h174 	:	o_val <= 16'b0101110100000000;
            9'h175 	:	o_val <= 16'b0101110101000000;
            9'h176 	:	o_val <= 16'b0101110110000000;
            9'h177 	:	o_val <= 16'b0101110111000000;
            9'h178 	:	o_val <= 16'b0101111000000000;
            9'h179 	:	o_val <= 16'b0101111001000000;
            9'h17a 	:	o_val <= 16'b0101111010000000;
            9'h17b 	:	o_val <= 16'b0101111011000000;
            9'h17c 	:	o_val <= 16'b0101111100000000;
            9'h17d 	:	o_val <= 16'b0101111101000000;
            9'h17e 	:	o_val <= 16'b0101111110000000;
            9'h17f 	:	o_val <= 16'b0101111111000000;
            9'h180 	:	o_val <= 16'b0110000000000000;
            9'h181 	:	o_val <= 16'b0110000001000000;
            9'h182 	:	o_val <= 16'b0110000010000000;
            9'h183 	:	o_val <= 16'b0110000011000000;
            9'h184 	:	o_val <= 16'b0110000100000000;
            9'h185 	:	o_val <= 16'b0110000101000000;
            9'h186 	:	o_val <= 16'b0110000110000000;
            9'h187 	:	o_val <= 16'b0110000111000000;
            9'h188 	:	o_val <= 16'b0110001000000000;
            9'h189 	:	o_val <= 16'b0110001001000000;
            9'h18a 	:	o_val <= 16'b0110001010000000;
            9'h18b 	:	o_val <= 16'b0110001011000000;
            9'h18c 	:	o_val <= 16'b0110001100000000;
            9'h18d 	:	o_val <= 16'b0110001101000000;
            9'h18e 	:	o_val <= 16'b0110001110000000;
            9'h18f 	:	o_val <= 16'b0110001111000000;
            9'h190 	:	o_val <= 16'b0110010000000000;
            9'h191 	:	o_val <= 16'b0110010001000000;
            9'h192 	:	o_val <= 16'b0110010010000000;
            9'h193 	:	o_val <= 16'b0110010011000000;
            9'h194 	:	o_val <= 16'b0110010100000000;
            9'h195 	:	o_val <= 16'b0110010101000000;
            9'h196 	:	o_val <= 16'b0110010110000000;
            9'h197 	:	o_val <= 16'b0110010111000000;
            9'h198 	:	o_val <= 16'b0110011000000000;
            9'h199 	:	o_val <= 16'b0110011001000000;
            9'h19a 	:	o_val <= 16'b0110011010000000;
            9'h19b 	:	o_val <= 16'b0110011011000000;
            9'h19c 	:	o_val <= 16'b0110011100000000;
            9'h19d 	:	o_val <= 16'b0110011101000000;
            9'h19e 	:	o_val <= 16'b0110011110000000;
            9'h19f 	:	o_val <= 16'b0110011111000000;
            9'h1a0 	:	o_val <= 16'b0110100000000000;
            9'h1a1 	:	o_val <= 16'b0110100001000000;
            9'h1a2 	:	o_val <= 16'b0110100010000000;
            9'h1a3 	:	o_val <= 16'b0110100011000000;
            9'h1a4 	:	o_val <= 16'b0110100100000000;
            9'h1a5 	:	o_val <= 16'b0110100101000000;
            9'h1a6 	:	o_val <= 16'b0110100110000000;
            9'h1a7 	:	o_val <= 16'b0110100111000000;
            9'h1a8 	:	o_val <= 16'b0110101000000000;
            9'h1a9 	:	o_val <= 16'b0110101001000000;
            9'h1aa 	:	o_val <= 16'b0110101010000000;
            9'h1ab 	:	o_val <= 16'b0110101011000000;
            9'h1ac 	:	o_val <= 16'b0110101100000000;
            9'h1ad 	:	o_val <= 16'b0110101101000000;
            9'h1ae 	:	o_val <= 16'b0110101110000000;
            9'h1af 	:	o_val <= 16'b0110101111000000;
            9'h1b0 	:	o_val <= 16'b0110110000000000;
            9'h1b1 	:	o_val <= 16'b0110110001000000;
            9'h1b2 	:	o_val <= 16'b0110110010000000;
            9'h1b3 	:	o_val <= 16'b0110110011000000;
            9'h1b4 	:	o_val <= 16'b0110110100000000;
            9'h1b5 	:	o_val <= 16'b0110110101000000;
            9'h1b6 	:	o_val <= 16'b0110110110000000;
            9'h1b7 	:	o_val <= 16'b0110110111000000;
            9'h1b8 	:	o_val <= 16'b0110111000000000;
            9'h1b9 	:	o_val <= 16'b0110111001000000;
            9'h1ba 	:	o_val <= 16'b0110111010000000;
            9'h1bb 	:	o_val <= 16'b0110111011000000;
            9'h1bc 	:	o_val <= 16'b0110111100000000;
            9'h1bd 	:	o_val <= 16'b0110111101000000;
            9'h1be 	:	o_val <= 16'b0110111110000000;
            9'h1bf 	:	o_val <= 16'b0110111111000000;
            9'h1c0 	:	o_val <= 16'b0111000000000000;
            9'h1c1 	:	o_val <= 16'b0111000001000000;
            9'h1c2 	:	o_val <= 16'b0111000010000000;
            9'h1c3 	:	o_val <= 16'b0111000011000000;
            9'h1c4 	:	o_val <= 16'b0111000100000000;
            9'h1c5 	:	o_val <= 16'b0111000101000000;
            9'h1c6 	:	o_val <= 16'b0111000110000000;
            9'h1c7 	:	o_val <= 16'b0111000111000000;
            9'h1c8 	:	o_val <= 16'b0111001000000000;
            9'h1c9 	:	o_val <= 16'b0111001001000000;
            9'h1ca 	:	o_val <= 16'b0111001010000000;
            9'h1cb 	:	o_val <= 16'b0111001011000000;
            9'h1cc 	:	o_val <= 16'b0111001100000000;
            9'h1cd 	:	o_val <= 16'b0111001101000000;
            9'h1ce 	:	o_val <= 16'b0111001110000000;
            9'h1cf 	:	o_val <= 16'b0111001111000000;
            9'h1d0 	:	o_val <= 16'b0111010000000000;
            9'h1d1 	:	o_val <= 16'b0111010001000000;
            9'h1d2 	:	o_val <= 16'b0111010010000000;
            9'h1d3 	:	o_val <= 16'b0111010011000000;
            9'h1d4 	:	o_val <= 16'b0111010100000000;
            9'h1d5 	:	o_val <= 16'b0111010101000000;
            9'h1d6 	:	o_val <= 16'b0111010110000000;
            9'h1d7 	:	o_val <= 16'b0111010111000000;
            9'h1d8 	:	o_val <= 16'b0111011000000000;
            9'h1d9 	:	o_val <= 16'b0111011001000000;
            9'h1da 	:	o_val <= 16'b0111011010000000;
            9'h1db 	:	o_val <= 16'b0111011011000000;
            9'h1dc 	:	o_val <= 16'b0111011100000000;
            9'h1dd 	:	o_val <= 16'b0111011101000000;
            9'h1de 	:	o_val <= 16'b0111011110000000;
            9'h1df 	:	o_val <= 16'b0111011111000000;
            9'h1e0 	:	o_val <= 16'b0111100000000000;
            9'h1e1 	:	o_val <= 16'b0111100001000000;
            9'h1e2 	:	o_val <= 16'b0111100010000000;
            9'h1e3 	:	o_val <= 16'b0111100011000000;
            9'h1e4 	:	o_val <= 16'b0111100100000000;
            9'h1e5 	:	o_val <= 16'b0111100101000000;
            9'h1e6 	:	o_val <= 16'b0111100110000000;
            9'h1e7 	:	o_val <= 16'b0111100111000000;
            9'h1e8 	:	o_val <= 16'b0111101000000000;
            9'h1e9 	:	o_val <= 16'b0111101001000000;
            9'h1ea 	:	o_val <= 16'b0111101010000000;
            9'h1eb 	:	o_val <= 16'b0111101011000000;
            9'h1ec 	:	o_val <= 16'b0111101100000000;
            9'h1ed 	:	o_val <= 16'b0111101101000000;
            9'h1ee 	:	o_val <= 16'b0111101110000000;
            9'h1ef 	:	o_val <= 16'b0111101111000000;
            9'h1f0 	:	o_val <= 16'b0111110000000000;
            9'h1f1 	:	o_val <= 16'b0111110001000000;
            9'h1f2 	:	o_val <= 16'b0111110010000000;
            9'h1f3 	:	o_val <= 16'b0111110011000000;
            9'h1f4 	:	o_val <= 16'b0111110100000000;
            9'h1f5 	:	o_val <= 16'b0111110101000000;
            9'h1f6 	:	o_val <= 16'b0111110110000000;
            9'h1f7 	:	o_val <= 16'b0111110111000000;
            9'h1f8 	:	o_val <= 16'b0111111000000000;
            9'h1f9 	:	o_val <= 16'b0111111001000000;
            9'h1fa 	:	o_val <= 16'b0111111010000000;
            9'h1fb 	:	o_val <= 16'b0111111011000000;
            9'h1fc 	:	o_val <= 16'b0111111100000000;
            9'h1fd 	:	o_val <= 16'b0111111101000000;
            9'h1fe 	:	o_val <= 16'b0111111110000000;
            9'h1ff 	:	o_val <= 16'b0111111111000000;
				default		:	o_val <= 16'b0;
			endcase
		end
endmodule
