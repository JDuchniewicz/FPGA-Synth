// modules for LUT's for multiple sinewaves for SIMPLE synthesis


//TODO: clock enable has to be given because it cannot be always enabled
// for now just A4 (440kHz) generating module (for phase calculation) 
module dummyA4(clk, val_out); // maybe different style of coding, everything in module declaration?
	input clk;
	output reg [15:0] val_out;
	reg [31:0] phase;
	// Phase increment can be precalculated = 188978561.024 (ignoring the truncated part) -> 2^32 * fd /fs
	
	wire [15:0] lut_out;
	assign lut_out = val_out;
	
	// for now wire it like this? can it be done simpler?
	sineLUT lut(.clk(clk), .index(phase[31:16]), .val_out(lut_out));
	
	always @(posedge clk)
		phase <= phase + 32'h0b43_9581;
	
endmodule

// for now let's assume 8192 samples = 2^13, generate four quarters of one cycle for now (simplify later, but requires more logic)
module sineLUT(clk, index, val_out);
	input clk;
	input [15:0] index; // has to be bus?
	output reg [15:0] val_out; //width?
	
	always @(posedge clk) begin
		case (index)
			4'h000 	:	val_out <= 4'h8000;
         4'h001 	:	val_out <= 4'h8000;
         4'h002 	:	val_out <= 4'h8000;
         4'h003 	:	val_out <= 4'h8000;
         4'h008 	:	val_out <= 4'h8019;
         4'h009 	:	val_out <= 4'h8019;
         4'h00a 	:	val_out <= 4'h8019;
         4'h00b 	:	val_out <= 4'h8019;
         4'h010 	:	val_out <= 4'h8032;
         4'h011 	:	val_out <= 4'h8032;
         4'h012 	:	val_out <= 4'h8032;
         4'h013 	:	val_out <= 4'h8032;
         4'h018 	:	val_out <= 4'h804b;
         4'h019 	:	val_out <= 4'h804b;
         4'h01a 	:	val_out <= 4'h804b;
         4'h01b 	:	val_out <= 4'h804b;
         4'h020 	:	val_out <= 4'h8064;
         4'h021 	:	val_out <= 4'h8064;
         4'h022 	:	val_out <= 4'h8064;
         4'h023 	:	val_out <= 4'h8064;
         4'h028 	:	val_out <= 4'h807d;
         4'h029 	:	val_out <= 4'h807d;
         4'h02a 	:	val_out <= 4'h807d;
         4'h02b 	:	val_out <= 4'h807d;
         4'h030 	:	val_out <= 4'h8096;
         4'h031 	:	val_out <= 4'h8096;
         4'h032 	:	val_out <= 4'h8096;
         4'h033 	:	val_out <= 4'h8096;
         4'h038 	:	val_out <= 4'h80af;
         4'h039 	:	val_out <= 4'h80af;
         4'h03a 	:	val_out <= 4'h80af;
         4'h03b 	:	val_out <= 4'h80af;
         4'h040 	:	val_out <= 4'h80c9;
         4'h041 	:	val_out <= 4'h80c9;
         4'h042 	:	val_out <= 4'h80c9;
         4'h043 	:	val_out <= 4'h80c9;
         4'h048 	:	val_out <= 4'h80e2;
         4'h049 	:	val_out <= 4'h80e2;
         4'h04a 	:	val_out <= 4'h80e2;
         4'h04b 	:	val_out <= 4'h80e2;
         4'h050 	:	val_out <= 4'h80fb;
         4'h051 	:	val_out <= 4'h80fb;
         4'h052 	:	val_out <= 4'h80fb;
         4'h053 	:	val_out <= 4'h80fb;
         4'h058 	:	val_out <= 4'h8114;
         4'h059 	:	val_out <= 4'h8114;
         4'h05a 	:	val_out <= 4'h8114;
         4'h05b 	:	val_out <= 4'h8114;
         4'h060 	:	val_out <= 4'h812d;
         4'h061 	:	val_out <= 4'h812d;
         4'h062 	:	val_out <= 4'h812d;
         4'h063 	:	val_out <= 4'h812d;
         4'h068 	:	val_out <= 4'h8146;
         4'h069 	:	val_out <= 4'h8146;
         4'h06a 	:	val_out <= 4'h8146;
         4'h06b 	:	val_out <= 4'h8146;
         4'h070 	:	val_out <= 4'h815f;
         4'h071 	:	val_out <= 4'h815f;
         4'h072 	:	val_out <= 4'h815f;
         4'h073 	:	val_out <= 4'h815f;
         4'h078 	:	val_out <= 4'h8178;
         4'h079 	:	val_out <= 4'h8178;
         4'h07a 	:	val_out <= 4'h8178;
         4'h07b 	:	val_out <= 4'h8178;
         4'h080 	:	val_out <= 4'h8192;
         4'h081 	:	val_out <= 4'h8192;
         4'h082 	:	val_out <= 4'h8192;
         4'h083 	:	val_out <= 4'h8192;
         4'h088 	:	val_out <= 4'h81ab;
         4'h089 	:	val_out <= 4'h81ab;
         4'h08a 	:	val_out <= 4'h81ab;
         4'h08b 	:	val_out <= 4'h81ab;
         4'h090 	:	val_out <= 4'h81c4;
         4'h091 	:	val_out <= 4'h81c4;
         4'h092 	:	val_out <= 4'h81c4;
         4'h093 	:	val_out <= 4'h81c4;
         4'h098 	:	val_out <= 4'h81dd;
         4'h099 	:	val_out <= 4'h81dd;
         4'h09a 	:	val_out <= 4'h81dd;
         4'h09b 	:	val_out <= 4'h81dd;
         4'h0a0 	:	val_out <= 4'h81f6;
         4'h0a1 	:	val_out <= 4'h81f6;
         4'h0a2 	:	val_out <= 4'h81f6;
         4'h0a3 	:	val_out <= 4'h81f6;
         4'h0a8 	:	val_out <= 4'h820f;
         4'h0a9 	:	val_out <= 4'h820f;
         4'h0aa 	:	val_out <= 4'h820f;
         4'h0ab 	:	val_out <= 4'h820f;
         4'h0b0 	:	val_out <= 4'h8228;
         4'h0b1 	:	val_out <= 4'h8228;
         4'h0b2 	:	val_out <= 4'h8228;
         4'h0b3 	:	val_out <= 4'h8228;
         4'h0b8 	:	val_out <= 4'h8242;
         4'h0b9 	:	val_out <= 4'h8242;
         4'h0ba 	:	val_out <= 4'h8242;
         4'h0bb 	:	val_out <= 4'h8242;
         4'h0c0 	:	val_out <= 4'h825b;
         4'h0c1 	:	val_out <= 4'h825b;
         4'h0c2 	:	val_out <= 4'h825b;
         4'h0c3 	:	val_out <= 4'h825b;
         4'h0c8 	:	val_out <= 4'h8274;
         4'h0c9 	:	val_out <= 4'h8274;
         4'h0ca 	:	val_out <= 4'h8274;
         4'h0cb 	:	val_out <= 4'h8274;
         4'h0d0 	:	val_out <= 4'h828d;
         4'h0d1 	:	val_out <= 4'h828d;
         4'h0d2 	:	val_out <= 4'h828d;
         4'h0d3 	:	val_out <= 4'h828d;
         4'h0d8 	:	val_out <= 4'h82a6;
         4'h0d9 	:	val_out <= 4'h82a6;
         4'h0da 	:	val_out <= 4'h82a6;
         4'h0db 	:	val_out <= 4'h82a6;
         4'h0e0 	:	val_out <= 4'h82bf;
         4'h0e1 	:	val_out <= 4'h82bf;
         4'h0e2 	:	val_out <= 4'h82bf;
         4'h0e3 	:	val_out <= 4'h82bf;
         4'h0e8 	:	val_out <= 4'h82d8;
         4'h0e9 	:	val_out <= 4'h82d8;
         4'h0ea 	:	val_out <= 4'h82d8;
         4'h0eb 	:	val_out <= 4'h82d8;
         4'h0f0 	:	val_out <= 4'h82f1;
         4'h0f1 	:	val_out <= 4'h82f1;
         4'h0f2 	:	val_out <= 4'h82f1;
         4'h0f3 	:	val_out <= 4'h82f1;
         4'h0f8 	:	val_out <= 4'h830b;
         4'h0f9 	:	val_out <= 4'h830b;
         4'h0fa 	:	val_out <= 4'h830b;
         4'h0fb 	:	val_out <= 4'h830b;
         4'h100 	:	val_out <= 4'h8324;
         4'h101 	:	val_out <= 4'h8324;
         4'h102 	:	val_out <= 4'h8324;
         4'h103 	:	val_out <= 4'h8324;
         4'h108 	:	val_out <= 4'h833d;
         4'h109 	:	val_out <= 4'h833d;
         4'h10a 	:	val_out <= 4'h833d;
         4'h10b 	:	val_out <= 4'h833d;
         4'h110 	:	val_out <= 4'h8356;
         4'h111 	:	val_out <= 4'h8356;
         4'h112 	:	val_out <= 4'h8356;
         4'h113 	:	val_out <= 4'h8356;
         4'h118 	:	val_out <= 4'h836f;
         4'h119 	:	val_out <= 4'h836f;
         4'h11a 	:	val_out <= 4'h836f;
         4'h11b 	:	val_out <= 4'h836f;
         4'h120 	:	val_out <= 4'h8388;
         4'h121 	:	val_out <= 4'h8388;
         4'h122 	:	val_out <= 4'h8388;
         4'h123 	:	val_out <= 4'h8388;
         4'h128 	:	val_out <= 4'h83a1;
         4'h129 	:	val_out <= 4'h83a1;
         4'h12a 	:	val_out <= 4'h83a1;
         4'h12b 	:	val_out <= 4'h83a1;
         4'h130 	:	val_out <= 4'h83ba;
         4'h131 	:	val_out <= 4'h83ba;
         4'h132 	:	val_out <= 4'h83ba;
         4'h133 	:	val_out <= 4'h83ba;
         4'h138 	:	val_out <= 4'h83d4;
         4'h139 	:	val_out <= 4'h83d4;
         4'h13a 	:	val_out <= 4'h83d4;
         4'h13b 	:	val_out <= 4'h83d4;
         4'h140 	:	val_out <= 4'h83ed;
         4'h141 	:	val_out <= 4'h83ed;
         4'h142 	:	val_out <= 4'h83ed;
         4'h143 	:	val_out <= 4'h83ed;
         4'h148 	:	val_out <= 4'h8406;
         4'h149 	:	val_out <= 4'h8406;
         4'h14a 	:	val_out <= 4'h8406;
         4'h14b 	:	val_out <= 4'h8406;
         4'h150 	:	val_out <= 4'h841f;
         4'h151 	:	val_out <= 4'h841f;
         4'h152 	:	val_out <= 4'h841f;
         4'h153 	:	val_out <= 4'h841f;
         4'h158 	:	val_out <= 4'h8438;
         4'h159 	:	val_out <= 4'h8438;
         4'h15a 	:	val_out <= 4'h8438;
         4'h15b 	:	val_out <= 4'h8438;
         4'h160 	:	val_out <= 4'h8451;
         4'h161 	:	val_out <= 4'h8451;
         4'h162 	:	val_out <= 4'h8451;
         4'h163 	:	val_out <= 4'h8451;
         4'h168 	:	val_out <= 4'h846a;
         4'h169 	:	val_out <= 4'h846a;
         4'h16a 	:	val_out <= 4'h846a;
         4'h16b 	:	val_out <= 4'h846a;
         4'h170 	:	val_out <= 4'h8483;
         4'h171 	:	val_out <= 4'h8483;
         4'h172 	:	val_out <= 4'h8483;
         4'h173 	:	val_out <= 4'h8483;
         4'h178 	:	val_out <= 4'h849c;
         4'h179 	:	val_out <= 4'h849c;
         4'h17a 	:	val_out <= 4'h849c;
         4'h17b 	:	val_out <= 4'h849c;
         4'h180 	:	val_out <= 4'h84b6;
         4'h181 	:	val_out <= 4'h84b6;
         4'h182 	:	val_out <= 4'h84b6;
         4'h183 	:	val_out <= 4'h84b6;
         4'h188 	:	val_out <= 4'h84cf;
         4'h189 	:	val_out <= 4'h84cf;
         4'h18a 	:	val_out <= 4'h84cf;
         4'h18b 	:	val_out <= 4'h84cf;
         4'h190 	:	val_out <= 4'h84e8;
         4'h191 	:	val_out <= 4'h84e8;
         4'h192 	:	val_out <= 4'h84e8;
         4'h193 	:	val_out <= 4'h84e8;
         4'h198 	:	val_out <= 4'h8501;
         4'h199 	:	val_out <= 4'h8501;
         4'h19a 	:	val_out <= 4'h8501;
         4'h19b 	:	val_out <= 4'h8501;
         4'h1a0 	:	val_out <= 4'h851a;
         4'h1a1 	:	val_out <= 4'h851a;
         4'h1a2 	:	val_out <= 4'h851a;
         4'h1a3 	:	val_out <= 4'h851a;
         4'h1a8 	:	val_out <= 4'h8533;
         4'h1a9 	:	val_out <= 4'h8533;
         4'h1aa 	:	val_out <= 4'h8533;
         4'h1ab 	:	val_out <= 4'h8533;
         4'h1b0 	:	val_out <= 4'h854c;
         4'h1b1 	:	val_out <= 4'h854c;
         4'h1b2 	:	val_out <= 4'h854c;
         4'h1b3 	:	val_out <= 4'h854c;
         4'h1b8 	:	val_out <= 4'h8565;
         4'h1b9 	:	val_out <= 4'h8565;
         4'h1ba 	:	val_out <= 4'h8565;
         4'h1bb 	:	val_out <= 4'h8565;
         4'h1c0 	:	val_out <= 4'h857f;
         4'h1c1 	:	val_out <= 4'h857f;
         4'h1c2 	:	val_out <= 4'h857f;
         4'h1c3 	:	val_out <= 4'h857f;
         4'h1c8 	:	val_out <= 4'h8598;
         4'h1c9 	:	val_out <= 4'h8598;
         4'h1ca 	:	val_out <= 4'h8598;
         4'h1cb 	:	val_out <= 4'h8598;
         4'h1d0 	:	val_out <= 4'h85b1;
         4'h1d1 	:	val_out <= 4'h85b1;
         4'h1d2 	:	val_out <= 4'h85b1;
         4'h1d3 	:	val_out <= 4'h85b1;
         4'h1d8 	:	val_out <= 4'h85ca;
         4'h1d9 	:	val_out <= 4'h85ca;
         4'h1da 	:	val_out <= 4'h85ca;
         4'h1db 	:	val_out <= 4'h85ca;
         4'h1e0 	:	val_out <= 4'h85e3;
         4'h1e1 	:	val_out <= 4'h85e3;
         4'h1e2 	:	val_out <= 4'h85e3;
         4'h1e3 	:	val_out <= 4'h85e3;
         4'h1e8 	:	val_out <= 4'h85fc;
         4'h1e9 	:	val_out <= 4'h85fc;
         4'h1ea 	:	val_out <= 4'h85fc;
         4'h1eb 	:	val_out <= 4'h85fc;
         4'h1f0 	:	val_out <= 4'h8615;
         4'h1f1 	:	val_out <= 4'h8615;
         4'h1f2 	:	val_out <= 4'h8615;
         4'h1f3 	:	val_out <= 4'h8615;
         4'h1f8 	:	val_out <= 4'h862e;
         4'h1f9 	:	val_out <= 4'h862e;
         4'h1fa 	:	val_out <= 4'h862e;
         4'h1fb 	:	val_out <= 4'h862e;
         4'h200 	:	val_out <= 4'h8647;
         4'h201 	:	val_out <= 4'h8647;
         4'h202 	:	val_out <= 4'h8647;
         4'h203 	:	val_out <= 4'h8647;
         4'h208 	:	val_out <= 4'h8660;
         4'h209 	:	val_out <= 4'h8660;
         4'h20a 	:	val_out <= 4'h8660;
         4'h20b 	:	val_out <= 4'h8660;
         4'h210 	:	val_out <= 4'h867a;
         4'h211 	:	val_out <= 4'h867a;
         4'h212 	:	val_out <= 4'h867a;
         4'h213 	:	val_out <= 4'h867a;
         4'h218 	:	val_out <= 4'h8693;
         4'h219 	:	val_out <= 4'h8693;
         4'h21a 	:	val_out <= 4'h8693;
         4'h21b 	:	val_out <= 4'h8693;
         4'h220 	:	val_out <= 4'h86ac;
         4'h221 	:	val_out <= 4'h86ac;
         4'h222 	:	val_out <= 4'h86ac;
         4'h223 	:	val_out <= 4'h86ac;
         4'h228 	:	val_out <= 4'h86c5;
         4'h229 	:	val_out <= 4'h86c5;
         4'h22a 	:	val_out <= 4'h86c5;
         4'h22b 	:	val_out <= 4'h86c5;
         4'h230 	:	val_out <= 4'h86de;
         4'h231 	:	val_out <= 4'h86de;
         4'h232 	:	val_out <= 4'h86de;
         4'h233 	:	val_out <= 4'h86de;
         4'h238 	:	val_out <= 4'h86f7;
         4'h239 	:	val_out <= 4'h86f7;
         4'h23a 	:	val_out <= 4'h86f7;
         4'h23b 	:	val_out <= 4'h86f7;
         4'h240 	:	val_out <= 4'h8710;
         4'h241 	:	val_out <= 4'h8710;
         4'h242 	:	val_out <= 4'h8710;
         4'h243 	:	val_out <= 4'h8710;
         4'h248 	:	val_out <= 4'h8729;
         4'h249 	:	val_out <= 4'h8729;
         4'h24a 	:	val_out <= 4'h8729;
         4'h24b 	:	val_out <= 4'h8729;
         4'h250 	:	val_out <= 4'h8742;
         4'h251 	:	val_out <= 4'h8742;
         4'h252 	:	val_out <= 4'h8742;
         4'h253 	:	val_out <= 4'h8742;
         4'h258 	:	val_out <= 4'h875b;
         4'h259 	:	val_out <= 4'h875b;
         4'h25a 	:	val_out <= 4'h875b;
         4'h25b 	:	val_out <= 4'h875b;
         4'h260 	:	val_out <= 4'h8775;
         4'h261 	:	val_out <= 4'h8775;
         4'h262 	:	val_out <= 4'h8775;
         4'h263 	:	val_out <= 4'h8775;
         4'h268 	:	val_out <= 4'h878e;
         4'h269 	:	val_out <= 4'h878e;
         4'h26a 	:	val_out <= 4'h878e;
         4'h26b 	:	val_out <= 4'h878e;
         4'h270 	:	val_out <= 4'h87a7;
         4'h271 	:	val_out <= 4'h87a7;
         4'h272 	:	val_out <= 4'h87a7;
         4'h273 	:	val_out <= 4'h87a7;
         4'h278 	:	val_out <= 4'h87c0;
         4'h279 	:	val_out <= 4'h87c0;
         4'h27a 	:	val_out <= 4'h87c0;
         4'h27b 	:	val_out <= 4'h87c0;
         4'h280 	:	val_out <= 4'h87d9;
         4'h281 	:	val_out <= 4'h87d9;
         4'h282 	:	val_out <= 4'h87d9;
         4'h283 	:	val_out <= 4'h87d9;
         4'h288 	:	val_out <= 4'h87f2;
         4'h289 	:	val_out <= 4'h87f2;
         4'h28a 	:	val_out <= 4'h87f2;
         4'h28b 	:	val_out <= 4'h87f2;
         4'h290 	:	val_out <= 4'h880b;
         4'h291 	:	val_out <= 4'h880b;
         4'h292 	:	val_out <= 4'h880b;
         4'h293 	:	val_out <= 4'h880b;
         4'h298 	:	val_out <= 4'h8824;
         4'h299 	:	val_out <= 4'h8824;
         4'h29a 	:	val_out <= 4'h8824;
         4'h29b 	:	val_out <= 4'h8824;
         4'h2a0 	:	val_out <= 4'h883d;
         4'h2a1 	:	val_out <= 4'h883d;
         4'h2a2 	:	val_out <= 4'h883d;
         4'h2a3 	:	val_out <= 4'h883d;
         4'h2a8 	:	val_out <= 4'h8856;
         4'h2a9 	:	val_out <= 4'h8856;
         4'h2aa 	:	val_out <= 4'h8856;
         4'h2ab 	:	val_out <= 4'h8856;
         4'h2b0 	:	val_out <= 4'h886f;
         4'h2b1 	:	val_out <= 4'h886f;
         4'h2b2 	:	val_out <= 4'h886f;
         4'h2b3 	:	val_out <= 4'h886f;
         4'h2b8 	:	val_out <= 4'h8888;
         4'h2b9 	:	val_out <= 4'h8888;
         4'h2ba 	:	val_out <= 4'h8888;
         4'h2bb 	:	val_out <= 4'h8888;
         4'h2c0 	:	val_out <= 4'h88a2;
         4'h2c1 	:	val_out <= 4'h88a2;
         4'h2c2 	:	val_out <= 4'h88a2;
         4'h2c3 	:	val_out <= 4'h88a2;
         4'h2c8 	:	val_out <= 4'h88bb;
         4'h2c9 	:	val_out <= 4'h88bb;
         4'h2ca 	:	val_out <= 4'h88bb;
         4'h2cb 	:	val_out <= 4'h88bb;
         4'h2d0 	:	val_out <= 4'h88d4;
         4'h2d1 	:	val_out <= 4'h88d4;
         4'h2d2 	:	val_out <= 4'h88d4;
         4'h2d3 	:	val_out <= 4'h88d4;
         4'h2d8 	:	val_out <= 4'h88ed;
         4'h2d9 	:	val_out <= 4'h88ed;
         4'h2da 	:	val_out <= 4'h88ed;
         4'h2db 	:	val_out <= 4'h88ed;
         4'h2e0 	:	val_out <= 4'h8906;
         4'h2e1 	:	val_out <= 4'h8906;
         4'h2e2 	:	val_out <= 4'h8906;
         4'h2e3 	:	val_out <= 4'h8906;
         4'h2e8 	:	val_out <= 4'h891f;
         4'h2e9 	:	val_out <= 4'h891f;
         4'h2ea 	:	val_out <= 4'h891f;
         4'h2eb 	:	val_out <= 4'h891f;
         4'h2f0 	:	val_out <= 4'h8938;
         4'h2f1 	:	val_out <= 4'h8938;
         4'h2f2 	:	val_out <= 4'h8938;
         4'h2f3 	:	val_out <= 4'h8938;
         4'h2f8 	:	val_out <= 4'h8951;
         4'h2f9 	:	val_out <= 4'h8951;
         4'h2fa 	:	val_out <= 4'h8951;
         4'h2fb 	:	val_out <= 4'h8951;
         4'h300 	:	val_out <= 4'h896a;
         4'h301 	:	val_out <= 4'h896a;
         4'h302 	:	val_out <= 4'h896a;
         4'h303 	:	val_out <= 4'h896a;
         4'h308 	:	val_out <= 4'h8983;
         4'h309 	:	val_out <= 4'h8983;
         4'h30a 	:	val_out <= 4'h8983;
         4'h30b 	:	val_out <= 4'h8983;
         4'h310 	:	val_out <= 4'h899c;
         4'h311 	:	val_out <= 4'h899c;
         4'h312 	:	val_out <= 4'h899c;
         4'h313 	:	val_out <= 4'h899c;
         4'h318 	:	val_out <= 4'h89b5;
         4'h319 	:	val_out <= 4'h89b5;
         4'h31a 	:	val_out <= 4'h89b5;
         4'h31b 	:	val_out <= 4'h89b5;
         4'h320 	:	val_out <= 4'h89ce;
         4'h321 	:	val_out <= 4'h89ce;
         4'h322 	:	val_out <= 4'h89ce;
         4'h323 	:	val_out <= 4'h89ce;
         4'h328 	:	val_out <= 4'h89e7;
         4'h329 	:	val_out <= 4'h89e7;
         4'h32a 	:	val_out <= 4'h89e7;
         4'h32b 	:	val_out <= 4'h89e7;
         4'h330 	:	val_out <= 4'h8a00;
         4'h331 	:	val_out <= 4'h8a00;
         4'h332 	:	val_out <= 4'h8a00;
         4'h333 	:	val_out <= 4'h8a00;
         4'h338 	:	val_out <= 4'h8a19;
         4'h339 	:	val_out <= 4'h8a19;
         4'h33a 	:	val_out <= 4'h8a19;
         4'h33b 	:	val_out <= 4'h8a19;
         4'h340 	:	val_out <= 4'h8a33;
         4'h341 	:	val_out <= 4'h8a33;
         4'h342 	:	val_out <= 4'h8a33;
         4'h343 	:	val_out <= 4'h8a33;
         4'h348 	:	val_out <= 4'h8a4c;
         4'h349 	:	val_out <= 4'h8a4c;
         4'h34a 	:	val_out <= 4'h8a4c;
         4'h34b 	:	val_out <= 4'h8a4c;
         4'h350 	:	val_out <= 4'h8a65;
         4'h351 	:	val_out <= 4'h8a65;
         4'h352 	:	val_out <= 4'h8a65;
         4'h353 	:	val_out <= 4'h8a65;
         4'h358 	:	val_out <= 4'h8a7e;
         4'h359 	:	val_out <= 4'h8a7e;
         4'h35a 	:	val_out <= 4'h8a7e;
         4'h35b 	:	val_out <= 4'h8a7e;
         4'h360 	:	val_out <= 4'h8a97;
         4'h361 	:	val_out <= 4'h8a97;
         4'h362 	:	val_out <= 4'h8a97;
         4'h363 	:	val_out <= 4'h8a97;
         4'h368 	:	val_out <= 4'h8ab0;
         4'h369 	:	val_out <= 4'h8ab0;
         4'h36a 	:	val_out <= 4'h8ab0;
         4'h36b 	:	val_out <= 4'h8ab0;
         4'h370 	:	val_out <= 4'h8ac9;
         4'h371 	:	val_out <= 4'h8ac9;
         4'h372 	:	val_out <= 4'h8ac9;
         4'h373 	:	val_out <= 4'h8ac9;
         4'h378 	:	val_out <= 4'h8ae2;
         4'h379 	:	val_out <= 4'h8ae2;
         4'h37a 	:	val_out <= 4'h8ae2;
         4'h37b 	:	val_out <= 4'h8ae2;
         4'h380 	:	val_out <= 4'h8afb;
         4'h381 	:	val_out <= 4'h8afb;
         4'h382 	:	val_out <= 4'h8afb;
         4'h383 	:	val_out <= 4'h8afb;
         4'h388 	:	val_out <= 4'h8b14;
         4'h389 	:	val_out <= 4'h8b14;
         4'h38a 	:	val_out <= 4'h8b14;
         4'h38b 	:	val_out <= 4'h8b14;
         4'h390 	:	val_out <= 4'h8b2d;
         4'h391 	:	val_out <= 4'h8b2d;
         4'h392 	:	val_out <= 4'h8b2d;
         4'h393 	:	val_out <= 4'h8b2d;
         4'h398 	:	val_out <= 4'h8b46;
         4'h399 	:	val_out <= 4'h8b46;
         4'h39a 	:	val_out <= 4'h8b46;
         4'h39b 	:	val_out <= 4'h8b46;
         4'h3a0 	:	val_out <= 4'h8b5f;
         4'h3a1 	:	val_out <= 4'h8b5f;
         4'h3a2 	:	val_out <= 4'h8b5f;
         4'h3a3 	:	val_out <= 4'h8b5f;
         4'h3a8 	:	val_out <= 4'h8b78;
         4'h3a9 	:	val_out <= 4'h8b78;
         4'h3aa 	:	val_out <= 4'h8b78;
         4'h3ab 	:	val_out <= 4'h8b78;
         4'h3b0 	:	val_out <= 4'h8b91;
         4'h3b1 	:	val_out <= 4'h8b91;
         4'h3b2 	:	val_out <= 4'h8b91;
         4'h3b3 	:	val_out <= 4'h8b91;
         4'h3b8 	:	val_out <= 4'h8baa;
         4'h3b9 	:	val_out <= 4'h8baa;
         4'h3ba 	:	val_out <= 4'h8baa;
         4'h3bb 	:	val_out <= 4'h8baa;
         4'h3c0 	:	val_out <= 4'h8bc3;
         4'h3c1 	:	val_out <= 4'h8bc3;
         4'h3c2 	:	val_out <= 4'h8bc3;
         4'h3c3 	:	val_out <= 4'h8bc3;
         4'h3c8 	:	val_out <= 4'h8bdc;
         4'h3c9 	:	val_out <= 4'h8bdc;
         4'h3ca 	:	val_out <= 4'h8bdc;
         4'h3cb 	:	val_out <= 4'h8bdc;
         4'h3d0 	:	val_out <= 4'h8bf5;
         4'h3d1 	:	val_out <= 4'h8bf5;
         4'h3d2 	:	val_out <= 4'h8bf5;
         4'h3d3 	:	val_out <= 4'h8bf5;
         4'h3d8 	:	val_out <= 4'h8c0e;
         4'h3d9 	:	val_out <= 4'h8c0e;
         4'h3da 	:	val_out <= 4'h8c0e;
         4'h3db 	:	val_out <= 4'h8c0e;
         4'h3e0 	:	val_out <= 4'h8c27;
         4'h3e1 	:	val_out <= 4'h8c27;
         4'h3e2 	:	val_out <= 4'h8c27;
         4'h3e3 	:	val_out <= 4'h8c27;
         4'h3e8 	:	val_out <= 4'h8c40;
         4'h3e9 	:	val_out <= 4'h8c40;
         4'h3ea 	:	val_out <= 4'h8c40;
         4'h3eb 	:	val_out <= 4'h8c40;
         4'h3f0 	:	val_out <= 4'h8c59;
         4'h3f1 	:	val_out <= 4'h8c59;
         4'h3f2 	:	val_out <= 4'h8c59;
         4'h3f3 	:	val_out <= 4'h8c59;
         4'h3f8 	:	val_out <= 4'h8c72;
         4'h3f9 	:	val_out <= 4'h8c72;
         4'h3fa 	:	val_out <= 4'h8c72;
         4'h3fb 	:	val_out <= 4'h8c72;
         4'h400 	:	val_out <= 4'h8c8b;
         4'h401 	:	val_out <= 4'h8c8b;
         4'h402 	:	val_out <= 4'h8c8b;
         4'h403 	:	val_out <= 4'h8c8b;
         4'h408 	:	val_out <= 4'h8ca4;
         4'h409 	:	val_out <= 4'h8ca4;
         4'h40a 	:	val_out <= 4'h8ca4;
         4'h40b 	:	val_out <= 4'h8ca4;
         4'h410 	:	val_out <= 4'h8cbd;
         4'h411 	:	val_out <= 4'h8cbd;
         4'h412 	:	val_out <= 4'h8cbd;
         4'h413 	:	val_out <= 4'h8cbd;
         4'h418 	:	val_out <= 4'h8cd6;
         4'h419 	:	val_out <= 4'h8cd6;
         4'h41a 	:	val_out <= 4'h8cd6;
         4'h41b 	:	val_out <= 4'h8cd6;
         4'h420 	:	val_out <= 4'h8cef;
         4'h421 	:	val_out <= 4'h8cef;
         4'h422 	:	val_out <= 4'h8cef;
         4'h423 	:	val_out <= 4'h8cef;
         4'h428 	:	val_out <= 4'h8d08;
         4'h429 	:	val_out <= 4'h8d08;
         4'h42a 	:	val_out <= 4'h8d08;
         4'h42b 	:	val_out <= 4'h8d08;
         4'h430 	:	val_out <= 4'h8d21;
         4'h431 	:	val_out <= 4'h8d21;
         4'h432 	:	val_out <= 4'h8d21;
         4'h433 	:	val_out <= 4'h8d21;
         4'h438 	:	val_out <= 4'h8d3a;
         4'h439 	:	val_out <= 4'h8d3a;
         4'h43a 	:	val_out <= 4'h8d3a;
         4'h43b 	:	val_out <= 4'h8d3a;
         4'h440 	:	val_out <= 4'h8d53;
         4'h441 	:	val_out <= 4'h8d53;
         4'h442 	:	val_out <= 4'h8d53;
         4'h443 	:	val_out <= 4'h8d53;
         4'h448 	:	val_out <= 4'h8d6c;
         4'h449 	:	val_out <= 4'h8d6c;
         4'h44a 	:	val_out <= 4'h8d6c;
         4'h44b 	:	val_out <= 4'h8d6c;
         4'h450 	:	val_out <= 4'h8d85;
         4'h451 	:	val_out <= 4'h8d85;
         4'h452 	:	val_out <= 4'h8d85;
         4'h453 	:	val_out <= 4'h8d85;
         4'h458 	:	val_out <= 4'h8d9e;
         4'h459 	:	val_out <= 4'h8d9e;
         4'h45a 	:	val_out <= 4'h8d9e;
         4'h45b 	:	val_out <= 4'h8d9e;
         4'h460 	:	val_out <= 4'h8db7;
         4'h461 	:	val_out <= 4'h8db7;
         4'h462 	:	val_out <= 4'h8db7;
         4'h463 	:	val_out <= 4'h8db7;
         4'h468 	:	val_out <= 4'h8dd0;
         4'h469 	:	val_out <= 4'h8dd0;
         4'h46a 	:	val_out <= 4'h8dd0;
         4'h46b 	:	val_out <= 4'h8dd0;
         4'h470 	:	val_out <= 4'h8de9;
         4'h471 	:	val_out <= 4'h8de9;
         4'h472 	:	val_out <= 4'h8de9;
         4'h473 	:	val_out <= 4'h8de9;
         4'h478 	:	val_out <= 4'h8e02;
         4'h479 	:	val_out <= 4'h8e02;
         4'h47a 	:	val_out <= 4'h8e02;
         4'h47b 	:	val_out <= 4'h8e02;
         4'h480 	:	val_out <= 4'h8e1b;
         4'h481 	:	val_out <= 4'h8e1b;
         4'h482 	:	val_out <= 4'h8e1b;
         4'h483 	:	val_out <= 4'h8e1b;
         4'h488 	:	val_out <= 4'h8e34;
         4'h489 	:	val_out <= 4'h8e34;
         4'h48a 	:	val_out <= 4'h8e34;
         4'h48b 	:	val_out <= 4'h8e34;
         4'h490 	:	val_out <= 4'h8e4d;
         4'h491 	:	val_out <= 4'h8e4d;
         4'h492 	:	val_out <= 4'h8e4d;
         4'h493 	:	val_out <= 4'h8e4d;
         4'h498 	:	val_out <= 4'h8e66;
         4'h499 	:	val_out <= 4'h8e66;
         4'h49a 	:	val_out <= 4'h8e66;
         4'h49b 	:	val_out <= 4'h8e66;
         4'h4a0 	:	val_out <= 4'h8e7f;
         4'h4a1 	:	val_out <= 4'h8e7f;
         4'h4a2 	:	val_out <= 4'h8e7f;
         4'h4a3 	:	val_out <= 4'h8e7f;
         4'h4a8 	:	val_out <= 4'h8e98;
         4'h4a9 	:	val_out <= 4'h8e98;
         4'h4aa 	:	val_out <= 4'h8e98;
         4'h4ab 	:	val_out <= 4'h8e98;
         4'h4b0 	:	val_out <= 4'h8eb1;
         4'h4b1 	:	val_out <= 4'h8eb1;
         4'h4b2 	:	val_out <= 4'h8eb1;
         4'h4b3 	:	val_out <= 4'h8eb1;
         4'h4b8 	:	val_out <= 4'h8eca;
         4'h4b9 	:	val_out <= 4'h8eca;
         4'h4ba 	:	val_out <= 4'h8eca;
         4'h4bb 	:	val_out <= 4'h8eca;
         4'h4c0 	:	val_out <= 4'h8ee3;
         4'h4c1 	:	val_out <= 4'h8ee3;
         4'h4c2 	:	val_out <= 4'h8ee3;
         4'h4c3 	:	val_out <= 4'h8ee3;
         4'h4c8 	:	val_out <= 4'h8efc;
         4'h4c9 	:	val_out <= 4'h8efc;
         4'h4ca 	:	val_out <= 4'h8efc;
         4'h4cb 	:	val_out <= 4'h8efc;
         4'h4d0 	:	val_out <= 4'h8f15;
         4'h4d1 	:	val_out <= 4'h8f15;
         4'h4d2 	:	val_out <= 4'h8f15;
         4'h4d3 	:	val_out <= 4'h8f15;
         4'h4d8 	:	val_out <= 4'h8f2e;
         4'h4d9 	:	val_out <= 4'h8f2e;
         4'h4da 	:	val_out <= 4'h8f2e;
         4'h4db 	:	val_out <= 4'h8f2e;
         4'h4e0 	:	val_out <= 4'h8f47;
         4'h4e1 	:	val_out <= 4'h8f47;
         4'h4e2 	:	val_out <= 4'h8f47;
         4'h4e3 	:	val_out <= 4'h8f47;
         4'h4e8 	:	val_out <= 4'h8f60;
         4'h4e9 	:	val_out <= 4'h8f60;
         4'h4ea 	:	val_out <= 4'h8f60;
         4'h4eb 	:	val_out <= 4'h8f60;
         4'h4f0 	:	val_out <= 4'h8f79;
         4'h4f1 	:	val_out <= 4'h8f79;
         4'h4f2 	:	val_out <= 4'h8f79;
         4'h4f3 	:	val_out <= 4'h8f79;
         4'h4f8 	:	val_out <= 4'h8f92;
         4'h4f9 	:	val_out <= 4'h8f92;
         4'h4fa 	:	val_out <= 4'h8f92;
         4'h4fb 	:	val_out <= 4'h8f92;
         4'h500 	:	val_out <= 4'h8fab;
         4'h501 	:	val_out <= 4'h8fab;
         4'h502 	:	val_out <= 4'h8fab;
         4'h503 	:	val_out <= 4'h8fab;
         4'h508 	:	val_out <= 4'h8fc4;
         4'h509 	:	val_out <= 4'h8fc4;
         4'h50a 	:	val_out <= 4'h8fc4;
         4'h50b 	:	val_out <= 4'h8fc4;
         4'h510 	:	val_out <= 4'h8fdd;
         4'h511 	:	val_out <= 4'h8fdd;
         4'h512 	:	val_out <= 4'h8fdd;
         4'h513 	:	val_out <= 4'h8fdd;
         4'h518 	:	val_out <= 4'h8ff5;
         4'h519 	:	val_out <= 4'h8ff5;
         4'h51a 	:	val_out <= 4'h8ff5;
         4'h51b 	:	val_out <= 4'h8ff5;
         4'h520 	:	val_out <= 4'h900e;
         4'h521 	:	val_out <= 4'h900e;
         4'h522 	:	val_out <= 4'h900e;
         4'h523 	:	val_out <= 4'h900e;
         4'h528 	:	val_out <= 4'h9027;
         4'h529 	:	val_out <= 4'h9027;
         4'h52a 	:	val_out <= 4'h9027;
         4'h52b 	:	val_out <= 4'h9027;
         4'h530 	:	val_out <= 4'h9040;
         4'h531 	:	val_out <= 4'h9040;
         4'h532 	:	val_out <= 4'h9040;
         4'h533 	:	val_out <= 4'h9040;
         4'h538 	:	val_out <= 4'h9059;
         4'h539 	:	val_out <= 4'h9059;
         4'h53a 	:	val_out <= 4'h9059;
         4'h53b 	:	val_out <= 4'h9059;
         4'h540 	:	val_out <= 4'h9072;
         4'h541 	:	val_out <= 4'h9072;
         4'h542 	:	val_out <= 4'h9072;
         4'h543 	:	val_out <= 4'h9072;
         4'h548 	:	val_out <= 4'h908b;
         4'h549 	:	val_out <= 4'h908b;
         4'h54a 	:	val_out <= 4'h908b;
         4'h54b 	:	val_out <= 4'h908b;
         4'h550 	:	val_out <= 4'h90a4;
         4'h551 	:	val_out <= 4'h90a4;
         4'h552 	:	val_out <= 4'h90a4;
         4'h553 	:	val_out <= 4'h90a4;
         4'h558 	:	val_out <= 4'h90bd;
         4'h559 	:	val_out <= 4'h90bd;
         4'h55a 	:	val_out <= 4'h90bd;
         4'h55b 	:	val_out <= 4'h90bd;
         4'h560 	:	val_out <= 4'h90d6;
         4'h561 	:	val_out <= 4'h90d6;
         4'h562 	:	val_out <= 4'h90d6;
         4'h563 	:	val_out <= 4'h90d6;
         4'h568 	:	val_out <= 4'h90ef;
         4'h569 	:	val_out <= 4'h90ef;
         4'h56a 	:	val_out <= 4'h90ef;
         4'h56b 	:	val_out <= 4'h90ef;
         4'h570 	:	val_out <= 4'h9108;
         4'h571 	:	val_out <= 4'h9108;
         4'h572 	:	val_out <= 4'h9108;
         4'h573 	:	val_out <= 4'h9108;
         4'h578 	:	val_out <= 4'h9121;
         4'h579 	:	val_out <= 4'h9121;
         4'h57a 	:	val_out <= 4'h9121;
         4'h57b 	:	val_out <= 4'h9121;
         4'h580 	:	val_out <= 4'h9139;
         4'h581 	:	val_out <= 4'h9139;
         4'h582 	:	val_out <= 4'h9139;
         4'h583 	:	val_out <= 4'h9139;
         4'h588 	:	val_out <= 4'h9152;
         4'h589 	:	val_out <= 4'h9152;
         4'h58a 	:	val_out <= 4'h9152;
         4'h58b 	:	val_out <= 4'h9152;
         4'h590 	:	val_out <= 4'h916b;
         4'h591 	:	val_out <= 4'h916b;
         4'h592 	:	val_out <= 4'h916b;
         4'h593 	:	val_out <= 4'h916b;
         4'h598 	:	val_out <= 4'h9184;
         4'h599 	:	val_out <= 4'h9184;
         4'h59a 	:	val_out <= 4'h9184;
         4'h59b 	:	val_out <= 4'h9184;
         4'h5a0 	:	val_out <= 4'h919d;
         4'h5a1 	:	val_out <= 4'h919d;
         4'h5a2 	:	val_out <= 4'h919d;
         4'h5a3 	:	val_out <= 4'h919d;
         4'h5a8 	:	val_out <= 4'h91b6;
         4'h5a9 	:	val_out <= 4'h91b6;
         4'h5aa 	:	val_out <= 4'h91b6;
         4'h5ab 	:	val_out <= 4'h91b6;
         4'h5b0 	:	val_out <= 4'h91cf;
         4'h5b1 	:	val_out <= 4'h91cf;
         4'h5b2 	:	val_out <= 4'h91cf;
         4'h5b3 	:	val_out <= 4'h91cf;
         4'h5b8 	:	val_out <= 4'h91e8;
         4'h5b9 	:	val_out <= 4'h91e8;
         4'h5ba 	:	val_out <= 4'h91e8;
         4'h5bb 	:	val_out <= 4'h91e8;
         4'h5c0 	:	val_out <= 4'h9201;
         4'h5c1 	:	val_out <= 4'h9201;
         4'h5c2 	:	val_out <= 4'h9201;
         4'h5c3 	:	val_out <= 4'h9201;
         4'h5c8 	:	val_out <= 4'h9219;
         4'h5c9 	:	val_out <= 4'h9219;
         4'h5ca 	:	val_out <= 4'h9219;
         4'h5cb 	:	val_out <= 4'h9219;
         4'h5d0 	:	val_out <= 4'h9232;
         4'h5d1 	:	val_out <= 4'h9232;
         4'h5d2 	:	val_out <= 4'h9232;
         4'h5d3 	:	val_out <= 4'h9232;
         4'h5d8 	:	val_out <= 4'h924b;
         4'h5d9 	:	val_out <= 4'h924b;
         4'h5da 	:	val_out <= 4'h924b;
         4'h5db 	:	val_out <= 4'h924b;
         4'h5e0 	:	val_out <= 4'h9264;
         4'h5e1 	:	val_out <= 4'h9264;
         4'h5e2 	:	val_out <= 4'h9264;
         4'h5e3 	:	val_out <= 4'h9264;
         4'h5e8 	:	val_out <= 4'h927d;
         4'h5e9 	:	val_out <= 4'h927d;
         4'h5ea 	:	val_out <= 4'h927d;
         4'h5eb 	:	val_out <= 4'h927d;
         4'h5f0 	:	val_out <= 4'h9296;
         4'h5f1 	:	val_out <= 4'h9296;
         4'h5f2 	:	val_out <= 4'h9296;
         4'h5f3 	:	val_out <= 4'h9296;
         4'h5f8 	:	val_out <= 4'h92af;
         4'h5f9 	:	val_out <= 4'h92af;
         4'h5fa 	:	val_out <= 4'h92af;
         4'h5fb 	:	val_out <= 4'h92af;
         4'h600 	:	val_out <= 4'h92c8;
         4'h601 	:	val_out <= 4'h92c8;
         4'h602 	:	val_out <= 4'h92c8;
         4'h603 	:	val_out <= 4'h92c8;
         4'h608 	:	val_out <= 4'h92e0;
         4'h609 	:	val_out <= 4'h92e0;
         4'h60a 	:	val_out <= 4'h92e0;
         4'h60b 	:	val_out <= 4'h92e0;
         4'h610 	:	val_out <= 4'h92f9;
         4'h611 	:	val_out <= 4'h92f9;
         4'h612 	:	val_out <= 4'h92f9;
         4'h613 	:	val_out <= 4'h92f9;
         4'h618 	:	val_out <= 4'h9312;
         4'h619 	:	val_out <= 4'h9312;
         4'h61a 	:	val_out <= 4'h9312;
         4'h61b 	:	val_out <= 4'h9312;
         4'h620 	:	val_out <= 4'h932b;
         4'h621 	:	val_out <= 4'h932b;
         4'h622 	:	val_out <= 4'h932b;
         4'h623 	:	val_out <= 4'h932b;
         4'h628 	:	val_out <= 4'h9344;
         4'h629 	:	val_out <= 4'h9344;
         4'h62a 	:	val_out <= 4'h9344;
         4'h62b 	:	val_out <= 4'h9344;
         4'h630 	:	val_out <= 4'h935d;
         4'h631 	:	val_out <= 4'h935d;
         4'h632 	:	val_out <= 4'h935d;
         4'h633 	:	val_out <= 4'h935d;
         4'h638 	:	val_out <= 4'h9376;
         4'h639 	:	val_out <= 4'h9376;
         4'h63a 	:	val_out <= 4'h9376;
         4'h63b 	:	val_out <= 4'h9376;
         4'h640 	:	val_out <= 4'h938e;
         4'h641 	:	val_out <= 4'h938e;
         4'h642 	:	val_out <= 4'h938e;
         4'h643 	:	val_out <= 4'h938e;
         4'h648 	:	val_out <= 4'h93a7;
         4'h649 	:	val_out <= 4'h93a7;
         4'h64a 	:	val_out <= 4'h93a7;
         4'h64b 	:	val_out <= 4'h93a7;
         4'h650 	:	val_out <= 4'h93c0;
         4'h651 	:	val_out <= 4'h93c0;
         4'h652 	:	val_out <= 4'h93c0;
         4'h653 	:	val_out <= 4'h93c0;
         4'h658 	:	val_out <= 4'h93d9;
         4'h659 	:	val_out <= 4'h93d9;
         4'h65a 	:	val_out <= 4'h93d9;
         4'h65b 	:	val_out <= 4'h93d9;
         4'h660 	:	val_out <= 4'h93f2;
         4'h661 	:	val_out <= 4'h93f2;
         4'h662 	:	val_out <= 4'h93f2;
         4'h663 	:	val_out <= 4'h93f2;
         4'h668 	:	val_out <= 4'h940b;
         4'h669 	:	val_out <= 4'h940b;
         4'h66a 	:	val_out <= 4'h940b;
         4'h66b 	:	val_out <= 4'h940b;
         4'h670 	:	val_out <= 4'h9423;
         4'h671 	:	val_out <= 4'h9423;
         4'h672 	:	val_out <= 4'h9423;
         4'h673 	:	val_out <= 4'h9423;
         4'h678 	:	val_out <= 4'h943c;
         4'h679 	:	val_out <= 4'h943c;
         4'h67a 	:	val_out <= 4'h943c;
         4'h67b 	:	val_out <= 4'h943c;
         4'h680 	:	val_out <= 4'h9455;
         4'h681 	:	val_out <= 4'h9455;
         4'h682 	:	val_out <= 4'h9455;
         4'h683 	:	val_out <= 4'h9455;
         4'h688 	:	val_out <= 4'h946e;
         4'h689 	:	val_out <= 4'h946e;
         4'h68a 	:	val_out <= 4'h946e;
         4'h68b 	:	val_out <= 4'h946e;
         4'h690 	:	val_out <= 4'h9487;
         4'h691 	:	val_out <= 4'h9487;
         4'h692 	:	val_out <= 4'h9487;
         4'h693 	:	val_out <= 4'h9487;
         4'h698 	:	val_out <= 4'h949f;
         4'h699 	:	val_out <= 4'h949f;
         4'h69a 	:	val_out <= 4'h949f;
         4'h69b 	:	val_out <= 4'h949f;
         4'h6a0 	:	val_out <= 4'h94b8;
         4'h6a1 	:	val_out <= 4'h94b8;
         4'h6a2 	:	val_out <= 4'h94b8;
         4'h6a3 	:	val_out <= 4'h94b8;
         4'h6a8 	:	val_out <= 4'h94d1;
         4'h6a9 	:	val_out <= 4'h94d1;
         4'h6aa 	:	val_out <= 4'h94d1;
         4'h6ab 	:	val_out <= 4'h94d1;
         4'h6b0 	:	val_out <= 4'h94ea;
         4'h6b1 	:	val_out <= 4'h94ea;
         4'h6b2 	:	val_out <= 4'h94ea;
         4'h6b3 	:	val_out <= 4'h94ea;
         4'h6b8 	:	val_out <= 4'h9503;
         4'h6b9 	:	val_out <= 4'h9503;
         4'h6ba 	:	val_out <= 4'h9503;
         4'h6bb 	:	val_out <= 4'h9503;
         4'h6c0 	:	val_out <= 4'h951b;
         4'h6c1 	:	val_out <= 4'h951b;
         4'h6c2 	:	val_out <= 4'h951b;
         4'h6c3 	:	val_out <= 4'h951b;
         4'h6c8 	:	val_out <= 4'h9534;
         4'h6c9 	:	val_out <= 4'h9534;
         4'h6ca 	:	val_out <= 4'h9534;
         4'h6cb 	:	val_out <= 4'h9534;
         4'h6d0 	:	val_out <= 4'h954d;
         4'h6d1 	:	val_out <= 4'h954d;
         4'h6d2 	:	val_out <= 4'h954d;
         4'h6d3 	:	val_out <= 4'h954d;
         4'h6d8 	:	val_out <= 4'h9566;
         4'h6d9 	:	val_out <= 4'h9566;
         4'h6da 	:	val_out <= 4'h9566;
         4'h6db 	:	val_out <= 4'h9566;
         4'h6e0 	:	val_out <= 4'h957f;
         4'h6e1 	:	val_out <= 4'h957f;
         4'h6e2 	:	val_out <= 4'h957f;
         4'h6e3 	:	val_out <= 4'h957f;
         4'h6e8 	:	val_out <= 4'h9597;
         4'h6e9 	:	val_out <= 4'h9597;
         4'h6ea 	:	val_out <= 4'h9597;
         4'h6eb 	:	val_out <= 4'h9597;
         4'h6f0 	:	val_out <= 4'h95b0;
         4'h6f1 	:	val_out <= 4'h95b0;
         4'h6f2 	:	val_out <= 4'h95b0;
         4'h6f3 	:	val_out <= 4'h95b0;
         4'h6f8 	:	val_out <= 4'h95c9;
         4'h6f9 	:	val_out <= 4'h95c9;
         4'h6fa 	:	val_out <= 4'h95c9;
         4'h6fb 	:	val_out <= 4'h95c9;
         4'h700 	:	val_out <= 4'h95e2;
         4'h701 	:	val_out <= 4'h95e2;
         4'h702 	:	val_out <= 4'h95e2;
         4'h703 	:	val_out <= 4'h95e2;
         4'h708 	:	val_out <= 4'h95fa;
         4'h709 	:	val_out <= 4'h95fa;
         4'h70a 	:	val_out <= 4'h95fa;
         4'h70b 	:	val_out <= 4'h95fa;
         4'h710 	:	val_out <= 4'h9613;
         4'h711 	:	val_out <= 4'h9613;
         4'h712 	:	val_out <= 4'h9613;
         4'h713 	:	val_out <= 4'h9613;
         4'h718 	:	val_out <= 4'h962c;
         4'h719 	:	val_out <= 4'h962c;
         4'h71a 	:	val_out <= 4'h962c;
         4'h71b 	:	val_out <= 4'h962c;
         4'h720 	:	val_out <= 4'h9645;
         4'h721 	:	val_out <= 4'h9645;
         4'h722 	:	val_out <= 4'h9645;
         4'h723 	:	val_out <= 4'h9645;
         4'h728 	:	val_out <= 4'h965d;
         4'h729 	:	val_out <= 4'h965d;
         4'h72a 	:	val_out <= 4'h965d;
         4'h72b 	:	val_out <= 4'h965d;
         4'h730 	:	val_out <= 4'h9676;
         4'h731 	:	val_out <= 4'h9676;
         4'h732 	:	val_out <= 4'h9676;
         4'h733 	:	val_out <= 4'h9676;
         4'h738 	:	val_out <= 4'h968f;
         4'h739 	:	val_out <= 4'h968f;
         4'h73a 	:	val_out <= 4'h968f;
         4'h73b 	:	val_out <= 4'h968f;
         4'h740 	:	val_out <= 4'h96a8;
         4'h741 	:	val_out <= 4'h96a8;
         4'h742 	:	val_out <= 4'h96a8;
         4'h743 	:	val_out <= 4'h96a8;
         4'h748 	:	val_out <= 4'h96c0;
         4'h749 	:	val_out <= 4'h96c0;
         4'h74a 	:	val_out <= 4'h96c0;
         4'h74b 	:	val_out <= 4'h96c0;
         4'h750 	:	val_out <= 4'h96d9;
         4'h751 	:	val_out <= 4'h96d9;
         4'h752 	:	val_out <= 4'h96d9;
         4'h753 	:	val_out <= 4'h96d9;
         4'h758 	:	val_out <= 4'h96f2;
         4'h759 	:	val_out <= 4'h96f2;
         4'h75a 	:	val_out <= 4'h96f2;
         4'h75b 	:	val_out <= 4'h96f2;
         4'h760 	:	val_out <= 4'h970a;
         4'h761 	:	val_out <= 4'h970a;
         4'h762 	:	val_out <= 4'h970a;
         4'h763 	:	val_out <= 4'h970a;
         4'h768 	:	val_out <= 4'h9723;
         4'h769 	:	val_out <= 4'h9723;
         4'h76a 	:	val_out <= 4'h9723;
         4'h76b 	:	val_out <= 4'h9723;
         4'h770 	:	val_out <= 4'h973c;
         4'h771 	:	val_out <= 4'h973c;
         4'h772 	:	val_out <= 4'h973c;
         4'h773 	:	val_out <= 4'h973c;
         4'h778 	:	val_out <= 4'h9755;
         4'h779 	:	val_out <= 4'h9755;
         4'h77a 	:	val_out <= 4'h9755;
         4'h77b 	:	val_out <= 4'h9755;
         4'h780 	:	val_out <= 4'h976d;
         4'h781 	:	val_out <= 4'h976d;
         4'h782 	:	val_out <= 4'h976d;
         4'h783 	:	val_out <= 4'h976d;
         4'h788 	:	val_out <= 4'h9786;
         4'h789 	:	val_out <= 4'h9786;
         4'h78a 	:	val_out <= 4'h9786;
         4'h78b 	:	val_out <= 4'h9786;
         4'h790 	:	val_out <= 4'h979f;
         4'h791 	:	val_out <= 4'h979f;
         4'h792 	:	val_out <= 4'h979f;
         4'h793 	:	val_out <= 4'h979f;
         4'h798 	:	val_out <= 4'h97b7;
         4'h799 	:	val_out <= 4'h97b7;
         4'h79a 	:	val_out <= 4'h97b7;
         4'h79b 	:	val_out <= 4'h97b7;
         4'h7a0 	:	val_out <= 4'h97d0;
         4'h7a1 	:	val_out <= 4'h97d0;
         4'h7a2 	:	val_out <= 4'h97d0;
         4'h7a3 	:	val_out <= 4'h97d0;
         4'h7a8 	:	val_out <= 4'h97e9;
         4'h7a9 	:	val_out <= 4'h97e9;
         4'h7aa 	:	val_out <= 4'h97e9;
         4'h7ab 	:	val_out <= 4'h97e9;
         4'h7b0 	:	val_out <= 4'h9802;
         4'h7b1 	:	val_out <= 4'h9802;
         4'h7b2 	:	val_out <= 4'h9802;
         4'h7b3 	:	val_out <= 4'h9802;
         4'h7b8 	:	val_out <= 4'h981a;
         4'h7b9 	:	val_out <= 4'h981a;
         4'h7ba 	:	val_out <= 4'h981a;
         4'h7bb 	:	val_out <= 4'h981a;
         4'h7c0 	:	val_out <= 4'h9833;
         4'h7c1 	:	val_out <= 4'h9833;
         4'h7c2 	:	val_out <= 4'h9833;
         4'h7c3 	:	val_out <= 4'h9833;
         4'h7c8 	:	val_out <= 4'h984c;
         4'h7c9 	:	val_out <= 4'h984c;
         4'h7ca 	:	val_out <= 4'h984c;
         4'h7cb 	:	val_out <= 4'h984c;
         4'h7d0 	:	val_out <= 4'h9864;
         4'h7d1 	:	val_out <= 4'h9864;
         4'h7d2 	:	val_out <= 4'h9864;
         4'h7d3 	:	val_out <= 4'h9864;
         4'h7d8 	:	val_out <= 4'h987d;
         4'h7d9 	:	val_out <= 4'h987d;
         4'h7da 	:	val_out <= 4'h987d;
         4'h7db 	:	val_out <= 4'h987d;
         4'h7e0 	:	val_out <= 4'h9896;
         4'h7e1 	:	val_out <= 4'h9896;
         4'h7e2 	:	val_out <= 4'h9896;
         4'h7e3 	:	val_out <= 4'h9896;
         4'h7e8 	:	val_out <= 4'h98ae;
         4'h7e9 	:	val_out <= 4'h98ae;
         4'h7ea 	:	val_out <= 4'h98ae;
         4'h7eb 	:	val_out <= 4'h98ae;
         4'h7f0 	:	val_out <= 4'h98c7;
         4'h7f1 	:	val_out <= 4'h98c7;
         4'h7f2 	:	val_out <= 4'h98c7;
         4'h7f3 	:	val_out <= 4'h98c7;
         4'h7f8 	:	val_out <= 4'h98e0;
         4'h7f9 	:	val_out <= 4'h98e0;
         4'h7fa 	:	val_out <= 4'h98e0;
         4'h7fb 	:	val_out <= 4'h98e0;
         4'h800 	:	val_out <= 4'h98f8;
         4'h801 	:	val_out <= 4'h98f8;
         4'h802 	:	val_out <= 4'h98f8;
         4'h803 	:	val_out <= 4'h98f8;
         4'h808 	:	val_out <= 4'h9911;
         4'h809 	:	val_out <= 4'h9911;
         4'h80a 	:	val_out <= 4'h9911;
         4'h80b 	:	val_out <= 4'h9911;
         4'h810 	:	val_out <= 4'h992a;
         4'h811 	:	val_out <= 4'h992a;
         4'h812 	:	val_out <= 4'h992a;
         4'h813 	:	val_out <= 4'h992a;
         4'h818 	:	val_out <= 4'h9942;
         4'h819 	:	val_out <= 4'h9942;
         4'h81a 	:	val_out <= 4'h9942;
         4'h81b 	:	val_out <= 4'h9942;
         4'h820 	:	val_out <= 4'h995b;
         4'h821 	:	val_out <= 4'h995b;
         4'h822 	:	val_out <= 4'h995b;
         4'h823 	:	val_out <= 4'h995b;
         4'h828 	:	val_out <= 4'h9973;
         4'h829 	:	val_out <= 4'h9973;
         4'h82a 	:	val_out <= 4'h9973;
         4'h82b 	:	val_out <= 4'h9973;
         4'h830 	:	val_out <= 4'h998c;
         4'h831 	:	val_out <= 4'h998c;
         4'h832 	:	val_out <= 4'h998c;
         4'h833 	:	val_out <= 4'h998c;
         4'h838 	:	val_out <= 4'h99a5;
         4'h839 	:	val_out <= 4'h99a5;
         4'h83a 	:	val_out <= 4'h99a5;
         4'h83b 	:	val_out <= 4'h99a5;
         4'h840 	:	val_out <= 4'h99bd;
         4'h841 	:	val_out <= 4'h99bd;
         4'h842 	:	val_out <= 4'h99bd;
         4'h843 	:	val_out <= 4'h99bd;
         4'h848 	:	val_out <= 4'h99d6;
         4'h849 	:	val_out <= 4'h99d6;
         4'h84a 	:	val_out <= 4'h99d6;
         4'h84b 	:	val_out <= 4'h99d6;
         4'h850 	:	val_out <= 4'h99ef;
         4'h851 	:	val_out <= 4'h99ef;
         4'h852 	:	val_out <= 4'h99ef;
         4'h853 	:	val_out <= 4'h99ef;
         4'h858 	:	val_out <= 4'h9a07;
         4'h859 	:	val_out <= 4'h9a07;
         4'h85a 	:	val_out <= 4'h9a07;
         4'h85b 	:	val_out <= 4'h9a07;
         4'h860 	:	val_out <= 4'h9a20;
         4'h861 	:	val_out <= 4'h9a20;
         4'h862 	:	val_out <= 4'h9a20;
         4'h863 	:	val_out <= 4'h9a20;
         4'h868 	:	val_out <= 4'h9a38;
         4'h869 	:	val_out <= 4'h9a38;
         4'h86a 	:	val_out <= 4'h9a38;
         4'h86b 	:	val_out <= 4'h9a38;
         4'h870 	:	val_out <= 4'h9a51;
         4'h871 	:	val_out <= 4'h9a51;
         4'h872 	:	val_out <= 4'h9a51;
         4'h873 	:	val_out <= 4'h9a51;
         4'h878 	:	val_out <= 4'h9a6a;
         4'h879 	:	val_out <= 4'h9a6a;
         4'h87a 	:	val_out <= 4'h9a6a;
         4'h87b 	:	val_out <= 4'h9a6a;
         4'h880 	:	val_out <= 4'h9a82;
         4'h881 	:	val_out <= 4'h9a82;
         4'h882 	:	val_out <= 4'h9a82;
         4'h883 	:	val_out <= 4'h9a82;
         4'h888 	:	val_out <= 4'h9a9b;
         4'h889 	:	val_out <= 4'h9a9b;
         4'h88a 	:	val_out <= 4'h9a9b;
         4'h88b 	:	val_out <= 4'h9a9b;
         4'h890 	:	val_out <= 4'h9ab3;
         4'h891 	:	val_out <= 4'h9ab3;
         4'h892 	:	val_out <= 4'h9ab3;
         4'h893 	:	val_out <= 4'h9ab3;
         4'h898 	:	val_out <= 4'h9acc;
         4'h899 	:	val_out <= 4'h9acc;
         4'h89a 	:	val_out <= 4'h9acc;
         4'h89b 	:	val_out <= 4'h9acc;
         4'h8a0 	:	val_out <= 4'h9ae4;
         4'h8a1 	:	val_out <= 4'h9ae4;
         4'h8a2 	:	val_out <= 4'h9ae4;
         4'h8a3 	:	val_out <= 4'h9ae4;
         4'h8a8 	:	val_out <= 4'h9afd;
         4'h8a9 	:	val_out <= 4'h9afd;
         4'h8aa 	:	val_out <= 4'h9afd;
         4'h8ab 	:	val_out <= 4'h9afd;
         4'h8b0 	:	val_out <= 4'h9b16;
         4'h8b1 	:	val_out <= 4'h9b16;
         4'h8b2 	:	val_out <= 4'h9b16;
         4'h8b3 	:	val_out <= 4'h9b16;
         4'h8b8 	:	val_out <= 4'h9b2e;
         4'h8b9 	:	val_out <= 4'h9b2e;
         4'h8ba 	:	val_out <= 4'h9b2e;
         4'h8bb 	:	val_out <= 4'h9b2e;
         4'h8c0 	:	val_out <= 4'h9b47;
         4'h8c1 	:	val_out <= 4'h9b47;
         4'h8c2 	:	val_out <= 4'h9b47;
         4'h8c3 	:	val_out <= 4'h9b47;
         4'h8c8 	:	val_out <= 4'h9b5f;
         4'h8c9 	:	val_out <= 4'h9b5f;
         4'h8ca 	:	val_out <= 4'h9b5f;
         4'h8cb 	:	val_out <= 4'h9b5f;
         4'h8d0 	:	val_out <= 4'h9b78;
         4'h8d1 	:	val_out <= 4'h9b78;
         4'h8d2 	:	val_out <= 4'h9b78;
         4'h8d3 	:	val_out <= 4'h9b78;
         4'h8d8 	:	val_out <= 4'h9b90;
         4'h8d9 	:	val_out <= 4'h9b90;
         4'h8da 	:	val_out <= 4'h9b90;
         4'h8db 	:	val_out <= 4'h9b90;
         4'h8e0 	:	val_out <= 4'h9ba9;
         4'h8e1 	:	val_out <= 4'h9ba9;
         4'h8e2 	:	val_out <= 4'h9ba9;
         4'h8e3 	:	val_out <= 4'h9ba9;
         4'h8e8 	:	val_out <= 4'h9bc1;
         4'h8e9 	:	val_out <= 4'h9bc1;
         4'h8ea 	:	val_out <= 4'h9bc1;
         4'h8eb 	:	val_out <= 4'h9bc1;
         4'h8f0 	:	val_out <= 4'h9bda;
         4'h8f1 	:	val_out <= 4'h9bda;
         4'h8f2 	:	val_out <= 4'h9bda;
         4'h8f3 	:	val_out <= 4'h9bda;
         4'h8f8 	:	val_out <= 4'h9bf2;
         4'h8f9 	:	val_out <= 4'h9bf2;
         4'h8fa 	:	val_out <= 4'h9bf2;
         4'h8fb 	:	val_out <= 4'h9bf2;
         4'h900 	:	val_out <= 4'h9c0b;
         4'h901 	:	val_out <= 4'h9c0b;
         4'h902 	:	val_out <= 4'h9c0b;
         4'h903 	:	val_out <= 4'h9c0b;
         4'h908 	:	val_out <= 4'h9c24;
         4'h909 	:	val_out <= 4'h9c24;
         4'h90a 	:	val_out <= 4'h9c24;
         4'h90b 	:	val_out <= 4'h9c24;
         4'h910 	:	val_out <= 4'h9c3c;
         4'h911 	:	val_out <= 4'h9c3c;
         4'h912 	:	val_out <= 4'h9c3c;
         4'h913 	:	val_out <= 4'h9c3c;
         4'h918 	:	val_out <= 4'h9c55;
         4'h919 	:	val_out <= 4'h9c55;
         4'h91a 	:	val_out <= 4'h9c55;
         4'h91b 	:	val_out <= 4'h9c55;
         4'h920 	:	val_out <= 4'h9c6d;
         4'h921 	:	val_out <= 4'h9c6d;
         4'h922 	:	val_out <= 4'h9c6d;
         4'h923 	:	val_out <= 4'h9c6d;
         4'h928 	:	val_out <= 4'h9c86;
         4'h929 	:	val_out <= 4'h9c86;
         4'h92a 	:	val_out <= 4'h9c86;
         4'h92b 	:	val_out <= 4'h9c86;
         4'h930 	:	val_out <= 4'h9c9e;
         4'h931 	:	val_out <= 4'h9c9e;
         4'h932 	:	val_out <= 4'h9c9e;
         4'h933 	:	val_out <= 4'h9c9e;
         4'h938 	:	val_out <= 4'h9cb7;
         4'h939 	:	val_out <= 4'h9cb7;
         4'h93a 	:	val_out <= 4'h9cb7;
         4'h93b 	:	val_out <= 4'h9cb7;
         4'h940 	:	val_out <= 4'h9ccf;
         4'h941 	:	val_out <= 4'h9ccf;
         4'h942 	:	val_out <= 4'h9ccf;
         4'h943 	:	val_out <= 4'h9ccf;
         4'h948 	:	val_out <= 4'h9ce8;
         4'h949 	:	val_out <= 4'h9ce8;
         4'h94a 	:	val_out <= 4'h9ce8;
         4'h94b 	:	val_out <= 4'h9ce8;
         4'h950 	:	val_out <= 4'h9d00;
         4'h951 	:	val_out <= 4'h9d00;
         4'h952 	:	val_out <= 4'h9d00;
         4'h953 	:	val_out <= 4'h9d00;
         4'h958 	:	val_out <= 4'h9d18;
         4'h959 	:	val_out <= 4'h9d18;
         4'h95a 	:	val_out <= 4'h9d18;
         4'h95b 	:	val_out <= 4'h9d18;
         4'h960 	:	val_out <= 4'h9d31;
         4'h961 	:	val_out <= 4'h9d31;
         4'h962 	:	val_out <= 4'h9d31;
         4'h963 	:	val_out <= 4'h9d31;
         4'h968 	:	val_out <= 4'h9d49;
         4'h969 	:	val_out <= 4'h9d49;
         4'h96a 	:	val_out <= 4'h9d49;
         4'h96b 	:	val_out <= 4'h9d49;
         4'h970 	:	val_out <= 4'h9d62;
         4'h971 	:	val_out <= 4'h9d62;
         4'h972 	:	val_out <= 4'h9d62;
         4'h973 	:	val_out <= 4'h9d62;
         4'h978 	:	val_out <= 4'h9d7a;
         4'h979 	:	val_out <= 4'h9d7a;
         4'h97a 	:	val_out <= 4'h9d7a;
         4'h97b 	:	val_out <= 4'h9d7a;
         4'h980 	:	val_out <= 4'h9d93;
         4'h981 	:	val_out <= 4'h9d93;
         4'h982 	:	val_out <= 4'h9d93;
         4'h983 	:	val_out <= 4'h9d93;
         4'h988 	:	val_out <= 4'h9dab;
         4'h989 	:	val_out <= 4'h9dab;
         4'h98a 	:	val_out <= 4'h9dab;
         4'h98b 	:	val_out <= 4'h9dab;
         4'h990 	:	val_out <= 4'h9dc4;
         4'h991 	:	val_out <= 4'h9dc4;
         4'h992 	:	val_out <= 4'h9dc4;
         4'h993 	:	val_out <= 4'h9dc4;
         4'h998 	:	val_out <= 4'h9ddc;
         4'h999 	:	val_out <= 4'h9ddc;
         4'h99a 	:	val_out <= 4'h9ddc;
         4'h99b 	:	val_out <= 4'h9ddc;
         4'h9a0 	:	val_out <= 4'h9df5;
         4'h9a1 	:	val_out <= 4'h9df5;
         4'h9a2 	:	val_out <= 4'h9df5;
         4'h9a3 	:	val_out <= 4'h9df5;
         4'h9a8 	:	val_out <= 4'h9e0d;
         4'h9a9 	:	val_out <= 4'h9e0d;
         4'h9aa 	:	val_out <= 4'h9e0d;
         4'h9ab 	:	val_out <= 4'h9e0d;
         4'h9b0 	:	val_out <= 4'h9e25;
         4'h9b1 	:	val_out <= 4'h9e25;
         4'h9b2 	:	val_out <= 4'h9e25;
         4'h9b3 	:	val_out <= 4'h9e25;
         4'h9b8 	:	val_out <= 4'h9e3e;
         4'h9b9 	:	val_out <= 4'h9e3e;
         4'h9ba 	:	val_out <= 4'h9e3e;
         4'h9bb 	:	val_out <= 4'h9e3e;
         4'h9c0 	:	val_out <= 4'h9e56;
         4'h9c1 	:	val_out <= 4'h9e56;
         4'h9c2 	:	val_out <= 4'h9e56;
         4'h9c3 	:	val_out <= 4'h9e56;
         4'h9c8 	:	val_out <= 4'h9e6f;
         4'h9c9 	:	val_out <= 4'h9e6f;
         4'h9ca 	:	val_out <= 4'h9e6f;
         4'h9cb 	:	val_out <= 4'h9e6f;
         4'h9d0 	:	val_out <= 4'h9e87;
         4'h9d1 	:	val_out <= 4'h9e87;
         4'h9d2 	:	val_out <= 4'h9e87;
         4'h9d3 	:	val_out <= 4'h9e87;
         4'h9d8 	:	val_out <= 4'h9ea0;
         4'h9d9 	:	val_out <= 4'h9ea0;
         4'h9da 	:	val_out <= 4'h9ea0;
         4'h9db 	:	val_out <= 4'h9ea0;
         4'h9e0 	:	val_out <= 4'h9eb8;
         4'h9e1 	:	val_out <= 4'h9eb8;
         4'h9e2 	:	val_out <= 4'h9eb8;
         4'h9e3 	:	val_out <= 4'h9eb8;
         4'h9e8 	:	val_out <= 4'h9ed0;
         4'h9e9 	:	val_out <= 4'h9ed0;
         4'h9ea 	:	val_out <= 4'h9ed0;
         4'h9eb 	:	val_out <= 4'h9ed0;
         4'h9f0 	:	val_out <= 4'h9ee9;
         4'h9f1 	:	val_out <= 4'h9ee9;
         4'h9f2 	:	val_out <= 4'h9ee9;
         4'h9f3 	:	val_out <= 4'h9ee9;
         4'h9f8 	:	val_out <= 4'h9f01;
         4'h9f9 	:	val_out <= 4'h9f01;
         4'h9fa 	:	val_out <= 4'h9f01;
         4'h9fb 	:	val_out <= 4'h9f01;
         4'ha00 	:	val_out <= 4'h9f19;
         4'ha01 	:	val_out <= 4'h9f19;
         4'ha02 	:	val_out <= 4'h9f19;
         4'ha03 	:	val_out <= 4'h9f19;
         4'ha08 	:	val_out <= 4'h9f32;
         4'ha09 	:	val_out <= 4'h9f32;
         4'ha0a 	:	val_out <= 4'h9f32;
         4'ha0b 	:	val_out <= 4'h9f32;
         4'ha10 	:	val_out <= 4'h9f4a;
         4'ha11 	:	val_out <= 4'h9f4a;
         4'ha12 	:	val_out <= 4'h9f4a;
         4'ha13 	:	val_out <= 4'h9f4a;
         4'ha18 	:	val_out <= 4'h9f63;
         4'ha19 	:	val_out <= 4'h9f63;
         4'ha1a 	:	val_out <= 4'h9f63;
         4'ha1b 	:	val_out <= 4'h9f63;
         4'ha20 	:	val_out <= 4'h9f7b;
         4'ha21 	:	val_out <= 4'h9f7b;
         4'ha22 	:	val_out <= 4'h9f7b;
         4'ha23 	:	val_out <= 4'h9f7b;
         4'ha28 	:	val_out <= 4'h9f93;
         4'ha29 	:	val_out <= 4'h9f93;
         4'ha2a 	:	val_out <= 4'h9f93;
         4'ha2b 	:	val_out <= 4'h9f93;
         4'ha30 	:	val_out <= 4'h9fac;
         4'ha31 	:	val_out <= 4'h9fac;
         4'ha32 	:	val_out <= 4'h9fac;
         4'ha33 	:	val_out <= 4'h9fac;
         4'ha38 	:	val_out <= 4'h9fc4;
         4'ha39 	:	val_out <= 4'h9fc4;
         4'ha3a 	:	val_out <= 4'h9fc4;
         4'ha3b 	:	val_out <= 4'h9fc4;
         4'ha40 	:	val_out <= 4'h9fdc;
         4'ha41 	:	val_out <= 4'h9fdc;
         4'ha42 	:	val_out <= 4'h9fdc;
         4'ha43 	:	val_out <= 4'h9fdc;
         4'ha48 	:	val_out <= 4'h9ff5;
         4'ha49 	:	val_out <= 4'h9ff5;
         4'ha4a 	:	val_out <= 4'h9ff5;
         4'ha4b 	:	val_out <= 4'h9ff5;
         4'ha50 	:	val_out <= 4'ha00d;
         4'ha51 	:	val_out <= 4'ha00d;
         4'ha52 	:	val_out <= 4'ha00d;
         4'ha53 	:	val_out <= 4'ha00d;
         4'ha58 	:	val_out <= 4'ha025;
         4'ha59 	:	val_out <= 4'ha025;
         4'ha5a 	:	val_out <= 4'ha025;
         4'ha5b 	:	val_out <= 4'ha025;
         4'ha60 	:	val_out <= 4'ha03e;
         4'ha61 	:	val_out <= 4'ha03e;
         4'ha62 	:	val_out <= 4'ha03e;
         4'ha63 	:	val_out <= 4'ha03e;
         4'ha68 	:	val_out <= 4'ha056;
         4'ha69 	:	val_out <= 4'ha056;
         4'ha6a 	:	val_out <= 4'ha056;
         4'ha6b 	:	val_out <= 4'ha056;
         4'ha70 	:	val_out <= 4'ha06e;
         4'ha71 	:	val_out <= 4'ha06e;
         4'ha72 	:	val_out <= 4'ha06e;
         4'ha73 	:	val_out <= 4'ha06e;
         4'ha78 	:	val_out <= 4'ha087;
         4'ha79 	:	val_out <= 4'ha087;
         4'ha7a 	:	val_out <= 4'ha087;
         4'ha7b 	:	val_out <= 4'ha087;
         4'ha80 	:	val_out <= 4'ha09f;
         4'ha81 	:	val_out <= 4'ha09f;
         4'ha82 	:	val_out <= 4'ha09f;
         4'ha83 	:	val_out <= 4'ha09f;
         4'ha88 	:	val_out <= 4'ha0b7;
         4'ha89 	:	val_out <= 4'ha0b7;
         4'ha8a 	:	val_out <= 4'ha0b7;
         4'ha8b 	:	val_out <= 4'ha0b7;
         4'ha90 	:	val_out <= 4'ha0d0;
         4'ha91 	:	val_out <= 4'ha0d0;
         4'ha92 	:	val_out <= 4'ha0d0;
         4'ha93 	:	val_out <= 4'ha0d0;
         4'ha98 	:	val_out <= 4'ha0e8;
         4'ha99 	:	val_out <= 4'ha0e8;
         4'ha9a 	:	val_out <= 4'ha0e8;
         4'ha9b 	:	val_out <= 4'ha0e8;
         4'haa0 	:	val_out <= 4'ha100;
         4'haa1 	:	val_out <= 4'ha100;
         4'haa2 	:	val_out <= 4'ha100;
         4'haa3 	:	val_out <= 4'ha100;
         4'haa8 	:	val_out <= 4'ha118;
         4'haa9 	:	val_out <= 4'ha118;
         4'haaa 	:	val_out <= 4'ha118;
         4'haab 	:	val_out <= 4'ha118;
         4'hab0 	:	val_out <= 4'ha131;
         4'hab1 	:	val_out <= 4'ha131;
         4'hab2 	:	val_out <= 4'ha131;
         4'hab3 	:	val_out <= 4'ha131;
         4'hab8 	:	val_out <= 4'ha149;
         4'hab9 	:	val_out <= 4'ha149;
         4'haba 	:	val_out <= 4'ha149;
         4'habb 	:	val_out <= 4'ha149;
         4'hac0 	:	val_out <= 4'ha161;
         4'hac1 	:	val_out <= 4'ha161;
         4'hac2 	:	val_out <= 4'ha161;
         4'hac3 	:	val_out <= 4'ha161;
         4'hac8 	:	val_out <= 4'ha179;
         4'hac9 	:	val_out <= 4'ha179;
         4'haca 	:	val_out <= 4'ha179;
         4'hacb 	:	val_out <= 4'ha179;
         4'had0 	:	val_out <= 4'ha192;
         4'had1 	:	val_out <= 4'ha192;
         4'had2 	:	val_out <= 4'ha192;
         4'had3 	:	val_out <= 4'ha192;
         4'had8 	:	val_out <= 4'ha1aa;
         4'had9 	:	val_out <= 4'ha1aa;
         4'hada 	:	val_out <= 4'ha1aa;
         4'hadb 	:	val_out <= 4'ha1aa;
         4'hae0 	:	val_out <= 4'ha1c2;
         4'hae1 	:	val_out <= 4'ha1c2;
         4'hae2 	:	val_out <= 4'ha1c2;
         4'hae3 	:	val_out <= 4'ha1c2;
         4'hae8 	:	val_out <= 4'ha1da;
         4'hae9 	:	val_out <= 4'ha1da;
         4'haea 	:	val_out <= 4'ha1da;
         4'haeb 	:	val_out <= 4'ha1da;
         4'haf0 	:	val_out <= 4'ha1f3;
         4'haf1 	:	val_out <= 4'ha1f3;
         4'haf2 	:	val_out <= 4'ha1f3;
         4'haf3 	:	val_out <= 4'ha1f3;
         4'haf8 	:	val_out <= 4'ha20b;
         4'haf9 	:	val_out <= 4'ha20b;
         4'hafa 	:	val_out <= 4'ha20b;
         4'hafb 	:	val_out <= 4'ha20b;
         4'hb00 	:	val_out <= 4'ha223;
         4'hb01 	:	val_out <= 4'ha223;
         4'hb02 	:	val_out <= 4'ha223;
         4'hb03 	:	val_out <= 4'ha223;
         4'hb08 	:	val_out <= 4'ha23b;
         4'hb09 	:	val_out <= 4'ha23b;
         4'hb0a 	:	val_out <= 4'ha23b;
         4'hb0b 	:	val_out <= 4'ha23b;
         4'hb10 	:	val_out <= 4'ha254;
         4'hb11 	:	val_out <= 4'ha254;
         4'hb12 	:	val_out <= 4'ha254;
         4'hb13 	:	val_out <= 4'ha254;
         4'hb18 	:	val_out <= 4'ha26c;
         4'hb19 	:	val_out <= 4'ha26c;
         4'hb1a 	:	val_out <= 4'ha26c;
         4'hb1b 	:	val_out <= 4'ha26c;
         4'hb20 	:	val_out <= 4'ha284;
         4'hb21 	:	val_out <= 4'ha284;
         4'hb22 	:	val_out <= 4'ha284;
         4'hb23 	:	val_out <= 4'ha284;
         4'hb28 	:	val_out <= 4'ha29c;
         4'hb29 	:	val_out <= 4'ha29c;
         4'hb2a 	:	val_out <= 4'ha29c;
         4'hb2b 	:	val_out <= 4'ha29c;
         4'hb30 	:	val_out <= 4'ha2b4;
         4'hb31 	:	val_out <= 4'ha2b4;
         4'hb32 	:	val_out <= 4'ha2b4;
         4'hb33 	:	val_out <= 4'ha2b4;
         4'hb38 	:	val_out <= 4'ha2cd;
         4'hb39 	:	val_out <= 4'ha2cd;
         4'hb3a 	:	val_out <= 4'ha2cd;
         4'hb3b 	:	val_out <= 4'ha2cd;
         4'hb40 	:	val_out <= 4'ha2e5;
         4'hb41 	:	val_out <= 4'ha2e5;
         4'hb42 	:	val_out <= 4'ha2e5;
         4'hb43 	:	val_out <= 4'ha2e5;
         4'hb48 	:	val_out <= 4'ha2fd;
         4'hb49 	:	val_out <= 4'ha2fd;
         4'hb4a 	:	val_out <= 4'ha2fd;
         4'hb4b 	:	val_out <= 4'ha2fd;
         4'hb50 	:	val_out <= 4'ha315;
         4'hb51 	:	val_out <= 4'ha315;
         4'hb52 	:	val_out <= 4'ha315;
         4'hb53 	:	val_out <= 4'ha315;
         4'hb58 	:	val_out <= 4'ha32d;
         4'hb59 	:	val_out <= 4'ha32d;
         4'hb5a 	:	val_out <= 4'ha32d;
         4'hb5b 	:	val_out <= 4'ha32d;
         4'hb60 	:	val_out <= 4'ha345;
         4'hb61 	:	val_out <= 4'ha345;
         4'hb62 	:	val_out <= 4'ha345;
         4'hb63 	:	val_out <= 4'ha345;
         4'hb68 	:	val_out <= 4'ha35e;
         4'hb69 	:	val_out <= 4'ha35e;
         4'hb6a 	:	val_out <= 4'ha35e;
         4'hb6b 	:	val_out <= 4'ha35e;
         4'hb70 	:	val_out <= 4'ha376;
         4'hb71 	:	val_out <= 4'ha376;
         4'hb72 	:	val_out <= 4'ha376;
         4'hb73 	:	val_out <= 4'ha376;
         4'hb78 	:	val_out <= 4'ha38e;
         4'hb79 	:	val_out <= 4'ha38e;
         4'hb7a 	:	val_out <= 4'ha38e;
         4'hb7b 	:	val_out <= 4'ha38e;
         4'hb80 	:	val_out <= 4'ha3a6;
         4'hb81 	:	val_out <= 4'ha3a6;
         4'hb82 	:	val_out <= 4'ha3a6;
         4'hb83 	:	val_out <= 4'ha3a6;
         4'hb88 	:	val_out <= 4'ha3be;
         4'hb89 	:	val_out <= 4'ha3be;
         4'hb8a 	:	val_out <= 4'ha3be;
         4'hb8b 	:	val_out <= 4'ha3be;
         4'hb90 	:	val_out <= 4'ha3d6;
         4'hb91 	:	val_out <= 4'ha3d6;
         4'hb92 	:	val_out <= 4'ha3d6;
         4'hb93 	:	val_out <= 4'ha3d6;
         4'hb98 	:	val_out <= 4'ha3ee;
         4'hb99 	:	val_out <= 4'ha3ee;
         4'hb9a 	:	val_out <= 4'ha3ee;
         4'hb9b 	:	val_out <= 4'ha3ee;
         4'hba0 	:	val_out <= 4'ha407;
         4'hba1 	:	val_out <= 4'ha407;
         4'hba2 	:	val_out <= 4'ha407;
         4'hba3 	:	val_out <= 4'ha407;
         4'hba8 	:	val_out <= 4'ha41f;
         4'hba9 	:	val_out <= 4'ha41f;
         4'hbaa 	:	val_out <= 4'ha41f;
         4'hbab 	:	val_out <= 4'ha41f;
         4'hbb0 	:	val_out <= 4'ha437;
         4'hbb1 	:	val_out <= 4'ha437;
         4'hbb2 	:	val_out <= 4'ha437;
         4'hbb3 	:	val_out <= 4'ha437;
         4'hbb8 	:	val_out <= 4'ha44f;
         4'hbb9 	:	val_out <= 4'ha44f;
         4'hbba 	:	val_out <= 4'ha44f;
         4'hbbb 	:	val_out <= 4'ha44f;
         4'hbc0 	:	val_out <= 4'ha467;
         4'hbc1 	:	val_out <= 4'ha467;
         4'hbc2 	:	val_out <= 4'ha467;
         4'hbc3 	:	val_out <= 4'ha467;
         4'hbc8 	:	val_out <= 4'ha47f;
         4'hbc9 	:	val_out <= 4'ha47f;
         4'hbca 	:	val_out <= 4'ha47f;
         4'hbcb 	:	val_out <= 4'ha47f;
         4'hbd0 	:	val_out <= 4'ha497;
         4'hbd1 	:	val_out <= 4'ha497;
         4'hbd2 	:	val_out <= 4'ha497;
         4'hbd3 	:	val_out <= 4'ha497;
         4'hbd8 	:	val_out <= 4'ha4af;
         4'hbd9 	:	val_out <= 4'ha4af;
         4'hbda 	:	val_out <= 4'ha4af;
         4'hbdb 	:	val_out <= 4'ha4af;
         4'hbe0 	:	val_out <= 4'ha4c7;
         4'hbe1 	:	val_out <= 4'ha4c7;
         4'hbe2 	:	val_out <= 4'ha4c7;
         4'hbe3 	:	val_out <= 4'ha4c7;
         4'hbe8 	:	val_out <= 4'ha4df;
         4'hbe9 	:	val_out <= 4'ha4df;
         4'hbea 	:	val_out <= 4'ha4df;
         4'hbeb 	:	val_out <= 4'ha4df;
         4'hbf0 	:	val_out <= 4'ha4f7;
         4'hbf1 	:	val_out <= 4'ha4f7;
         4'hbf2 	:	val_out <= 4'ha4f7;
         4'hbf3 	:	val_out <= 4'ha4f7;
         4'hbf8 	:	val_out <= 4'ha50f;
         4'hbf9 	:	val_out <= 4'ha50f;
         4'hbfa 	:	val_out <= 4'ha50f;
         4'hbfb 	:	val_out <= 4'ha50f;
         4'hc00 	:	val_out <= 4'ha528;
         4'hc01 	:	val_out <= 4'ha528;
         4'hc02 	:	val_out <= 4'ha528;
         4'hc03 	:	val_out <= 4'ha528;
         4'hc08 	:	val_out <= 4'ha540;
         4'hc09 	:	val_out <= 4'ha540;
         4'hc0a 	:	val_out <= 4'ha540;
         4'hc0b 	:	val_out <= 4'ha540;
         4'hc10 	:	val_out <= 4'ha558;
         4'hc11 	:	val_out <= 4'ha558;
         4'hc12 	:	val_out <= 4'ha558;
         4'hc13 	:	val_out <= 4'ha558;
         4'hc18 	:	val_out <= 4'ha570;
         4'hc19 	:	val_out <= 4'ha570;
         4'hc1a 	:	val_out <= 4'ha570;
         4'hc1b 	:	val_out <= 4'ha570;
         4'hc20 	:	val_out <= 4'ha588;
         4'hc21 	:	val_out <= 4'ha588;
         4'hc22 	:	val_out <= 4'ha588;
         4'hc23 	:	val_out <= 4'ha588;
         4'hc28 	:	val_out <= 4'ha5a0;
         4'hc29 	:	val_out <= 4'ha5a0;
         4'hc2a 	:	val_out <= 4'ha5a0;
         4'hc2b 	:	val_out <= 4'ha5a0;
         4'hc30 	:	val_out <= 4'ha5b8;
         4'hc31 	:	val_out <= 4'ha5b8;
         4'hc32 	:	val_out <= 4'ha5b8;
         4'hc33 	:	val_out <= 4'ha5b8;
         4'hc38 	:	val_out <= 4'ha5d0;
         4'hc39 	:	val_out <= 4'ha5d0;
         4'hc3a 	:	val_out <= 4'ha5d0;
         4'hc3b 	:	val_out <= 4'ha5d0;
         4'hc40 	:	val_out <= 4'ha5e8;
         4'hc41 	:	val_out <= 4'ha5e8;
         4'hc42 	:	val_out <= 4'ha5e8;
         4'hc43 	:	val_out <= 4'ha5e8;
         4'hc48 	:	val_out <= 4'ha600;
         4'hc49 	:	val_out <= 4'ha600;
         4'hc4a 	:	val_out <= 4'ha600;
         4'hc4b 	:	val_out <= 4'ha600;
         4'hc50 	:	val_out <= 4'ha618;
         4'hc51 	:	val_out <= 4'ha618;
         4'hc52 	:	val_out <= 4'ha618;
         4'hc53 	:	val_out <= 4'ha618;
         4'hc58 	:	val_out <= 4'ha630;
         4'hc59 	:	val_out <= 4'ha630;
         4'hc5a 	:	val_out <= 4'ha630;
         4'hc5b 	:	val_out <= 4'ha630;
         4'hc60 	:	val_out <= 4'ha648;
         4'hc61 	:	val_out <= 4'ha648;
         4'hc62 	:	val_out <= 4'ha648;
         4'hc63 	:	val_out <= 4'ha648;
         4'hc68 	:	val_out <= 4'ha660;
         4'hc69 	:	val_out <= 4'ha660;
         4'hc6a 	:	val_out <= 4'ha660;
         4'hc6b 	:	val_out <= 4'ha660;
         4'hc70 	:	val_out <= 4'ha678;
         4'hc71 	:	val_out <= 4'ha678;
         4'hc72 	:	val_out <= 4'ha678;
         4'hc73 	:	val_out <= 4'ha678;
         4'hc78 	:	val_out <= 4'ha690;
         4'hc79 	:	val_out <= 4'ha690;
         4'hc7a 	:	val_out <= 4'ha690;
         4'hc7b 	:	val_out <= 4'ha690;
         4'hc80 	:	val_out <= 4'ha6a8;
         4'hc81 	:	val_out <= 4'ha6a8;
         4'hc82 	:	val_out <= 4'ha6a8;
         4'hc83 	:	val_out <= 4'ha6a8;
         4'hc88 	:	val_out <= 4'ha6c0;
         4'hc89 	:	val_out <= 4'ha6c0;
         4'hc8a 	:	val_out <= 4'ha6c0;
         4'hc8b 	:	val_out <= 4'ha6c0;
         4'hc90 	:	val_out <= 4'ha6d8;
         4'hc91 	:	val_out <= 4'ha6d8;
         4'hc92 	:	val_out <= 4'ha6d8;
         4'hc93 	:	val_out <= 4'ha6d8;
         4'hc98 	:	val_out <= 4'ha6ef;
         4'hc99 	:	val_out <= 4'ha6ef;
         4'hc9a 	:	val_out <= 4'ha6ef;
         4'hc9b 	:	val_out <= 4'ha6ef;
         4'hca0 	:	val_out <= 4'ha707;
         4'hca1 	:	val_out <= 4'ha707;
         4'hca2 	:	val_out <= 4'ha707;
         4'hca3 	:	val_out <= 4'ha707;
         4'hca8 	:	val_out <= 4'ha71f;
         4'hca9 	:	val_out <= 4'ha71f;
         4'hcaa 	:	val_out <= 4'ha71f;
         4'hcab 	:	val_out <= 4'ha71f;
         4'hcb0 	:	val_out <= 4'ha737;
         4'hcb1 	:	val_out <= 4'ha737;
         4'hcb2 	:	val_out <= 4'ha737;
         4'hcb3 	:	val_out <= 4'ha737;
         4'hcb8 	:	val_out <= 4'ha74f;
         4'hcb9 	:	val_out <= 4'ha74f;
         4'hcba 	:	val_out <= 4'ha74f;
         4'hcbb 	:	val_out <= 4'ha74f;
         4'hcc0 	:	val_out <= 4'ha767;
         4'hcc1 	:	val_out <= 4'ha767;
         4'hcc2 	:	val_out <= 4'ha767;
         4'hcc3 	:	val_out <= 4'ha767;
         4'hcc8 	:	val_out <= 4'ha77f;
         4'hcc9 	:	val_out <= 4'ha77f;
         4'hcca 	:	val_out <= 4'ha77f;
         4'hccb 	:	val_out <= 4'ha77f;
         4'hcd0 	:	val_out <= 4'ha797;
         4'hcd1 	:	val_out <= 4'ha797;
         4'hcd2 	:	val_out <= 4'ha797;
         4'hcd3 	:	val_out <= 4'ha797;
         4'hcd8 	:	val_out <= 4'ha7af;
         4'hcd9 	:	val_out <= 4'ha7af;
         4'hcda 	:	val_out <= 4'ha7af;
         4'hcdb 	:	val_out <= 4'ha7af;
         4'hce0 	:	val_out <= 4'ha7c7;
         4'hce1 	:	val_out <= 4'ha7c7;
         4'hce2 	:	val_out <= 4'ha7c7;
         4'hce3 	:	val_out <= 4'ha7c7;
         4'hce8 	:	val_out <= 4'ha7df;
         4'hce9 	:	val_out <= 4'ha7df;
         4'hcea 	:	val_out <= 4'ha7df;
         4'hceb 	:	val_out <= 4'ha7df;
         4'hcf0 	:	val_out <= 4'ha7f6;
         4'hcf1 	:	val_out <= 4'ha7f6;
         4'hcf2 	:	val_out <= 4'ha7f6;
         4'hcf3 	:	val_out <= 4'ha7f6;
         4'hcf8 	:	val_out <= 4'ha80e;
         4'hcf9 	:	val_out <= 4'ha80e;
         4'hcfa 	:	val_out <= 4'ha80e;
         4'hcfb 	:	val_out <= 4'ha80e;
         4'hd00 	:	val_out <= 4'ha826;
         4'hd01 	:	val_out <= 4'ha826;
         4'hd02 	:	val_out <= 4'ha826;
         4'hd03 	:	val_out <= 4'ha826;
         4'hd08 	:	val_out <= 4'ha83e;
         4'hd09 	:	val_out <= 4'ha83e;
         4'hd0a 	:	val_out <= 4'ha83e;
         4'hd0b 	:	val_out <= 4'ha83e;
         4'hd10 	:	val_out <= 4'ha856;
         4'hd11 	:	val_out <= 4'ha856;
         4'hd12 	:	val_out <= 4'ha856;
         4'hd13 	:	val_out <= 4'ha856;
         4'hd18 	:	val_out <= 4'ha86e;
         4'hd19 	:	val_out <= 4'ha86e;
         4'hd1a 	:	val_out <= 4'ha86e;
         4'hd1b 	:	val_out <= 4'ha86e;
         4'hd20 	:	val_out <= 4'ha886;
         4'hd21 	:	val_out <= 4'ha886;
         4'hd22 	:	val_out <= 4'ha886;
         4'hd23 	:	val_out <= 4'ha886;
         4'hd28 	:	val_out <= 4'ha89d;
         4'hd29 	:	val_out <= 4'ha89d;
         4'hd2a 	:	val_out <= 4'ha89d;
         4'hd2b 	:	val_out <= 4'ha89d;
         4'hd30 	:	val_out <= 4'ha8b5;
         4'hd31 	:	val_out <= 4'ha8b5;
         4'hd32 	:	val_out <= 4'ha8b5;
         4'hd33 	:	val_out <= 4'ha8b5;
         4'hd38 	:	val_out <= 4'ha8cd;
         4'hd39 	:	val_out <= 4'ha8cd;
         4'hd3a 	:	val_out <= 4'ha8cd;
         4'hd3b 	:	val_out <= 4'ha8cd;
         4'hd40 	:	val_out <= 4'ha8e5;
         4'hd41 	:	val_out <= 4'ha8e5;
         4'hd42 	:	val_out <= 4'ha8e5;
         4'hd43 	:	val_out <= 4'ha8e5;
         4'hd48 	:	val_out <= 4'ha8fd;
         4'hd49 	:	val_out <= 4'ha8fd;
         4'hd4a 	:	val_out <= 4'ha8fd;
         4'hd4b 	:	val_out <= 4'ha8fd;
         4'hd50 	:	val_out <= 4'ha915;
         4'hd51 	:	val_out <= 4'ha915;
         4'hd52 	:	val_out <= 4'ha915;
         4'hd53 	:	val_out <= 4'ha915;
         4'hd58 	:	val_out <= 4'ha92c;
         4'hd59 	:	val_out <= 4'ha92c;
         4'hd5a 	:	val_out <= 4'ha92c;
         4'hd5b 	:	val_out <= 4'ha92c;
         4'hd60 	:	val_out <= 4'ha944;
         4'hd61 	:	val_out <= 4'ha944;
         4'hd62 	:	val_out <= 4'ha944;
         4'hd63 	:	val_out <= 4'ha944;
         4'hd68 	:	val_out <= 4'ha95c;
         4'hd69 	:	val_out <= 4'ha95c;
         4'hd6a 	:	val_out <= 4'ha95c;
         4'hd6b 	:	val_out <= 4'ha95c;
         4'hd70 	:	val_out <= 4'ha974;
         4'hd71 	:	val_out <= 4'ha974;
         4'hd72 	:	val_out <= 4'ha974;
         4'hd73 	:	val_out <= 4'ha974;
         4'hd78 	:	val_out <= 4'ha98b;
         4'hd79 	:	val_out <= 4'ha98b;
         4'hd7a 	:	val_out <= 4'ha98b;
         4'hd7b 	:	val_out <= 4'ha98b;
         4'hd80 	:	val_out <= 4'ha9a3;
         4'hd81 	:	val_out <= 4'ha9a3;
         4'hd82 	:	val_out <= 4'ha9a3;
         4'hd83 	:	val_out <= 4'ha9a3;
         4'hd88 	:	val_out <= 4'ha9bb;
         4'hd89 	:	val_out <= 4'ha9bb;
         4'hd8a 	:	val_out <= 4'ha9bb;
         4'hd8b 	:	val_out <= 4'ha9bb;
         4'hd90 	:	val_out <= 4'ha9d3;
         4'hd91 	:	val_out <= 4'ha9d3;
         4'hd92 	:	val_out <= 4'ha9d3;
         4'hd93 	:	val_out <= 4'ha9d3;
         4'hd98 	:	val_out <= 4'ha9eb;
         4'hd99 	:	val_out <= 4'ha9eb;
         4'hd9a 	:	val_out <= 4'ha9eb;
         4'hd9b 	:	val_out <= 4'ha9eb;
         4'hda0 	:	val_out <= 4'haa02;
         4'hda1 	:	val_out <= 4'haa02;
         4'hda2 	:	val_out <= 4'haa02;
         4'hda3 	:	val_out <= 4'haa02;
         4'hda8 	:	val_out <= 4'haa1a;
         4'hda9 	:	val_out <= 4'haa1a;
         4'hdaa 	:	val_out <= 4'haa1a;
         4'hdab 	:	val_out <= 4'haa1a;
         4'hdb0 	:	val_out <= 4'haa32;
         4'hdb1 	:	val_out <= 4'haa32;
         4'hdb2 	:	val_out <= 4'haa32;
         4'hdb3 	:	val_out <= 4'haa32;
         4'hdb8 	:	val_out <= 4'haa49;
         4'hdb9 	:	val_out <= 4'haa49;
         4'hdba 	:	val_out <= 4'haa49;
         4'hdbb 	:	val_out <= 4'haa49;
         4'hdc0 	:	val_out <= 4'haa61;
         4'hdc1 	:	val_out <= 4'haa61;
         4'hdc2 	:	val_out <= 4'haa61;
         4'hdc3 	:	val_out <= 4'haa61;
         4'hdc8 	:	val_out <= 4'haa79;
         4'hdc9 	:	val_out <= 4'haa79;
         4'hdca 	:	val_out <= 4'haa79;
         4'hdcb 	:	val_out <= 4'haa79;
         4'hdd0 	:	val_out <= 4'haa91;
         4'hdd1 	:	val_out <= 4'haa91;
         4'hdd2 	:	val_out <= 4'haa91;
         4'hdd3 	:	val_out <= 4'haa91;
         4'hdd8 	:	val_out <= 4'haaa8;
         4'hdd9 	:	val_out <= 4'haaa8;
         4'hdda 	:	val_out <= 4'haaa8;
         4'hddb 	:	val_out <= 4'haaa8;
         4'hde0 	:	val_out <= 4'haac0;
         4'hde1 	:	val_out <= 4'haac0;
         4'hde2 	:	val_out <= 4'haac0;
         4'hde3 	:	val_out <= 4'haac0;
         4'hde8 	:	val_out <= 4'haad8;
         4'hde9 	:	val_out <= 4'haad8;
         4'hdea 	:	val_out <= 4'haad8;
         4'hdeb 	:	val_out <= 4'haad8;
         4'hdf0 	:	val_out <= 4'haaef;
         4'hdf1 	:	val_out <= 4'haaef;
         4'hdf2 	:	val_out <= 4'haaef;
         4'hdf3 	:	val_out <= 4'haaef;
         4'hdf8 	:	val_out <= 4'hab07;
         4'hdf9 	:	val_out <= 4'hab07;
         4'hdfa 	:	val_out <= 4'hab07;
         4'hdfb 	:	val_out <= 4'hab07;
         4'he00 	:	val_out <= 4'hab1f;
         4'he01 	:	val_out <= 4'hab1f;
         4'he02 	:	val_out <= 4'hab1f;
         4'he03 	:	val_out <= 4'hab1f;
         4'he08 	:	val_out <= 4'hab36;
         4'he09 	:	val_out <= 4'hab36;
         4'he0a 	:	val_out <= 4'hab36;
         4'he0b 	:	val_out <= 4'hab36;
         4'he10 	:	val_out <= 4'hab4e;
         4'he11 	:	val_out <= 4'hab4e;
         4'he12 	:	val_out <= 4'hab4e;
         4'he13 	:	val_out <= 4'hab4e;
         4'he18 	:	val_out <= 4'hab66;
         4'he19 	:	val_out <= 4'hab66;
         4'he1a 	:	val_out <= 4'hab66;
         4'he1b 	:	val_out <= 4'hab66;
         4'he20 	:	val_out <= 4'hab7d;
         4'he21 	:	val_out <= 4'hab7d;
         4'he22 	:	val_out <= 4'hab7d;
         4'he23 	:	val_out <= 4'hab7d;
         4'he28 	:	val_out <= 4'hab95;
         4'he29 	:	val_out <= 4'hab95;
         4'he2a 	:	val_out <= 4'hab95;
         4'he2b 	:	val_out <= 4'hab95;
         4'he30 	:	val_out <= 4'habad;
         4'he31 	:	val_out <= 4'habad;
         4'he32 	:	val_out <= 4'habad;
         4'he33 	:	val_out <= 4'habad;
         4'he38 	:	val_out <= 4'habc4;
         4'he39 	:	val_out <= 4'habc4;
         4'he3a 	:	val_out <= 4'habc4;
         4'he3b 	:	val_out <= 4'habc4;
         4'he40 	:	val_out <= 4'habdc;
         4'he41 	:	val_out <= 4'habdc;
         4'he42 	:	val_out <= 4'habdc;
         4'he43 	:	val_out <= 4'habdc;
         4'he48 	:	val_out <= 4'habf3;
         4'he49 	:	val_out <= 4'habf3;
         4'he4a 	:	val_out <= 4'habf3;
         4'he4b 	:	val_out <= 4'habf3;
         4'he50 	:	val_out <= 4'hac0b;
         4'he51 	:	val_out <= 4'hac0b;
         4'he52 	:	val_out <= 4'hac0b;
         4'he53 	:	val_out <= 4'hac0b;
         4'he58 	:	val_out <= 4'hac23;
         4'he59 	:	val_out <= 4'hac23;
         4'he5a 	:	val_out <= 4'hac23;
         4'he5b 	:	val_out <= 4'hac23;
         4'he60 	:	val_out <= 4'hac3a;
         4'he61 	:	val_out <= 4'hac3a;
         4'he62 	:	val_out <= 4'hac3a;
         4'he63 	:	val_out <= 4'hac3a;
         4'he68 	:	val_out <= 4'hac52;
         4'he69 	:	val_out <= 4'hac52;
         4'he6a 	:	val_out <= 4'hac52;
         4'he6b 	:	val_out <= 4'hac52;
         4'he70 	:	val_out <= 4'hac69;
         4'he71 	:	val_out <= 4'hac69;
         4'he72 	:	val_out <= 4'hac69;
         4'he73 	:	val_out <= 4'hac69;
         4'he78 	:	val_out <= 4'hac81;
         4'he79 	:	val_out <= 4'hac81;
         4'he7a 	:	val_out <= 4'hac81;
         4'he7b 	:	val_out <= 4'hac81;
         4'he80 	:	val_out <= 4'hac98;
         4'he81 	:	val_out <= 4'hac98;
         4'he82 	:	val_out <= 4'hac98;
         4'he83 	:	val_out <= 4'hac98;
         4'he88 	:	val_out <= 4'hacb0;
         4'he89 	:	val_out <= 4'hacb0;
         4'he8a 	:	val_out <= 4'hacb0;
         4'he8b 	:	val_out <= 4'hacb0;
         4'he90 	:	val_out <= 4'hacc8;
         4'he91 	:	val_out <= 4'hacc8;
         4'he92 	:	val_out <= 4'hacc8;
         4'he93 	:	val_out <= 4'hacc8;
         4'he98 	:	val_out <= 4'hacdf;
         4'he99 	:	val_out <= 4'hacdf;
         4'he9a 	:	val_out <= 4'hacdf;
         4'he9b 	:	val_out <= 4'hacdf;
         4'hea0 	:	val_out <= 4'hacf7;
         4'hea1 	:	val_out <= 4'hacf7;
         4'hea2 	:	val_out <= 4'hacf7;
         4'hea3 	:	val_out <= 4'hacf7;
         4'hea8 	:	val_out <= 4'had0e;
         4'hea9 	:	val_out <= 4'had0e;
         4'heaa 	:	val_out <= 4'had0e;
         4'heab 	:	val_out <= 4'had0e;
         4'heb0 	:	val_out <= 4'had26;
         4'heb1 	:	val_out <= 4'had26;
         4'heb2 	:	val_out <= 4'had26;
         4'heb3 	:	val_out <= 4'had26;
         4'heb8 	:	val_out <= 4'had3d;
         4'heb9 	:	val_out <= 4'had3d;
         4'heba 	:	val_out <= 4'had3d;
         4'hebb 	:	val_out <= 4'had3d;
         4'hec0 	:	val_out <= 4'had55;
         4'hec1 	:	val_out <= 4'had55;
         4'hec2 	:	val_out <= 4'had55;
         4'hec3 	:	val_out <= 4'had55;
         4'hec8 	:	val_out <= 4'had6c;
         4'hec9 	:	val_out <= 4'had6c;
         4'heca 	:	val_out <= 4'had6c;
         4'hecb 	:	val_out <= 4'had6c;
         4'hed0 	:	val_out <= 4'had84;
         4'hed1 	:	val_out <= 4'had84;
         4'hed2 	:	val_out <= 4'had84;
         4'hed3 	:	val_out <= 4'had84;
         4'hed8 	:	val_out <= 4'had9b;
         4'hed9 	:	val_out <= 4'had9b;
         4'heda 	:	val_out <= 4'had9b;
         4'hedb 	:	val_out <= 4'had9b;
         4'hee0 	:	val_out <= 4'hadb3;
         4'hee1 	:	val_out <= 4'hadb3;
         4'hee2 	:	val_out <= 4'hadb3;
         4'hee3 	:	val_out <= 4'hadb3;
         4'hee8 	:	val_out <= 4'hadca;
         4'hee9 	:	val_out <= 4'hadca;
         4'heea 	:	val_out <= 4'hadca;
         4'heeb 	:	val_out <= 4'hadca;
         4'hef0 	:	val_out <= 4'hade2;
         4'hef1 	:	val_out <= 4'hade2;
         4'hef2 	:	val_out <= 4'hade2;
         4'hef3 	:	val_out <= 4'hade2;
         4'hef8 	:	val_out <= 4'hadf9;
         4'hef9 	:	val_out <= 4'hadf9;
         4'hefa 	:	val_out <= 4'hadf9;
         4'hefb 	:	val_out <= 4'hadf9;
         4'hf00 	:	val_out <= 4'hae11;
         4'hf01 	:	val_out <= 4'hae11;
         4'hf02 	:	val_out <= 4'hae11;
         4'hf03 	:	val_out <= 4'hae11;
         4'hf08 	:	val_out <= 4'hae28;
         4'hf09 	:	val_out <= 4'hae28;
         4'hf0a 	:	val_out <= 4'hae28;
         4'hf0b 	:	val_out <= 4'hae28;
         4'hf10 	:	val_out <= 4'hae3f;
         4'hf11 	:	val_out <= 4'hae3f;
         4'hf12 	:	val_out <= 4'hae3f;
         4'hf13 	:	val_out <= 4'hae3f;
         4'hf18 	:	val_out <= 4'hae57;
         4'hf19 	:	val_out <= 4'hae57;
         4'hf1a 	:	val_out <= 4'hae57;
         4'hf1b 	:	val_out <= 4'hae57;
         4'hf20 	:	val_out <= 4'hae6e;
         4'hf21 	:	val_out <= 4'hae6e;
         4'hf22 	:	val_out <= 4'hae6e;
         4'hf23 	:	val_out <= 4'hae6e;
         4'hf28 	:	val_out <= 4'hae86;
         4'hf29 	:	val_out <= 4'hae86;
         4'hf2a 	:	val_out <= 4'hae86;
         4'hf2b 	:	val_out <= 4'hae86;
         4'hf30 	:	val_out <= 4'hae9d;
         4'hf31 	:	val_out <= 4'hae9d;
         4'hf32 	:	val_out <= 4'hae9d;
         4'hf33 	:	val_out <= 4'hae9d;
         4'hf38 	:	val_out <= 4'haeb5;
         4'hf39 	:	val_out <= 4'haeb5;
         4'hf3a 	:	val_out <= 4'haeb5;
         4'hf3b 	:	val_out <= 4'haeb5;
         4'hf40 	:	val_out <= 4'haecc;
         4'hf41 	:	val_out <= 4'haecc;
         4'hf42 	:	val_out <= 4'haecc;
         4'hf43 	:	val_out <= 4'haecc;
         4'hf48 	:	val_out <= 4'haee3;
         4'hf49 	:	val_out <= 4'haee3;
         4'hf4a 	:	val_out <= 4'haee3;
         4'hf4b 	:	val_out <= 4'haee3;
         4'hf50 	:	val_out <= 4'haefb;
         4'hf51 	:	val_out <= 4'haefb;
         4'hf52 	:	val_out <= 4'haefb;
         4'hf53 	:	val_out <= 4'haefb;
         4'hf58 	:	val_out <= 4'haf12;
         4'hf59 	:	val_out <= 4'haf12;
         4'hf5a 	:	val_out <= 4'haf12;
         4'hf5b 	:	val_out <= 4'haf12;
         4'hf60 	:	val_out <= 4'haf29;
         4'hf61 	:	val_out <= 4'haf29;
         4'hf62 	:	val_out <= 4'haf29;
         4'hf63 	:	val_out <= 4'haf29;
         4'hf68 	:	val_out <= 4'haf41;
         4'hf69 	:	val_out <= 4'haf41;
         4'hf6a 	:	val_out <= 4'haf41;
         4'hf6b 	:	val_out <= 4'haf41;
         4'hf70 	:	val_out <= 4'haf58;
         4'hf71 	:	val_out <= 4'haf58;
         4'hf72 	:	val_out <= 4'haf58;
         4'hf73 	:	val_out <= 4'haf58;
         4'hf78 	:	val_out <= 4'haf6f;
         4'hf79 	:	val_out <= 4'haf6f;
         4'hf7a 	:	val_out <= 4'haf6f;
         4'hf7b 	:	val_out <= 4'haf6f;
         4'hf80 	:	val_out <= 4'haf87;
         4'hf81 	:	val_out <= 4'haf87;
         4'hf82 	:	val_out <= 4'haf87;
         4'hf83 	:	val_out <= 4'haf87;
         4'hf88 	:	val_out <= 4'haf9e;
         4'hf89 	:	val_out <= 4'haf9e;
         4'hf8a 	:	val_out <= 4'haf9e;
         4'hf8b 	:	val_out <= 4'haf9e;
         4'hf90 	:	val_out <= 4'hafb5;
         4'hf91 	:	val_out <= 4'hafb5;
         4'hf92 	:	val_out <= 4'hafb5;
         4'hf93 	:	val_out <= 4'hafb5;
         4'hf98 	:	val_out <= 4'hafcd;
         4'hf99 	:	val_out <= 4'hafcd;
         4'hf9a 	:	val_out <= 4'hafcd;
         4'hf9b 	:	val_out <= 4'hafcd;
         4'hfa0 	:	val_out <= 4'hafe4;
         4'hfa1 	:	val_out <= 4'hafe4;
         4'hfa2 	:	val_out <= 4'hafe4;
         4'hfa3 	:	val_out <= 4'hafe4;
         4'hfa8 	:	val_out <= 4'haffb;
         4'hfa9 	:	val_out <= 4'haffb;
         4'hfaa 	:	val_out <= 4'haffb;
         4'hfab 	:	val_out <= 4'haffb;
         4'hfb0 	:	val_out <= 4'hb013;
         4'hfb1 	:	val_out <= 4'hb013;
         4'hfb2 	:	val_out <= 4'hb013;
         4'hfb3 	:	val_out <= 4'hb013;
         4'hfb8 	:	val_out <= 4'hb02a;
         4'hfb9 	:	val_out <= 4'hb02a;
         4'hfba 	:	val_out <= 4'hb02a;
         4'hfbb 	:	val_out <= 4'hb02a;
         4'hfc0 	:	val_out <= 4'hb041;
         4'hfc1 	:	val_out <= 4'hb041;
         4'hfc2 	:	val_out <= 4'hb041;
         4'hfc3 	:	val_out <= 4'hb041;
         4'hfc8 	:	val_out <= 4'hb059;
         4'hfc9 	:	val_out <= 4'hb059;
         4'hfca 	:	val_out <= 4'hb059;
         4'hfcb 	:	val_out <= 4'hb059;
         4'hfd0 	:	val_out <= 4'hb070;
         4'hfd1 	:	val_out <= 4'hb070;
         4'hfd2 	:	val_out <= 4'hb070;
         4'hfd3 	:	val_out <= 4'hb070;
         4'hfd8 	:	val_out <= 4'hb087;
         4'hfd9 	:	val_out <= 4'hb087;
         4'hfda 	:	val_out <= 4'hb087;
         4'hfdb 	:	val_out <= 4'hb087;
         4'hfe0 	:	val_out <= 4'hb09e;
         4'hfe1 	:	val_out <= 4'hb09e;
         4'hfe2 	:	val_out <= 4'hb09e;
         4'hfe3 	:	val_out <= 4'hb09e;
         4'hfe8 	:	val_out <= 4'hb0b6;
         4'hfe9 	:	val_out <= 4'hb0b6;
         4'hfea 	:	val_out <= 4'hb0b6;
         4'hfeb 	:	val_out <= 4'hb0b6;
         4'hff0 	:	val_out <= 4'hb0cd;
         4'hff1 	:	val_out <= 4'hb0cd;
         4'hff2 	:	val_out <= 4'hb0cd;
         4'hff3 	:	val_out <= 4'hb0cd;
         4'hff8 	:	val_out <= 4'hb0e4;
         4'hff9 	:	val_out <= 4'hb0e4;
         4'hffa 	:	val_out <= 4'hb0e4;
         4'hffb 	:	val_out <= 4'hb0e4;
         4'h1000 	:	val_out <= 4'hb0fb;
         4'h1001 	:	val_out <= 4'hb0fb;
         4'h1002 	:	val_out <= 4'hb0fb;
         4'h1003 	:	val_out <= 4'hb0fb;
         4'h1008 	:	val_out <= 4'hb112;
         4'h1009 	:	val_out <= 4'hb112;
         4'h100a 	:	val_out <= 4'hb112;
         4'h100b 	:	val_out <= 4'hb112;
         4'h1010 	:	val_out <= 4'hb12a;
         4'h1011 	:	val_out <= 4'hb12a;
         4'h1012 	:	val_out <= 4'hb12a;
         4'h1013 	:	val_out <= 4'hb12a;
         4'h1018 	:	val_out <= 4'hb141;
         4'h1019 	:	val_out <= 4'hb141;
         4'h101a 	:	val_out <= 4'hb141;
         4'h101b 	:	val_out <= 4'hb141;
         4'h1020 	:	val_out <= 4'hb158;
         4'h1021 	:	val_out <= 4'hb158;
         4'h1022 	:	val_out <= 4'hb158;
         4'h1023 	:	val_out <= 4'hb158;
         4'h1028 	:	val_out <= 4'hb16f;
         4'h1029 	:	val_out <= 4'hb16f;
         4'h102a 	:	val_out <= 4'hb16f;
         4'h102b 	:	val_out <= 4'hb16f;
         4'h1030 	:	val_out <= 4'hb186;
         4'h1031 	:	val_out <= 4'hb186;
         4'h1032 	:	val_out <= 4'hb186;
         4'h1033 	:	val_out <= 4'hb186;
         4'h1038 	:	val_out <= 4'hb19e;
         4'h1039 	:	val_out <= 4'hb19e;
         4'h103a 	:	val_out <= 4'hb19e;
         4'h103b 	:	val_out <= 4'hb19e;
         4'h1040 	:	val_out <= 4'hb1b5;
         4'h1041 	:	val_out <= 4'hb1b5;
         4'h1042 	:	val_out <= 4'hb1b5;
         4'h1043 	:	val_out <= 4'hb1b5;
         4'h1048 	:	val_out <= 4'hb1cc;
         4'h1049 	:	val_out <= 4'hb1cc;
         4'h104a 	:	val_out <= 4'hb1cc;
         4'h104b 	:	val_out <= 4'hb1cc;
         4'h1050 	:	val_out <= 4'hb1e3;
         4'h1051 	:	val_out <= 4'hb1e3;
         4'h1052 	:	val_out <= 4'hb1e3;
         4'h1053 	:	val_out <= 4'hb1e3;
         4'h1058 	:	val_out <= 4'hb1fa;
         4'h1059 	:	val_out <= 4'hb1fa;
         4'h105a 	:	val_out <= 4'hb1fa;
         4'h105b 	:	val_out <= 4'hb1fa;
         4'h1060 	:	val_out <= 4'hb211;
         4'h1061 	:	val_out <= 4'hb211;
         4'h1062 	:	val_out <= 4'hb211;
         4'h1063 	:	val_out <= 4'hb211;
         4'h1068 	:	val_out <= 4'hb228;
         4'h1069 	:	val_out <= 4'hb228;
         4'h106a 	:	val_out <= 4'hb228;
         4'h106b 	:	val_out <= 4'hb228;
         4'h1070 	:	val_out <= 4'hb240;
         4'h1071 	:	val_out <= 4'hb240;
         4'h1072 	:	val_out <= 4'hb240;
         4'h1073 	:	val_out <= 4'hb240;
         4'h1078 	:	val_out <= 4'hb257;
         4'h1079 	:	val_out <= 4'hb257;
         4'h107a 	:	val_out <= 4'hb257;
         4'h107b 	:	val_out <= 4'hb257;
         4'h1080 	:	val_out <= 4'hb26e;
         4'h1081 	:	val_out <= 4'hb26e;
         4'h1082 	:	val_out <= 4'hb26e;
         4'h1083 	:	val_out <= 4'hb26e;
         4'h1088 	:	val_out <= 4'hb285;
         4'h1089 	:	val_out <= 4'hb285;
         4'h108a 	:	val_out <= 4'hb285;
         4'h108b 	:	val_out <= 4'hb285;
         4'h1090 	:	val_out <= 4'hb29c;
         4'h1091 	:	val_out <= 4'hb29c;
         4'h1092 	:	val_out <= 4'hb29c;
         4'h1093 	:	val_out <= 4'hb29c;
         4'h1098 	:	val_out <= 4'hb2b3;
         4'h1099 	:	val_out <= 4'hb2b3;
         4'h109a 	:	val_out <= 4'hb2b3;
         4'h109b 	:	val_out <= 4'hb2b3;
         4'h10a0 	:	val_out <= 4'hb2ca;
         4'h10a1 	:	val_out <= 4'hb2ca;
         4'h10a2 	:	val_out <= 4'hb2ca;
         4'h10a3 	:	val_out <= 4'hb2ca;
         4'h10a8 	:	val_out <= 4'hb2e1;
         4'h10a9 	:	val_out <= 4'hb2e1;
         4'h10aa 	:	val_out <= 4'hb2e1;
         4'h10ab 	:	val_out <= 4'hb2e1;
         4'h10b0 	:	val_out <= 4'hb2f8;
         4'h10b1 	:	val_out <= 4'hb2f8;
         4'h10b2 	:	val_out <= 4'hb2f8;
         4'h10b3 	:	val_out <= 4'hb2f8;
         4'h10b8 	:	val_out <= 4'hb30f;
         4'h10b9 	:	val_out <= 4'hb30f;
         4'h10ba 	:	val_out <= 4'hb30f;
         4'h10bb 	:	val_out <= 4'hb30f;
         4'h10c0 	:	val_out <= 4'hb326;
         4'h10c1 	:	val_out <= 4'hb326;
         4'h10c2 	:	val_out <= 4'hb326;
         4'h10c3 	:	val_out <= 4'hb326;
         4'h10c8 	:	val_out <= 4'hb33d;
         4'h10c9 	:	val_out <= 4'hb33d;
         4'h10ca 	:	val_out <= 4'hb33d;
         4'h10cb 	:	val_out <= 4'hb33d;
         4'h10d0 	:	val_out <= 4'hb354;
         4'h10d1 	:	val_out <= 4'hb354;
         4'h10d2 	:	val_out <= 4'hb354;
         4'h10d3 	:	val_out <= 4'hb354;
         4'h10d8 	:	val_out <= 4'hb36b;
         4'h10d9 	:	val_out <= 4'hb36b;
         4'h10da 	:	val_out <= 4'hb36b;
         4'h10db 	:	val_out <= 4'hb36b;
         4'h10e0 	:	val_out <= 4'hb382;
         4'h10e1 	:	val_out <= 4'hb382;
         4'h10e2 	:	val_out <= 4'hb382;
         4'h10e3 	:	val_out <= 4'hb382;
         4'h10e8 	:	val_out <= 4'hb399;
         4'h10e9 	:	val_out <= 4'hb399;
         4'h10ea 	:	val_out <= 4'hb399;
         4'h10eb 	:	val_out <= 4'hb399;
         4'h10f0 	:	val_out <= 4'hb3b0;
         4'h10f1 	:	val_out <= 4'hb3b0;
         4'h10f2 	:	val_out <= 4'hb3b0;
         4'h10f3 	:	val_out <= 4'hb3b0;
         4'h10f8 	:	val_out <= 4'hb3c7;
         4'h10f9 	:	val_out <= 4'hb3c7;
         4'h10fa 	:	val_out <= 4'hb3c7;
         4'h10fb 	:	val_out <= 4'hb3c7;
         4'h1100 	:	val_out <= 4'hb3de;
         4'h1101 	:	val_out <= 4'hb3de;
         4'h1102 	:	val_out <= 4'hb3de;
         4'h1103 	:	val_out <= 4'hb3de;
         4'h1108 	:	val_out <= 4'hb3f5;
         4'h1109 	:	val_out <= 4'hb3f5;
         4'h110a 	:	val_out <= 4'hb3f5;
         4'h110b 	:	val_out <= 4'hb3f5;
         4'h1110 	:	val_out <= 4'hb40c;
         4'h1111 	:	val_out <= 4'hb40c;
         4'h1112 	:	val_out <= 4'hb40c;
         4'h1113 	:	val_out <= 4'hb40c;
         4'h1118 	:	val_out <= 4'hb423;
         4'h1119 	:	val_out <= 4'hb423;
         4'h111a 	:	val_out <= 4'hb423;
         4'h111b 	:	val_out <= 4'hb423;
         4'h1120 	:	val_out <= 4'hb43a;
         4'h1121 	:	val_out <= 4'hb43a;
         4'h1122 	:	val_out <= 4'hb43a;
         4'h1123 	:	val_out <= 4'hb43a;
         4'h1128 	:	val_out <= 4'hb451;
         4'h1129 	:	val_out <= 4'hb451;
         4'h112a 	:	val_out <= 4'hb451;
         4'h112b 	:	val_out <= 4'hb451;
         4'h1130 	:	val_out <= 4'hb468;
         4'h1131 	:	val_out <= 4'hb468;
         4'h1132 	:	val_out <= 4'hb468;
         4'h1133 	:	val_out <= 4'hb468;
         4'h1138 	:	val_out <= 4'hb47f;
         4'h1139 	:	val_out <= 4'hb47f;
         4'h113a 	:	val_out <= 4'hb47f;
         4'h113b 	:	val_out <= 4'hb47f;
         4'h1140 	:	val_out <= 4'hb496;
         4'h1141 	:	val_out <= 4'hb496;
         4'h1142 	:	val_out <= 4'hb496;
         4'h1143 	:	val_out <= 4'hb496;
         4'h1148 	:	val_out <= 4'hb4ad;
         4'h1149 	:	val_out <= 4'hb4ad;
         4'h114a 	:	val_out <= 4'hb4ad;
         4'h114b 	:	val_out <= 4'hb4ad;
         4'h1150 	:	val_out <= 4'hb4c4;
         4'h1151 	:	val_out <= 4'hb4c4;
         4'h1152 	:	val_out <= 4'hb4c4;
         4'h1153 	:	val_out <= 4'hb4c4;
         4'h1158 	:	val_out <= 4'hb4db;
         4'h1159 	:	val_out <= 4'hb4db;
         4'h115a 	:	val_out <= 4'hb4db;
         4'h115b 	:	val_out <= 4'hb4db;
         4'h1160 	:	val_out <= 4'hb4f2;
         4'h1161 	:	val_out <= 4'hb4f2;
         4'h1162 	:	val_out <= 4'hb4f2;
         4'h1163 	:	val_out <= 4'hb4f2;
         4'h1168 	:	val_out <= 4'hb508;
         4'h1169 	:	val_out <= 4'hb508;
         4'h116a 	:	val_out <= 4'hb508;
         4'h116b 	:	val_out <= 4'hb508;
         4'h1170 	:	val_out <= 4'hb51f;
         4'h1171 	:	val_out <= 4'hb51f;
         4'h1172 	:	val_out <= 4'hb51f;
         4'h1173 	:	val_out <= 4'hb51f;
         4'h1178 	:	val_out <= 4'hb536;
         4'h1179 	:	val_out <= 4'hb536;
         4'h117a 	:	val_out <= 4'hb536;
         4'h117b 	:	val_out <= 4'hb536;
         4'h1180 	:	val_out <= 4'hb54d;
         4'h1181 	:	val_out <= 4'hb54d;
         4'h1182 	:	val_out <= 4'hb54d;
         4'h1183 	:	val_out <= 4'hb54d;
         4'h1188 	:	val_out <= 4'hb564;
         4'h1189 	:	val_out <= 4'hb564;
         4'h118a 	:	val_out <= 4'hb564;
         4'h118b 	:	val_out <= 4'hb564;
         4'h1190 	:	val_out <= 4'hb57b;
         4'h1191 	:	val_out <= 4'hb57b;
         4'h1192 	:	val_out <= 4'hb57b;
         4'h1193 	:	val_out <= 4'hb57b;
         4'h1198 	:	val_out <= 4'hb592;
         4'h1199 	:	val_out <= 4'hb592;
         4'h119a 	:	val_out <= 4'hb592;
         4'h119b 	:	val_out <= 4'hb592;
         4'h11a0 	:	val_out <= 4'hb5a8;
         4'h11a1 	:	val_out <= 4'hb5a8;
         4'h11a2 	:	val_out <= 4'hb5a8;
         4'h11a3 	:	val_out <= 4'hb5a8;
         4'h11a8 	:	val_out <= 4'hb5bf;
         4'h11a9 	:	val_out <= 4'hb5bf;
         4'h11aa 	:	val_out <= 4'hb5bf;
         4'h11ab 	:	val_out <= 4'hb5bf;
         4'h11b0 	:	val_out <= 4'hb5d6;
         4'h11b1 	:	val_out <= 4'hb5d6;
         4'h11b2 	:	val_out <= 4'hb5d6;
         4'h11b3 	:	val_out <= 4'hb5d6;
         4'h11b8 	:	val_out <= 4'hb5ed;
         4'h11b9 	:	val_out <= 4'hb5ed;
         4'h11ba 	:	val_out <= 4'hb5ed;
         4'h11bb 	:	val_out <= 4'hb5ed;
         4'h11c0 	:	val_out <= 4'hb604;
         4'h11c1 	:	val_out <= 4'hb604;
         4'h11c2 	:	val_out <= 4'hb604;
         4'h11c3 	:	val_out <= 4'hb604;
         4'h11c8 	:	val_out <= 4'hb61a;
         4'h11c9 	:	val_out <= 4'hb61a;
         4'h11ca 	:	val_out <= 4'hb61a;
         4'h11cb 	:	val_out <= 4'hb61a;
         4'h11d0 	:	val_out <= 4'hb631;
         4'h11d1 	:	val_out <= 4'hb631;
         4'h11d2 	:	val_out <= 4'hb631;
         4'h11d3 	:	val_out <= 4'hb631;
         4'h11d8 	:	val_out <= 4'hb648;
         4'h11d9 	:	val_out <= 4'hb648;
         4'h11da 	:	val_out <= 4'hb648;
         4'h11db 	:	val_out <= 4'hb648;
         4'h11e0 	:	val_out <= 4'hb65f;
         4'h11e1 	:	val_out <= 4'hb65f;
         4'h11e2 	:	val_out <= 4'hb65f;
         4'h11e3 	:	val_out <= 4'hb65f;
         4'h11e8 	:	val_out <= 4'hb675;
         4'h11e9 	:	val_out <= 4'hb675;
         4'h11ea 	:	val_out <= 4'hb675;
         4'h11eb 	:	val_out <= 4'hb675;
         4'h11f0 	:	val_out <= 4'hb68c;
         4'h11f1 	:	val_out <= 4'hb68c;
         4'h11f2 	:	val_out <= 4'hb68c;
         4'h11f3 	:	val_out <= 4'hb68c;
         4'h11f8 	:	val_out <= 4'hb6a3;
         4'h11f9 	:	val_out <= 4'hb6a3;
         4'h11fa 	:	val_out <= 4'hb6a3;
         4'h11fb 	:	val_out <= 4'hb6a3;
         4'h1200 	:	val_out <= 4'hb6ba;
         4'h1201 	:	val_out <= 4'hb6ba;
         4'h1202 	:	val_out <= 4'hb6ba;
         4'h1203 	:	val_out <= 4'hb6ba;
         4'h1208 	:	val_out <= 4'hb6d0;
         4'h1209 	:	val_out <= 4'hb6d0;
         4'h120a 	:	val_out <= 4'hb6d0;
         4'h120b 	:	val_out <= 4'hb6d0;
         4'h1210 	:	val_out <= 4'hb6e7;
         4'h1211 	:	val_out <= 4'hb6e7;
         4'h1212 	:	val_out <= 4'hb6e7;
         4'h1213 	:	val_out <= 4'hb6e7;
         4'h1218 	:	val_out <= 4'hb6fe;
         4'h1219 	:	val_out <= 4'hb6fe;
         4'h121a 	:	val_out <= 4'hb6fe;
         4'h121b 	:	val_out <= 4'hb6fe;
         4'h1220 	:	val_out <= 4'hb714;
         4'h1221 	:	val_out <= 4'hb714;
         4'h1222 	:	val_out <= 4'hb714;
         4'h1223 	:	val_out <= 4'hb714;
         4'h1228 	:	val_out <= 4'hb72b;
         4'h1229 	:	val_out <= 4'hb72b;
         4'h122a 	:	val_out <= 4'hb72b;
         4'h122b 	:	val_out <= 4'hb72b;
         4'h1230 	:	val_out <= 4'hb742;
         4'h1231 	:	val_out <= 4'hb742;
         4'h1232 	:	val_out <= 4'hb742;
         4'h1233 	:	val_out <= 4'hb742;
         4'h1238 	:	val_out <= 4'hb758;
         4'h1239 	:	val_out <= 4'hb758;
         4'h123a 	:	val_out <= 4'hb758;
         4'h123b 	:	val_out <= 4'hb758;
         4'h1240 	:	val_out <= 4'hb76f;
         4'h1241 	:	val_out <= 4'hb76f;
         4'h1242 	:	val_out <= 4'hb76f;
         4'h1243 	:	val_out <= 4'hb76f;
         4'h1248 	:	val_out <= 4'hb786;
         4'h1249 	:	val_out <= 4'hb786;
         4'h124a 	:	val_out <= 4'hb786;
         4'h124b 	:	val_out <= 4'hb786;
         4'h1250 	:	val_out <= 4'hb79c;
         4'h1251 	:	val_out <= 4'hb79c;
         4'h1252 	:	val_out <= 4'hb79c;
         4'h1253 	:	val_out <= 4'hb79c;
         4'h1258 	:	val_out <= 4'hb7b3;
         4'h1259 	:	val_out <= 4'hb7b3;
         4'h125a 	:	val_out <= 4'hb7b3;
         4'h125b 	:	val_out <= 4'hb7b3;
         4'h1260 	:	val_out <= 4'hb7ca;
         4'h1261 	:	val_out <= 4'hb7ca;
         4'h1262 	:	val_out <= 4'hb7ca;
         4'h1263 	:	val_out <= 4'hb7ca;
         4'h1268 	:	val_out <= 4'hb7e0;
         4'h1269 	:	val_out <= 4'hb7e0;
         4'h126a 	:	val_out <= 4'hb7e0;
         4'h126b 	:	val_out <= 4'hb7e0;
         4'h1270 	:	val_out <= 4'hb7f7;
         4'h1271 	:	val_out <= 4'hb7f7;
         4'h1272 	:	val_out <= 4'hb7f7;
         4'h1273 	:	val_out <= 4'hb7f7;
         4'h1278 	:	val_out <= 4'hb80d;
         4'h1279 	:	val_out <= 4'hb80d;
         4'h127a 	:	val_out <= 4'hb80d;
         4'h127b 	:	val_out <= 4'hb80d;
         4'h1280 	:	val_out <= 4'hb824;
         4'h1281 	:	val_out <= 4'hb824;
         4'h1282 	:	val_out <= 4'hb824;
         4'h1283 	:	val_out <= 4'hb824;
         4'h1288 	:	val_out <= 4'hb83b;
         4'h1289 	:	val_out <= 4'hb83b;
         4'h128a 	:	val_out <= 4'hb83b;
         4'h128b 	:	val_out <= 4'hb83b;
         4'h1290 	:	val_out <= 4'hb851;
         4'h1291 	:	val_out <= 4'hb851;
         4'h1292 	:	val_out <= 4'hb851;
         4'h1293 	:	val_out <= 4'hb851;
         4'h1298 	:	val_out <= 4'hb868;
         4'h1299 	:	val_out <= 4'hb868;
         4'h129a 	:	val_out <= 4'hb868;
         4'h129b 	:	val_out <= 4'hb868;
         4'h12a0 	:	val_out <= 4'hb87e;
         4'h12a1 	:	val_out <= 4'hb87e;
         4'h12a2 	:	val_out <= 4'hb87e;
         4'h12a3 	:	val_out <= 4'hb87e;
         4'h12a8 	:	val_out <= 4'hb895;
         4'h12a9 	:	val_out <= 4'hb895;
         4'h12aa 	:	val_out <= 4'hb895;
         4'h12ab 	:	val_out <= 4'hb895;
         4'h12b0 	:	val_out <= 4'hb8ab;
         4'h12b1 	:	val_out <= 4'hb8ab;
         4'h12b2 	:	val_out <= 4'hb8ab;
         4'h12b3 	:	val_out <= 4'hb8ab;
         4'h12b8 	:	val_out <= 4'hb8c2;
         4'h12b9 	:	val_out <= 4'hb8c2;
         4'h12ba 	:	val_out <= 4'hb8c2;
         4'h12bb 	:	val_out <= 4'hb8c2;
         4'h12c0 	:	val_out <= 4'hb8d8;
         4'h12c1 	:	val_out <= 4'hb8d8;
         4'h12c2 	:	val_out <= 4'hb8d8;
         4'h12c3 	:	val_out <= 4'hb8d8;
         4'h12c8 	:	val_out <= 4'hb8ef;
         4'h12c9 	:	val_out <= 4'hb8ef;
         4'h12ca 	:	val_out <= 4'hb8ef;
         4'h12cb 	:	val_out <= 4'hb8ef;
         4'h12d0 	:	val_out <= 4'hb906;
         4'h12d1 	:	val_out <= 4'hb906;
         4'h12d2 	:	val_out <= 4'hb906;
         4'h12d3 	:	val_out <= 4'hb906;
         4'h12d8 	:	val_out <= 4'hb91c;
         4'h12d9 	:	val_out <= 4'hb91c;
         4'h12da 	:	val_out <= 4'hb91c;
         4'h12db 	:	val_out <= 4'hb91c;
         4'h12e0 	:	val_out <= 4'hb932;
         4'h12e1 	:	val_out <= 4'hb932;
         4'h12e2 	:	val_out <= 4'hb932;
         4'h12e3 	:	val_out <= 4'hb932;
         4'h12e8 	:	val_out <= 4'hb949;
         4'h12e9 	:	val_out <= 4'hb949;
         4'h12ea 	:	val_out <= 4'hb949;
         4'h12eb 	:	val_out <= 4'hb949;
         4'h12f0 	:	val_out <= 4'hb95f;
         4'h12f1 	:	val_out <= 4'hb95f;
         4'h12f2 	:	val_out <= 4'hb95f;
         4'h12f3 	:	val_out <= 4'hb95f;
         4'h12f8 	:	val_out <= 4'hb976;
         4'h12f9 	:	val_out <= 4'hb976;
         4'h12fa 	:	val_out <= 4'hb976;
         4'h12fb 	:	val_out <= 4'hb976;
         4'h1300 	:	val_out <= 4'hb98c;
         4'h1301 	:	val_out <= 4'hb98c;
         4'h1302 	:	val_out <= 4'hb98c;
         4'h1303 	:	val_out <= 4'hb98c;
         4'h1308 	:	val_out <= 4'hb9a3;
         4'h1309 	:	val_out <= 4'hb9a3;
         4'h130a 	:	val_out <= 4'hb9a3;
         4'h130b 	:	val_out <= 4'hb9a3;
         4'h1310 	:	val_out <= 4'hb9b9;
         4'h1311 	:	val_out <= 4'hb9b9;
         4'h1312 	:	val_out <= 4'hb9b9;
         4'h1313 	:	val_out <= 4'hb9b9;
         4'h1318 	:	val_out <= 4'hb9d0;
         4'h1319 	:	val_out <= 4'hb9d0;
         4'h131a 	:	val_out <= 4'hb9d0;
         4'h131b 	:	val_out <= 4'hb9d0;
         4'h1320 	:	val_out <= 4'hb9e6;
         4'h1321 	:	val_out <= 4'hb9e6;
         4'h1322 	:	val_out <= 4'hb9e6;
         4'h1323 	:	val_out <= 4'hb9e6;
         4'h1328 	:	val_out <= 4'hb9fd;
         4'h1329 	:	val_out <= 4'hb9fd;
         4'h132a 	:	val_out <= 4'hb9fd;
         4'h132b 	:	val_out <= 4'hb9fd;
         4'h1330 	:	val_out <= 4'hba13;
         4'h1331 	:	val_out <= 4'hba13;
         4'h1332 	:	val_out <= 4'hba13;
         4'h1333 	:	val_out <= 4'hba13;
         4'h1338 	:	val_out <= 4'hba29;
         4'h1339 	:	val_out <= 4'hba29;
         4'h133a 	:	val_out <= 4'hba29;
         4'h133b 	:	val_out <= 4'hba29;
         4'h1340 	:	val_out <= 4'hba40;
         4'h1341 	:	val_out <= 4'hba40;
         4'h1342 	:	val_out <= 4'hba40;
         4'h1343 	:	val_out <= 4'hba40;
         4'h1348 	:	val_out <= 4'hba56;
         4'h1349 	:	val_out <= 4'hba56;
         4'h134a 	:	val_out <= 4'hba56;
         4'h134b 	:	val_out <= 4'hba56;
         4'h1350 	:	val_out <= 4'hba6c;
         4'h1351 	:	val_out <= 4'hba6c;
         4'h1352 	:	val_out <= 4'hba6c;
         4'h1353 	:	val_out <= 4'hba6c;
         4'h1358 	:	val_out <= 4'hba83;
         4'h1359 	:	val_out <= 4'hba83;
         4'h135a 	:	val_out <= 4'hba83;
         4'h135b 	:	val_out <= 4'hba83;
         4'h1360 	:	val_out <= 4'hba99;
         4'h1361 	:	val_out <= 4'hba99;
         4'h1362 	:	val_out <= 4'hba99;
         4'h1363 	:	val_out <= 4'hba99;
         4'h1368 	:	val_out <= 4'hbaaf;
         4'h1369 	:	val_out <= 4'hbaaf;
         4'h136a 	:	val_out <= 4'hbaaf;
         4'h136b 	:	val_out <= 4'hbaaf;
         4'h1370 	:	val_out <= 4'hbac6;
         4'h1371 	:	val_out <= 4'hbac6;
         4'h1372 	:	val_out <= 4'hbac6;
         4'h1373 	:	val_out <= 4'hbac6;
         4'h1378 	:	val_out <= 4'hbadc;
         4'h1379 	:	val_out <= 4'hbadc;
         4'h137a 	:	val_out <= 4'hbadc;
         4'h137b 	:	val_out <= 4'hbadc;
         4'h1380 	:	val_out <= 4'hbaf2;
         4'h1381 	:	val_out <= 4'hbaf2;
         4'h1382 	:	val_out <= 4'hbaf2;
         4'h1383 	:	val_out <= 4'hbaf2;
         4'h1388 	:	val_out <= 4'hbb09;
         4'h1389 	:	val_out <= 4'hbb09;
         4'h138a 	:	val_out <= 4'hbb09;
         4'h138b 	:	val_out <= 4'hbb09;
         4'h1390 	:	val_out <= 4'hbb1f;
         4'h1391 	:	val_out <= 4'hbb1f;
         4'h1392 	:	val_out <= 4'hbb1f;
         4'h1393 	:	val_out <= 4'hbb1f;
         4'h1398 	:	val_out <= 4'hbb35;
         4'h1399 	:	val_out <= 4'hbb35;
         4'h139a 	:	val_out <= 4'hbb35;
         4'h139b 	:	val_out <= 4'hbb35;
         4'h13a0 	:	val_out <= 4'hbb4c;
         4'h13a1 	:	val_out <= 4'hbb4c;
         4'h13a2 	:	val_out <= 4'hbb4c;
         4'h13a3 	:	val_out <= 4'hbb4c;
         4'h13a8 	:	val_out <= 4'hbb62;
         4'h13a9 	:	val_out <= 4'hbb62;
         4'h13aa 	:	val_out <= 4'hbb62;
         4'h13ab 	:	val_out <= 4'hbb62;
         4'h13b0 	:	val_out <= 4'hbb78;
         4'h13b1 	:	val_out <= 4'hbb78;
         4'h13b2 	:	val_out <= 4'hbb78;
         4'h13b3 	:	val_out <= 4'hbb78;
         4'h13b8 	:	val_out <= 4'hbb8e;
         4'h13b9 	:	val_out <= 4'hbb8e;
         4'h13ba 	:	val_out <= 4'hbb8e;
         4'h13bb 	:	val_out <= 4'hbb8e;
         4'h13c0 	:	val_out <= 4'hbba5;
         4'h13c1 	:	val_out <= 4'hbba5;
         4'h13c2 	:	val_out <= 4'hbba5;
         4'h13c3 	:	val_out <= 4'hbba5;
         4'h13c8 	:	val_out <= 4'hbbbb;
         4'h13c9 	:	val_out <= 4'hbbbb;
         4'h13ca 	:	val_out <= 4'hbbbb;
         4'h13cb 	:	val_out <= 4'hbbbb;
         4'h13d0 	:	val_out <= 4'hbbd1;
         4'h13d1 	:	val_out <= 4'hbbd1;
         4'h13d2 	:	val_out <= 4'hbbd1;
         4'h13d3 	:	val_out <= 4'hbbd1;
         4'h13d8 	:	val_out <= 4'hbbe7;
         4'h13d9 	:	val_out <= 4'hbbe7;
         4'h13da 	:	val_out <= 4'hbbe7;
         4'h13db 	:	val_out <= 4'hbbe7;
         4'h13e0 	:	val_out <= 4'hbbfd;
         4'h13e1 	:	val_out <= 4'hbbfd;
         4'h13e2 	:	val_out <= 4'hbbfd;
         4'h13e3 	:	val_out <= 4'hbbfd;
         4'h13e8 	:	val_out <= 4'hbc14;
         4'h13e9 	:	val_out <= 4'hbc14;
         4'h13ea 	:	val_out <= 4'hbc14;
         4'h13eb 	:	val_out <= 4'hbc14;
         4'h13f0 	:	val_out <= 4'hbc2a;
         4'h13f1 	:	val_out <= 4'hbc2a;
         4'h13f2 	:	val_out <= 4'hbc2a;
         4'h13f3 	:	val_out <= 4'hbc2a;
         4'h13f8 	:	val_out <= 4'hbc40;
         4'h13f9 	:	val_out <= 4'hbc40;
         4'h13fa 	:	val_out <= 4'hbc40;
         4'h13fb 	:	val_out <= 4'hbc40;
         4'h1400 	:	val_out <= 4'hbc56;
         4'h1401 	:	val_out <= 4'hbc56;
         4'h1402 	:	val_out <= 4'hbc56;
         4'h1403 	:	val_out <= 4'hbc56;
         4'h1408 	:	val_out <= 4'hbc6c;
         4'h1409 	:	val_out <= 4'hbc6c;
         4'h140a 	:	val_out <= 4'hbc6c;
         4'h140b 	:	val_out <= 4'hbc6c;
         4'h1410 	:	val_out <= 4'hbc83;
         4'h1411 	:	val_out <= 4'hbc83;
         4'h1412 	:	val_out <= 4'hbc83;
         4'h1413 	:	val_out <= 4'hbc83;
         4'h1418 	:	val_out <= 4'hbc99;
         4'h1419 	:	val_out <= 4'hbc99;
         4'h141a 	:	val_out <= 4'hbc99;
         4'h141b 	:	val_out <= 4'hbc99;
         4'h1420 	:	val_out <= 4'hbcaf;
         4'h1421 	:	val_out <= 4'hbcaf;
         4'h1422 	:	val_out <= 4'hbcaf;
         4'h1423 	:	val_out <= 4'hbcaf;
         4'h1428 	:	val_out <= 4'hbcc5;
         4'h1429 	:	val_out <= 4'hbcc5;
         4'h142a 	:	val_out <= 4'hbcc5;
         4'h142b 	:	val_out <= 4'hbcc5;
         4'h1430 	:	val_out <= 4'hbcdb;
         4'h1431 	:	val_out <= 4'hbcdb;
         4'h1432 	:	val_out <= 4'hbcdb;
         4'h1433 	:	val_out <= 4'hbcdb;
         4'h1438 	:	val_out <= 4'hbcf1;
         4'h1439 	:	val_out <= 4'hbcf1;
         4'h143a 	:	val_out <= 4'hbcf1;
         4'h143b 	:	val_out <= 4'hbcf1;
         4'h1440 	:	val_out <= 4'hbd07;
         4'h1441 	:	val_out <= 4'hbd07;
         4'h1442 	:	val_out <= 4'hbd07;
         4'h1443 	:	val_out <= 4'hbd07;
         4'h1448 	:	val_out <= 4'hbd1d;
         4'h1449 	:	val_out <= 4'hbd1d;
         4'h144a 	:	val_out <= 4'hbd1d;
         4'h144b 	:	val_out <= 4'hbd1d;
         4'h1450 	:	val_out <= 4'hbd33;
         4'h1451 	:	val_out <= 4'hbd33;
         4'h1452 	:	val_out <= 4'hbd33;
         4'h1453 	:	val_out <= 4'hbd33;
         4'h1458 	:	val_out <= 4'hbd49;
         4'h1459 	:	val_out <= 4'hbd49;
         4'h145a 	:	val_out <= 4'hbd49;
         4'h145b 	:	val_out <= 4'hbd49;
         4'h1460 	:	val_out <= 4'hbd60;
         4'h1461 	:	val_out <= 4'hbd60;
         4'h1462 	:	val_out <= 4'hbd60;
         4'h1463 	:	val_out <= 4'hbd60;
         4'h1468 	:	val_out <= 4'hbd76;
         4'h1469 	:	val_out <= 4'hbd76;
         4'h146a 	:	val_out <= 4'hbd76;
         4'h146b 	:	val_out <= 4'hbd76;
         4'h1470 	:	val_out <= 4'hbd8c;
         4'h1471 	:	val_out <= 4'hbd8c;
         4'h1472 	:	val_out <= 4'hbd8c;
         4'h1473 	:	val_out <= 4'hbd8c;
         4'h1478 	:	val_out <= 4'hbda2;
         4'h1479 	:	val_out <= 4'hbda2;
         4'h147a 	:	val_out <= 4'hbda2;
         4'h147b 	:	val_out <= 4'hbda2;
         4'h1480 	:	val_out <= 4'hbdb8;
         4'h1481 	:	val_out <= 4'hbdb8;
         4'h1482 	:	val_out <= 4'hbdb8;
         4'h1483 	:	val_out <= 4'hbdb8;
         4'h1488 	:	val_out <= 4'hbdce;
         4'h1489 	:	val_out <= 4'hbdce;
         4'h148a 	:	val_out <= 4'hbdce;
         4'h148b 	:	val_out <= 4'hbdce;
         4'h1490 	:	val_out <= 4'hbde4;
         4'h1491 	:	val_out <= 4'hbde4;
         4'h1492 	:	val_out <= 4'hbde4;
         4'h1493 	:	val_out <= 4'hbde4;
         4'h1498 	:	val_out <= 4'hbdfa;
         4'h1499 	:	val_out <= 4'hbdfa;
         4'h149a 	:	val_out <= 4'hbdfa;
         4'h149b 	:	val_out <= 4'hbdfa;
         4'h14a0 	:	val_out <= 4'hbe10;
         4'h14a1 	:	val_out <= 4'hbe10;
         4'h14a2 	:	val_out <= 4'hbe10;
         4'h14a3 	:	val_out <= 4'hbe10;
         4'h14a8 	:	val_out <= 4'hbe26;
         4'h14a9 	:	val_out <= 4'hbe26;
         4'h14aa 	:	val_out <= 4'hbe26;
         4'h14ab 	:	val_out <= 4'hbe26;
         4'h14b0 	:	val_out <= 4'hbe3c;
         4'h14b1 	:	val_out <= 4'hbe3c;
         4'h14b2 	:	val_out <= 4'hbe3c;
         4'h14b3 	:	val_out <= 4'hbe3c;
         4'h14b8 	:	val_out <= 4'hbe52;
         4'h14b9 	:	val_out <= 4'hbe52;
         4'h14ba 	:	val_out <= 4'hbe52;
         4'h14bb 	:	val_out <= 4'hbe52;
         4'h14c0 	:	val_out <= 4'hbe68;
         4'h14c1 	:	val_out <= 4'hbe68;
         4'h14c2 	:	val_out <= 4'hbe68;
         4'h14c3 	:	val_out <= 4'hbe68;
         4'h14c8 	:	val_out <= 4'hbe7d;
         4'h14c9 	:	val_out <= 4'hbe7d;
         4'h14ca 	:	val_out <= 4'hbe7d;
         4'h14cb 	:	val_out <= 4'hbe7d;
         4'h14d0 	:	val_out <= 4'hbe93;
         4'h14d1 	:	val_out <= 4'hbe93;
         4'h14d2 	:	val_out <= 4'hbe93;
         4'h14d3 	:	val_out <= 4'hbe93;
         4'h14d8 	:	val_out <= 4'hbea9;
         4'h14d9 	:	val_out <= 4'hbea9;
         4'h14da 	:	val_out <= 4'hbea9;
         4'h14db 	:	val_out <= 4'hbea9;
         4'h14e0 	:	val_out <= 4'hbebf;
         4'h14e1 	:	val_out <= 4'hbebf;
         4'h14e2 	:	val_out <= 4'hbebf;
         4'h14e3 	:	val_out <= 4'hbebf;
         4'h14e8 	:	val_out <= 4'hbed5;
         4'h14e9 	:	val_out <= 4'hbed5;
         4'h14ea 	:	val_out <= 4'hbed5;
         4'h14eb 	:	val_out <= 4'hbed5;
         4'h14f0 	:	val_out <= 4'hbeeb;
         4'h14f1 	:	val_out <= 4'hbeeb;
         4'h14f2 	:	val_out <= 4'hbeeb;
         4'h14f3 	:	val_out <= 4'hbeeb;
         4'h14f8 	:	val_out <= 4'hbf01;
         4'h14f9 	:	val_out <= 4'hbf01;
         4'h14fa 	:	val_out <= 4'hbf01;
         4'h14fb 	:	val_out <= 4'hbf01;
         4'h1500 	:	val_out <= 4'hbf17;
         4'h1501 	:	val_out <= 4'hbf17;
         4'h1502 	:	val_out <= 4'hbf17;
         4'h1503 	:	val_out <= 4'hbf17;
         4'h1508 	:	val_out <= 4'hbf2d;
         4'h1509 	:	val_out <= 4'hbf2d;
         4'h150a 	:	val_out <= 4'hbf2d;
         4'h150b 	:	val_out <= 4'hbf2d;
         4'h1510 	:	val_out <= 4'hbf43;
         4'h1511 	:	val_out <= 4'hbf43;
         4'h1512 	:	val_out <= 4'hbf43;
         4'h1513 	:	val_out <= 4'hbf43;
         4'h1518 	:	val_out <= 4'hbf58;
         4'h1519 	:	val_out <= 4'hbf58;
         4'h151a 	:	val_out <= 4'hbf58;
         4'h151b 	:	val_out <= 4'hbf58;
         4'h1520 	:	val_out <= 4'hbf6e;
         4'h1521 	:	val_out <= 4'hbf6e;
         4'h1522 	:	val_out <= 4'hbf6e;
         4'h1523 	:	val_out <= 4'hbf6e;
         4'h1528 	:	val_out <= 4'hbf84;
         4'h1529 	:	val_out <= 4'hbf84;
         4'h152a 	:	val_out <= 4'hbf84;
         4'h152b 	:	val_out <= 4'hbf84;
         4'h1530 	:	val_out <= 4'hbf9a;
         4'h1531 	:	val_out <= 4'hbf9a;
         4'h1532 	:	val_out <= 4'hbf9a;
         4'h1533 	:	val_out <= 4'hbf9a;
         4'h1538 	:	val_out <= 4'hbfb0;
         4'h1539 	:	val_out <= 4'hbfb0;
         4'h153a 	:	val_out <= 4'hbfb0;
         4'h153b 	:	val_out <= 4'hbfb0;
         4'h1540 	:	val_out <= 4'hbfc5;
         4'h1541 	:	val_out <= 4'hbfc5;
         4'h1542 	:	val_out <= 4'hbfc5;
         4'h1543 	:	val_out <= 4'hbfc5;
         4'h1548 	:	val_out <= 4'hbfdb;
         4'h1549 	:	val_out <= 4'hbfdb;
         4'h154a 	:	val_out <= 4'hbfdb;
         4'h154b 	:	val_out <= 4'hbfdb;
         4'h1550 	:	val_out <= 4'hbff1;
         4'h1551 	:	val_out <= 4'hbff1;
         4'h1552 	:	val_out <= 4'hbff1;
         4'h1553 	:	val_out <= 4'hbff1;
         4'h1558 	:	val_out <= 4'hc007;
         4'h1559 	:	val_out <= 4'hc007;
         4'h155a 	:	val_out <= 4'hc007;
         4'h155b 	:	val_out <= 4'hc007;
         4'h1560 	:	val_out <= 4'hc01d;
         4'h1561 	:	val_out <= 4'hc01d;
         4'h1562 	:	val_out <= 4'hc01d;
         4'h1563 	:	val_out <= 4'hc01d;
         4'h1568 	:	val_out <= 4'hc032;
         4'h1569 	:	val_out <= 4'hc032;
         4'h156a 	:	val_out <= 4'hc032;
         4'h156b 	:	val_out <= 4'hc032;
         4'h1570 	:	val_out <= 4'hc048;
         4'h1571 	:	val_out <= 4'hc048;
         4'h1572 	:	val_out <= 4'hc048;
         4'h1573 	:	val_out <= 4'hc048;
         4'h1578 	:	val_out <= 4'hc05e;
         4'h1579 	:	val_out <= 4'hc05e;
         4'h157a 	:	val_out <= 4'hc05e;
         4'h157b 	:	val_out <= 4'hc05e;
         4'h1580 	:	val_out <= 4'hc073;
         4'h1581 	:	val_out <= 4'hc073;
         4'h1582 	:	val_out <= 4'hc073;
         4'h1583 	:	val_out <= 4'hc073;
         4'h1588 	:	val_out <= 4'hc089;
         4'h1589 	:	val_out <= 4'hc089;
         4'h158a 	:	val_out <= 4'hc089;
         4'h158b 	:	val_out <= 4'hc089;
         4'h1590 	:	val_out <= 4'hc09f;
         4'h1591 	:	val_out <= 4'hc09f;
         4'h1592 	:	val_out <= 4'hc09f;
         4'h1593 	:	val_out <= 4'hc09f;
         4'h1598 	:	val_out <= 4'hc0b5;
         4'h1599 	:	val_out <= 4'hc0b5;
         4'h159a 	:	val_out <= 4'hc0b5;
         4'h159b 	:	val_out <= 4'hc0b5;
         4'h15a0 	:	val_out <= 4'hc0ca;
         4'h15a1 	:	val_out <= 4'hc0ca;
         4'h15a2 	:	val_out <= 4'hc0ca;
         4'h15a3 	:	val_out <= 4'hc0ca;
         4'h15a8 	:	val_out <= 4'hc0e0;
         4'h15a9 	:	val_out <= 4'hc0e0;
         4'h15aa 	:	val_out <= 4'hc0e0;
         4'h15ab 	:	val_out <= 4'hc0e0;
         4'h15b0 	:	val_out <= 4'hc0f6;
         4'h15b1 	:	val_out <= 4'hc0f6;
         4'h15b2 	:	val_out <= 4'hc0f6;
         4'h15b3 	:	val_out <= 4'hc0f6;
         4'h15b8 	:	val_out <= 4'hc10b;
         4'h15b9 	:	val_out <= 4'hc10b;
         4'h15ba 	:	val_out <= 4'hc10b;
         4'h15bb 	:	val_out <= 4'hc10b;
         4'h15c0 	:	val_out <= 4'hc121;
         4'h15c1 	:	val_out <= 4'hc121;
         4'h15c2 	:	val_out <= 4'hc121;
         4'h15c3 	:	val_out <= 4'hc121;
         4'h15c8 	:	val_out <= 4'hc136;
         4'h15c9 	:	val_out <= 4'hc136;
         4'h15ca 	:	val_out <= 4'hc136;
         4'h15cb 	:	val_out <= 4'hc136;
         4'h15d0 	:	val_out <= 4'hc14c;
         4'h15d1 	:	val_out <= 4'hc14c;
         4'h15d2 	:	val_out <= 4'hc14c;
         4'h15d3 	:	val_out <= 4'hc14c;
         4'h15d8 	:	val_out <= 4'hc162;
         4'h15d9 	:	val_out <= 4'hc162;
         4'h15da 	:	val_out <= 4'hc162;
         4'h15db 	:	val_out <= 4'hc162;
         4'h15e0 	:	val_out <= 4'hc177;
         4'h15e1 	:	val_out <= 4'hc177;
         4'h15e2 	:	val_out <= 4'hc177;
         4'h15e3 	:	val_out <= 4'hc177;
         4'h15e8 	:	val_out <= 4'hc18d;
         4'h15e9 	:	val_out <= 4'hc18d;
         4'h15ea 	:	val_out <= 4'hc18d;
         4'h15eb 	:	val_out <= 4'hc18d;
         4'h15f0 	:	val_out <= 4'hc1a2;
         4'h15f1 	:	val_out <= 4'hc1a2;
         4'h15f2 	:	val_out <= 4'hc1a2;
         4'h15f3 	:	val_out <= 4'hc1a2;
         4'h15f8 	:	val_out <= 4'hc1b8;
         4'h15f9 	:	val_out <= 4'hc1b8;
         4'h15fa 	:	val_out <= 4'hc1b8;
         4'h15fb 	:	val_out <= 4'hc1b8;
         4'h1600 	:	val_out <= 4'hc1ce;
         4'h1601 	:	val_out <= 4'hc1ce;
         4'h1602 	:	val_out <= 4'hc1ce;
         4'h1603 	:	val_out <= 4'hc1ce;
         4'h1608 	:	val_out <= 4'hc1e3;
         4'h1609 	:	val_out <= 4'hc1e3;
         4'h160a 	:	val_out <= 4'hc1e3;
         4'h160b 	:	val_out <= 4'hc1e3;
         4'h1610 	:	val_out <= 4'hc1f9;
         4'h1611 	:	val_out <= 4'hc1f9;
         4'h1612 	:	val_out <= 4'hc1f9;
         4'h1613 	:	val_out <= 4'hc1f9;
         4'h1618 	:	val_out <= 4'hc20e;
         4'h1619 	:	val_out <= 4'hc20e;
         4'h161a 	:	val_out <= 4'hc20e;
         4'h161b 	:	val_out <= 4'hc20e;
         4'h1620 	:	val_out <= 4'hc224;
         4'h1621 	:	val_out <= 4'hc224;
         4'h1622 	:	val_out <= 4'hc224;
         4'h1623 	:	val_out <= 4'hc224;
         4'h1628 	:	val_out <= 4'hc239;
         4'h1629 	:	val_out <= 4'hc239;
         4'h162a 	:	val_out <= 4'hc239;
         4'h162b 	:	val_out <= 4'hc239;
         4'h1630 	:	val_out <= 4'hc24f;
         4'h1631 	:	val_out <= 4'hc24f;
         4'h1632 	:	val_out <= 4'hc24f;
         4'h1633 	:	val_out <= 4'hc24f;
         4'h1638 	:	val_out <= 4'hc264;
         4'h1639 	:	val_out <= 4'hc264;
         4'h163a 	:	val_out <= 4'hc264;
         4'h163b 	:	val_out <= 4'hc264;
         4'h1640 	:	val_out <= 4'hc27a;
         4'h1641 	:	val_out <= 4'hc27a;
         4'h1642 	:	val_out <= 4'hc27a;
         4'h1643 	:	val_out <= 4'hc27a;
         4'h1648 	:	val_out <= 4'hc28f;
         4'h1649 	:	val_out <= 4'hc28f;
         4'h164a 	:	val_out <= 4'hc28f;
         4'h164b 	:	val_out <= 4'hc28f;
         4'h1650 	:	val_out <= 4'hc2a5;
         4'h1651 	:	val_out <= 4'hc2a5;
         4'h1652 	:	val_out <= 4'hc2a5;
         4'h1653 	:	val_out <= 4'hc2a5;
         4'h1658 	:	val_out <= 4'hc2ba;
         4'h1659 	:	val_out <= 4'hc2ba;
         4'h165a 	:	val_out <= 4'hc2ba;
         4'h165b 	:	val_out <= 4'hc2ba;
         4'h1660 	:	val_out <= 4'hc2d0;
         4'h1661 	:	val_out <= 4'hc2d0;
         4'h1662 	:	val_out <= 4'hc2d0;
         4'h1663 	:	val_out <= 4'hc2d0;
         4'h1668 	:	val_out <= 4'hc2e5;
         4'h1669 	:	val_out <= 4'hc2e5;
         4'h166a 	:	val_out <= 4'hc2e5;
         4'h166b 	:	val_out <= 4'hc2e5;
         4'h1670 	:	val_out <= 4'hc2fa;
         4'h1671 	:	val_out <= 4'hc2fa;
         4'h1672 	:	val_out <= 4'hc2fa;
         4'h1673 	:	val_out <= 4'hc2fa;
         4'h1678 	:	val_out <= 4'hc310;
         4'h1679 	:	val_out <= 4'hc310;
         4'h167a 	:	val_out <= 4'hc310;
         4'h167b 	:	val_out <= 4'hc310;
         4'h1680 	:	val_out <= 4'hc325;
         4'h1681 	:	val_out <= 4'hc325;
         4'h1682 	:	val_out <= 4'hc325;
         4'h1683 	:	val_out <= 4'hc325;
         4'h1688 	:	val_out <= 4'hc33b;
         4'h1689 	:	val_out <= 4'hc33b;
         4'h168a 	:	val_out <= 4'hc33b;
         4'h168b 	:	val_out <= 4'hc33b;
         4'h1690 	:	val_out <= 4'hc350;
         4'h1691 	:	val_out <= 4'hc350;
         4'h1692 	:	val_out <= 4'hc350;
         4'h1693 	:	val_out <= 4'hc350;
         4'h1698 	:	val_out <= 4'hc365;
         4'h1699 	:	val_out <= 4'hc365;
         4'h169a 	:	val_out <= 4'hc365;
         4'h169b 	:	val_out <= 4'hc365;
         4'h16a0 	:	val_out <= 4'hc37b;
         4'h16a1 	:	val_out <= 4'hc37b;
         4'h16a2 	:	val_out <= 4'hc37b;
         4'h16a3 	:	val_out <= 4'hc37b;
         4'h16a8 	:	val_out <= 4'hc390;
         4'h16a9 	:	val_out <= 4'hc390;
         4'h16aa 	:	val_out <= 4'hc390;
         4'h16ab 	:	val_out <= 4'hc390;
         4'h16b0 	:	val_out <= 4'hc3a5;
         4'h16b1 	:	val_out <= 4'hc3a5;
         4'h16b2 	:	val_out <= 4'hc3a5;
         4'h16b3 	:	val_out <= 4'hc3a5;
         4'h16b8 	:	val_out <= 4'hc3bb;
         4'h16b9 	:	val_out <= 4'hc3bb;
         4'h16ba 	:	val_out <= 4'hc3bb;
         4'h16bb 	:	val_out <= 4'hc3bb;
         4'h16c0 	:	val_out <= 4'hc3d0;
         4'h16c1 	:	val_out <= 4'hc3d0;
         4'h16c2 	:	val_out <= 4'hc3d0;
         4'h16c3 	:	val_out <= 4'hc3d0;
         4'h16c8 	:	val_out <= 4'hc3e5;
         4'h16c9 	:	val_out <= 4'hc3e5;
         4'h16ca 	:	val_out <= 4'hc3e5;
         4'h16cb 	:	val_out <= 4'hc3e5;
         4'h16d0 	:	val_out <= 4'hc3fb;
         4'h16d1 	:	val_out <= 4'hc3fb;
         4'h16d2 	:	val_out <= 4'hc3fb;
         4'h16d3 	:	val_out <= 4'hc3fb;
         4'h16d8 	:	val_out <= 4'hc410;
         4'h16d9 	:	val_out <= 4'hc410;
         4'h16da 	:	val_out <= 4'hc410;
         4'h16db 	:	val_out <= 4'hc410;
         4'h16e0 	:	val_out <= 4'hc425;
         4'h16e1 	:	val_out <= 4'hc425;
         4'h16e2 	:	val_out <= 4'hc425;
         4'h16e3 	:	val_out <= 4'hc425;
         4'h16e8 	:	val_out <= 4'hc43b;
         4'h16e9 	:	val_out <= 4'hc43b;
         4'h16ea 	:	val_out <= 4'hc43b;
         4'h16eb 	:	val_out <= 4'hc43b;
         4'h16f0 	:	val_out <= 4'hc450;
         4'h16f1 	:	val_out <= 4'hc450;
         4'h16f2 	:	val_out <= 4'hc450;
         4'h16f3 	:	val_out <= 4'hc450;
         4'h16f8 	:	val_out <= 4'hc465;
         4'h16f9 	:	val_out <= 4'hc465;
         4'h16fa 	:	val_out <= 4'hc465;
         4'h16fb 	:	val_out <= 4'hc465;
         4'h1700 	:	val_out <= 4'hc47a;
         4'h1701 	:	val_out <= 4'hc47a;
         4'h1702 	:	val_out <= 4'hc47a;
         4'h1703 	:	val_out <= 4'hc47a;
         4'h1708 	:	val_out <= 4'hc490;
         4'h1709 	:	val_out <= 4'hc490;
         4'h170a 	:	val_out <= 4'hc490;
         4'h170b 	:	val_out <= 4'hc490;
         4'h1710 	:	val_out <= 4'hc4a5;
         4'h1711 	:	val_out <= 4'hc4a5;
         4'h1712 	:	val_out <= 4'hc4a5;
         4'h1713 	:	val_out <= 4'hc4a5;
         4'h1718 	:	val_out <= 4'hc4ba;
         4'h1719 	:	val_out <= 4'hc4ba;
         4'h171a 	:	val_out <= 4'hc4ba;
         4'h171b 	:	val_out <= 4'hc4ba;
         4'h1720 	:	val_out <= 4'hc4cf;
         4'h1721 	:	val_out <= 4'hc4cf;
         4'h1722 	:	val_out <= 4'hc4cf;
         4'h1723 	:	val_out <= 4'hc4cf;
         4'h1728 	:	val_out <= 4'hc4e4;
         4'h1729 	:	val_out <= 4'hc4e4;
         4'h172a 	:	val_out <= 4'hc4e4;
         4'h172b 	:	val_out <= 4'hc4e4;
         4'h1730 	:	val_out <= 4'hc4fa;
         4'h1731 	:	val_out <= 4'hc4fa;
         4'h1732 	:	val_out <= 4'hc4fa;
         4'h1733 	:	val_out <= 4'hc4fa;
         4'h1738 	:	val_out <= 4'hc50f;
         4'h1739 	:	val_out <= 4'hc50f;
         4'h173a 	:	val_out <= 4'hc50f;
         4'h173b 	:	val_out <= 4'hc50f;
         4'h1740 	:	val_out <= 4'hc524;
         4'h1741 	:	val_out <= 4'hc524;
         4'h1742 	:	val_out <= 4'hc524;
         4'h1743 	:	val_out <= 4'hc524;
         4'h1748 	:	val_out <= 4'hc539;
         4'h1749 	:	val_out <= 4'hc539;
         4'h174a 	:	val_out <= 4'hc539;
         4'h174b 	:	val_out <= 4'hc539;
         4'h1750 	:	val_out <= 4'hc54e;
         4'h1751 	:	val_out <= 4'hc54e;
         4'h1752 	:	val_out <= 4'hc54e;
         4'h1753 	:	val_out <= 4'hc54e;
         4'h1758 	:	val_out <= 4'hc563;
         4'h1759 	:	val_out <= 4'hc563;
         4'h175a 	:	val_out <= 4'hc563;
         4'h175b 	:	val_out <= 4'hc563;
         4'h1760 	:	val_out <= 4'hc578;
         4'h1761 	:	val_out <= 4'hc578;
         4'h1762 	:	val_out <= 4'hc578;
         4'h1763 	:	val_out <= 4'hc578;
         4'h1768 	:	val_out <= 4'hc58d;
         4'h1769 	:	val_out <= 4'hc58d;
         4'h176a 	:	val_out <= 4'hc58d;
         4'h176b 	:	val_out <= 4'hc58d;
         4'h1770 	:	val_out <= 4'hc5a3;
         4'h1771 	:	val_out <= 4'hc5a3;
         4'h1772 	:	val_out <= 4'hc5a3;
         4'h1773 	:	val_out <= 4'hc5a3;
         4'h1778 	:	val_out <= 4'hc5b8;
         4'h1779 	:	val_out <= 4'hc5b8;
         4'h177a 	:	val_out <= 4'hc5b8;
         4'h177b 	:	val_out <= 4'hc5b8;
         4'h1780 	:	val_out <= 4'hc5cd;
         4'h1781 	:	val_out <= 4'hc5cd;
         4'h1782 	:	val_out <= 4'hc5cd;
         4'h1783 	:	val_out <= 4'hc5cd;
         4'h1788 	:	val_out <= 4'hc5e2;
         4'h1789 	:	val_out <= 4'hc5e2;
         4'h178a 	:	val_out <= 4'hc5e2;
         4'h178b 	:	val_out <= 4'hc5e2;
         4'h1790 	:	val_out <= 4'hc5f7;
         4'h1791 	:	val_out <= 4'hc5f7;
         4'h1792 	:	val_out <= 4'hc5f7;
         4'h1793 	:	val_out <= 4'hc5f7;
         4'h1798 	:	val_out <= 4'hc60c;
         4'h1799 	:	val_out <= 4'hc60c;
         4'h179a 	:	val_out <= 4'hc60c;
         4'h179b 	:	val_out <= 4'hc60c;
         4'h17a0 	:	val_out <= 4'hc621;
         4'h17a1 	:	val_out <= 4'hc621;
         4'h17a2 	:	val_out <= 4'hc621;
         4'h17a3 	:	val_out <= 4'hc621;
         4'h17a8 	:	val_out <= 4'hc636;
         4'h17a9 	:	val_out <= 4'hc636;
         4'h17aa 	:	val_out <= 4'hc636;
         4'h17ab 	:	val_out <= 4'hc636;
         4'h17b0 	:	val_out <= 4'hc64b;
         4'h17b1 	:	val_out <= 4'hc64b;
         4'h17b2 	:	val_out <= 4'hc64b;
         4'h17b3 	:	val_out <= 4'hc64b;
         4'h17b8 	:	val_out <= 4'hc660;
         4'h17b9 	:	val_out <= 4'hc660;
         4'h17ba 	:	val_out <= 4'hc660;
         4'h17bb 	:	val_out <= 4'hc660;
         4'h17c0 	:	val_out <= 4'hc675;
         4'h17c1 	:	val_out <= 4'hc675;
         4'h17c2 	:	val_out <= 4'hc675;
         4'h17c3 	:	val_out <= 4'hc675;
         4'h17c8 	:	val_out <= 4'hc68a;
         4'h17c9 	:	val_out <= 4'hc68a;
         4'h17ca 	:	val_out <= 4'hc68a;
         4'h17cb 	:	val_out <= 4'hc68a;
         4'h17d0 	:	val_out <= 4'hc69f;
         4'h17d1 	:	val_out <= 4'hc69f;
         4'h17d2 	:	val_out <= 4'hc69f;
         4'h17d3 	:	val_out <= 4'hc69f;
         4'h17d8 	:	val_out <= 4'hc6b4;
         4'h17d9 	:	val_out <= 4'hc6b4;
         4'h17da 	:	val_out <= 4'hc6b4;
         4'h17db 	:	val_out <= 4'hc6b4;
         4'h17e0 	:	val_out <= 4'hc6c9;
         4'h17e1 	:	val_out <= 4'hc6c9;
         4'h17e2 	:	val_out <= 4'hc6c9;
         4'h17e3 	:	val_out <= 4'hc6c9;
         4'h17e8 	:	val_out <= 4'hc6de;
         4'h17e9 	:	val_out <= 4'hc6de;
         4'h17ea 	:	val_out <= 4'hc6de;
         4'h17eb 	:	val_out <= 4'hc6de;
         4'h17f0 	:	val_out <= 4'hc6f3;
         4'h17f1 	:	val_out <= 4'hc6f3;
         4'h17f2 	:	val_out <= 4'hc6f3;
         4'h17f3 	:	val_out <= 4'hc6f3;
         4'h17f8 	:	val_out <= 4'hc708;
         4'h17f9 	:	val_out <= 4'hc708;
         4'h17fa 	:	val_out <= 4'hc708;
         4'h17fb 	:	val_out <= 4'hc708;
         4'h1800 	:	val_out <= 4'hc71c;
         4'h1801 	:	val_out <= 4'hc71c;
         4'h1802 	:	val_out <= 4'hc71c;
         4'h1803 	:	val_out <= 4'hc71c;
         4'h1808 	:	val_out <= 4'hc731;
         4'h1809 	:	val_out <= 4'hc731;
         4'h180a 	:	val_out <= 4'hc731;
         4'h180b 	:	val_out <= 4'hc731;
         4'h1810 	:	val_out <= 4'hc746;
         4'h1811 	:	val_out <= 4'hc746;
         4'h1812 	:	val_out <= 4'hc746;
         4'h1813 	:	val_out <= 4'hc746;
         4'h1818 	:	val_out <= 4'hc75b;
         4'h1819 	:	val_out <= 4'hc75b;
         4'h181a 	:	val_out <= 4'hc75b;
         4'h181b 	:	val_out <= 4'hc75b;
         4'h1820 	:	val_out <= 4'hc770;
         4'h1821 	:	val_out <= 4'hc770;
         4'h1822 	:	val_out <= 4'hc770;
         4'h1823 	:	val_out <= 4'hc770;
         4'h1828 	:	val_out <= 4'hc785;
         4'h1829 	:	val_out <= 4'hc785;
         4'h182a 	:	val_out <= 4'hc785;
         4'h182b 	:	val_out <= 4'hc785;
         4'h1830 	:	val_out <= 4'hc79a;
         4'h1831 	:	val_out <= 4'hc79a;
         4'h1832 	:	val_out <= 4'hc79a;
         4'h1833 	:	val_out <= 4'hc79a;
         4'h1838 	:	val_out <= 4'hc7ae;
         4'h1839 	:	val_out <= 4'hc7ae;
         4'h183a 	:	val_out <= 4'hc7ae;
         4'h183b 	:	val_out <= 4'hc7ae;
         4'h1840 	:	val_out <= 4'hc7c3;
         4'h1841 	:	val_out <= 4'hc7c3;
         4'h1842 	:	val_out <= 4'hc7c3;
         4'h1843 	:	val_out <= 4'hc7c3;
         4'h1848 	:	val_out <= 4'hc7d8;
         4'h1849 	:	val_out <= 4'hc7d8;
         4'h184a 	:	val_out <= 4'hc7d8;
         4'h184b 	:	val_out <= 4'hc7d8;
         4'h1850 	:	val_out <= 4'hc7ed;
         4'h1851 	:	val_out <= 4'hc7ed;
         4'h1852 	:	val_out <= 4'hc7ed;
         4'h1853 	:	val_out <= 4'hc7ed;
         4'h1858 	:	val_out <= 4'hc802;
         4'h1859 	:	val_out <= 4'hc802;
         4'h185a 	:	val_out <= 4'hc802;
         4'h185b 	:	val_out <= 4'hc802;
         4'h1860 	:	val_out <= 4'hc816;
         4'h1861 	:	val_out <= 4'hc816;
         4'h1862 	:	val_out <= 4'hc816;
         4'h1863 	:	val_out <= 4'hc816;
         4'h1868 	:	val_out <= 4'hc82b;
         4'h1869 	:	val_out <= 4'hc82b;
         4'h186a 	:	val_out <= 4'hc82b;
         4'h186b 	:	val_out <= 4'hc82b;
         4'h1870 	:	val_out <= 4'hc840;
         4'h1871 	:	val_out <= 4'hc840;
         4'h1872 	:	val_out <= 4'hc840;
         4'h1873 	:	val_out <= 4'hc840;
         4'h1878 	:	val_out <= 4'hc855;
         4'h1879 	:	val_out <= 4'hc855;
         4'h187a 	:	val_out <= 4'hc855;
         4'h187b 	:	val_out <= 4'hc855;
         4'h1880 	:	val_out <= 4'hc869;
         4'h1881 	:	val_out <= 4'hc869;
         4'h1882 	:	val_out <= 4'hc869;
         4'h1883 	:	val_out <= 4'hc869;
         4'h1888 	:	val_out <= 4'hc87e;
         4'h1889 	:	val_out <= 4'hc87e;
         4'h188a 	:	val_out <= 4'hc87e;
         4'h188b 	:	val_out <= 4'hc87e;
         4'h1890 	:	val_out <= 4'hc893;
         4'h1891 	:	val_out <= 4'hc893;
         4'h1892 	:	val_out <= 4'hc893;
         4'h1893 	:	val_out <= 4'hc893;
         4'h1898 	:	val_out <= 4'hc8a8;
         4'h1899 	:	val_out <= 4'hc8a8;
         4'h189a 	:	val_out <= 4'hc8a8;
         4'h189b 	:	val_out <= 4'hc8a8;
         4'h18a0 	:	val_out <= 4'hc8bc;
         4'h18a1 	:	val_out <= 4'hc8bc;
         4'h18a2 	:	val_out <= 4'hc8bc;
         4'h18a3 	:	val_out <= 4'hc8bc;
         4'h18a8 	:	val_out <= 4'hc8d1;
         4'h18a9 	:	val_out <= 4'hc8d1;
         4'h18aa 	:	val_out <= 4'hc8d1;
         4'h18ab 	:	val_out <= 4'hc8d1;
         4'h18b0 	:	val_out <= 4'hc8e6;
         4'h18b1 	:	val_out <= 4'hc8e6;
         4'h18b2 	:	val_out <= 4'hc8e6;
         4'h18b3 	:	val_out <= 4'hc8e6;
         4'h18b8 	:	val_out <= 4'hc8fa;
         4'h18b9 	:	val_out <= 4'hc8fa;
         4'h18ba 	:	val_out <= 4'hc8fa;
         4'h18bb 	:	val_out <= 4'hc8fa;
         4'h18c0 	:	val_out <= 4'hc90f;
         4'h18c1 	:	val_out <= 4'hc90f;
         4'h18c2 	:	val_out <= 4'hc90f;
         4'h18c3 	:	val_out <= 4'hc90f;
         4'h18c8 	:	val_out <= 4'hc923;
         4'h18c9 	:	val_out <= 4'hc923;
         4'h18ca 	:	val_out <= 4'hc923;
         4'h18cb 	:	val_out <= 4'hc923;
         4'h18d0 	:	val_out <= 4'hc938;
         4'h18d1 	:	val_out <= 4'hc938;
         4'h18d2 	:	val_out <= 4'hc938;
         4'h18d3 	:	val_out <= 4'hc938;
         4'h18d8 	:	val_out <= 4'hc94d;
         4'h18d9 	:	val_out <= 4'hc94d;
         4'h18da 	:	val_out <= 4'hc94d;
         4'h18db 	:	val_out <= 4'hc94d;
         4'h18e0 	:	val_out <= 4'hc961;
         4'h18e1 	:	val_out <= 4'hc961;
         4'h18e2 	:	val_out <= 4'hc961;
         4'h18e3 	:	val_out <= 4'hc961;
         4'h18e8 	:	val_out <= 4'hc976;
         4'h18e9 	:	val_out <= 4'hc976;
         4'h18ea 	:	val_out <= 4'hc976;
         4'h18eb 	:	val_out <= 4'hc976;
         4'h18f0 	:	val_out <= 4'hc98a;
         4'h18f1 	:	val_out <= 4'hc98a;
         4'h18f2 	:	val_out <= 4'hc98a;
         4'h18f3 	:	val_out <= 4'hc98a;
         4'h18f8 	:	val_out <= 4'hc99f;
         4'h18f9 	:	val_out <= 4'hc99f;
         4'h18fa 	:	val_out <= 4'hc99f;
         4'h18fb 	:	val_out <= 4'hc99f;
         4'h1900 	:	val_out <= 4'hc9b4;
         4'h1901 	:	val_out <= 4'hc9b4;
         4'h1902 	:	val_out <= 4'hc9b4;
         4'h1903 	:	val_out <= 4'hc9b4;
         4'h1908 	:	val_out <= 4'hc9c8;
         4'h1909 	:	val_out <= 4'hc9c8;
         4'h190a 	:	val_out <= 4'hc9c8;
         4'h190b 	:	val_out <= 4'hc9c8;
         4'h1910 	:	val_out <= 4'hc9dd;
         4'h1911 	:	val_out <= 4'hc9dd;
         4'h1912 	:	val_out <= 4'hc9dd;
         4'h1913 	:	val_out <= 4'hc9dd;
         4'h1918 	:	val_out <= 4'hc9f1;
         4'h1919 	:	val_out <= 4'hc9f1;
         4'h191a 	:	val_out <= 4'hc9f1;
         4'h191b 	:	val_out <= 4'hc9f1;
         4'h1920 	:	val_out <= 4'hca06;
         4'h1921 	:	val_out <= 4'hca06;
         4'h1922 	:	val_out <= 4'hca06;
         4'h1923 	:	val_out <= 4'hca06;
         4'h1928 	:	val_out <= 4'hca1a;
         4'h1929 	:	val_out <= 4'hca1a;
         4'h192a 	:	val_out <= 4'hca1a;
         4'h192b 	:	val_out <= 4'hca1a;
         4'h1930 	:	val_out <= 4'hca2f;
         4'h1931 	:	val_out <= 4'hca2f;
         4'h1932 	:	val_out <= 4'hca2f;
         4'h1933 	:	val_out <= 4'hca2f;
         4'h1938 	:	val_out <= 4'hca43;
         4'h1939 	:	val_out <= 4'hca43;
         4'h193a 	:	val_out <= 4'hca43;
         4'h193b 	:	val_out <= 4'hca43;
         4'h1940 	:	val_out <= 4'hca58;
         4'h1941 	:	val_out <= 4'hca58;
         4'h1942 	:	val_out <= 4'hca58;
         4'h1943 	:	val_out <= 4'hca58;
         4'h1948 	:	val_out <= 4'hca6c;
         4'h1949 	:	val_out <= 4'hca6c;
         4'h194a 	:	val_out <= 4'hca6c;
         4'h194b 	:	val_out <= 4'hca6c;
         4'h1950 	:	val_out <= 4'hca81;
         4'h1951 	:	val_out <= 4'hca81;
         4'h1952 	:	val_out <= 4'hca81;
         4'h1953 	:	val_out <= 4'hca81;
         4'h1958 	:	val_out <= 4'hca95;
         4'h1959 	:	val_out <= 4'hca95;
         4'h195a 	:	val_out <= 4'hca95;
         4'h195b 	:	val_out <= 4'hca95;
         4'h1960 	:	val_out <= 4'hcaa9;
         4'h1961 	:	val_out <= 4'hcaa9;
         4'h1962 	:	val_out <= 4'hcaa9;
         4'h1963 	:	val_out <= 4'hcaa9;
         4'h1968 	:	val_out <= 4'hcabe;
         4'h1969 	:	val_out <= 4'hcabe;
         4'h196a 	:	val_out <= 4'hcabe;
         4'h196b 	:	val_out <= 4'hcabe;
         4'h1970 	:	val_out <= 4'hcad2;
         4'h1971 	:	val_out <= 4'hcad2;
         4'h1972 	:	val_out <= 4'hcad2;
         4'h1973 	:	val_out <= 4'hcad2;
         4'h1978 	:	val_out <= 4'hcae7;
         4'h1979 	:	val_out <= 4'hcae7;
         4'h197a 	:	val_out <= 4'hcae7;
         4'h197b 	:	val_out <= 4'hcae7;
         4'h1980 	:	val_out <= 4'hcafb;
         4'h1981 	:	val_out <= 4'hcafb;
         4'h1982 	:	val_out <= 4'hcafb;
         4'h1983 	:	val_out <= 4'hcafb;
         4'h1988 	:	val_out <= 4'hcb0f;
         4'h1989 	:	val_out <= 4'hcb0f;
         4'h198a 	:	val_out <= 4'hcb0f;
         4'h198b 	:	val_out <= 4'hcb0f;
         4'h1990 	:	val_out <= 4'hcb24;
         4'h1991 	:	val_out <= 4'hcb24;
         4'h1992 	:	val_out <= 4'hcb24;
         4'h1993 	:	val_out <= 4'hcb24;
         4'h1998 	:	val_out <= 4'hcb38;
         4'h1999 	:	val_out <= 4'hcb38;
         4'h199a 	:	val_out <= 4'hcb38;
         4'h199b 	:	val_out <= 4'hcb38;
         4'h19a0 	:	val_out <= 4'hcb4c;
         4'h19a1 	:	val_out <= 4'hcb4c;
         4'h19a2 	:	val_out <= 4'hcb4c;
         4'h19a3 	:	val_out <= 4'hcb4c;
         4'h19a8 	:	val_out <= 4'hcb61;
         4'h19a9 	:	val_out <= 4'hcb61;
         4'h19aa 	:	val_out <= 4'hcb61;
         4'h19ab 	:	val_out <= 4'hcb61;
         4'h19b0 	:	val_out <= 4'hcb75;
         4'h19b1 	:	val_out <= 4'hcb75;
         4'h19b2 	:	val_out <= 4'hcb75;
         4'h19b3 	:	val_out <= 4'hcb75;
         4'h19b8 	:	val_out <= 4'hcb89;
         4'h19b9 	:	val_out <= 4'hcb89;
         4'h19ba 	:	val_out <= 4'hcb89;
         4'h19bb 	:	val_out <= 4'hcb89;
         4'h19c0 	:	val_out <= 4'hcb9e;
         4'h19c1 	:	val_out <= 4'hcb9e;
         4'h19c2 	:	val_out <= 4'hcb9e;
         4'h19c3 	:	val_out <= 4'hcb9e;
         4'h19c8 	:	val_out <= 4'hcbb2;
         4'h19c9 	:	val_out <= 4'hcbb2;
         4'h19ca 	:	val_out <= 4'hcbb2;
         4'h19cb 	:	val_out <= 4'hcbb2;
         4'h19d0 	:	val_out <= 4'hcbc6;
         4'h19d1 	:	val_out <= 4'hcbc6;
         4'h19d2 	:	val_out <= 4'hcbc6;
         4'h19d3 	:	val_out <= 4'hcbc6;
         4'h19d8 	:	val_out <= 4'hcbda;
         4'h19d9 	:	val_out <= 4'hcbda;
         4'h19da 	:	val_out <= 4'hcbda;
         4'h19db 	:	val_out <= 4'hcbda;
         4'h19e0 	:	val_out <= 4'hcbef;
         4'h19e1 	:	val_out <= 4'hcbef;
         4'h19e2 	:	val_out <= 4'hcbef;
         4'h19e3 	:	val_out <= 4'hcbef;
         4'h19e8 	:	val_out <= 4'hcc03;
         4'h19e9 	:	val_out <= 4'hcc03;
         4'h19ea 	:	val_out <= 4'hcc03;
         4'h19eb 	:	val_out <= 4'hcc03;
         4'h19f0 	:	val_out <= 4'hcc17;
         4'h19f1 	:	val_out <= 4'hcc17;
         4'h19f2 	:	val_out <= 4'hcc17;
         4'h19f3 	:	val_out <= 4'hcc17;
         4'h19f8 	:	val_out <= 4'hcc2b;
         4'h19f9 	:	val_out <= 4'hcc2b;
         4'h19fa 	:	val_out <= 4'hcc2b;
         4'h19fb 	:	val_out <= 4'hcc2b;
         4'h1a00 	:	val_out <= 4'hcc3f;
         4'h1a01 	:	val_out <= 4'hcc3f;
         4'h1a02 	:	val_out <= 4'hcc3f;
         4'h1a03 	:	val_out <= 4'hcc3f;
         4'h1a08 	:	val_out <= 4'hcc54;
         4'h1a09 	:	val_out <= 4'hcc54;
         4'h1a0a 	:	val_out <= 4'hcc54;
         4'h1a0b 	:	val_out <= 4'hcc54;
         4'h1a10 	:	val_out <= 4'hcc68;
         4'h1a11 	:	val_out <= 4'hcc68;
         4'h1a12 	:	val_out <= 4'hcc68;
         4'h1a13 	:	val_out <= 4'hcc68;
         4'h1a18 	:	val_out <= 4'hcc7c;
         4'h1a19 	:	val_out <= 4'hcc7c;
         4'h1a1a 	:	val_out <= 4'hcc7c;
         4'h1a1b 	:	val_out <= 4'hcc7c;
         4'h1a20 	:	val_out <= 4'hcc90;
         4'h1a21 	:	val_out <= 4'hcc90;
         4'h1a22 	:	val_out <= 4'hcc90;
         4'h1a23 	:	val_out <= 4'hcc90;
         4'h1a28 	:	val_out <= 4'hcca4;
         4'h1a29 	:	val_out <= 4'hcca4;
         4'h1a2a 	:	val_out <= 4'hcca4;
         4'h1a2b 	:	val_out <= 4'hcca4;
         4'h1a30 	:	val_out <= 4'hccb8;
         4'h1a31 	:	val_out <= 4'hccb8;
         4'h1a32 	:	val_out <= 4'hccb8;
         4'h1a33 	:	val_out <= 4'hccb8;
         4'h1a38 	:	val_out <= 4'hcccc;
         4'h1a39 	:	val_out <= 4'hcccc;
         4'h1a3a 	:	val_out <= 4'hcccc;
         4'h1a3b 	:	val_out <= 4'hcccc;
         4'h1a40 	:	val_out <= 4'hcce1;
         4'h1a41 	:	val_out <= 4'hcce1;
         4'h1a42 	:	val_out <= 4'hcce1;
         4'h1a43 	:	val_out <= 4'hcce1;
         4'h1a48 	:	val_out <= 4'hccf5;
         4'h1a49 	:	val_out <= 4'hccf5;
         4'h1a4a 	:	val_out <= 4'hccf5;
         4'h1a4b 	:	val_out <= 4'hccf5;
         4'h1a50 	:	val_out <= 4'hcd09;
         4'h1a51 	:	val_out <= 4'hcd09;
         4'h1a52 	:	val_out <= 4'hcd09;
         4'h1a53 	:	val_out <= 4'hcd09;
         4'h1a58 	:	val_out <= 4'hcd1d;
         4'h1a59 	:	val_out <= 4'hcd1d;
         4'h1a5a 	:	val_out <= 4'hcd1d;
         4'h1a5b 	:	val_out <= 4'hcd1d;
         4'h1a60 	:	val_out <= 4'hcd31;
         4'h1a61 	:	val_out <= 4'hcd31;
         4'h1a62 	:	val_out <= 4'hcd31;
         4'h1a63 	:	val_out <= 4'hcd31;
         4'h1a68 	:	val_out <= 4'hcd45;
         4'h1a69 	:	val_out <= 4'hcd45;
         4'h1a6a 	:	val_out <= 4'hcd45;
         4'h1a6b 	:	val_out <= 4'hcd45;
         4'h1a70 	:	val_out <= 4'hcd59;
         4'h1a71 	:	val_out <= 4'hcd59;
         4'h1a72 	:	val_out <= 4'hcd59;
         4'h1a73 	:	val_out <= 4'hcd59;
         4'h1a78 	:	val_out <= 4'hcd6d;
         4'h1a79 	:	val_out <= 4'hcd6d;
         4'h1a7a 	:	val_out <= 4'hcd6d;
         4'h1a7b 	:	val_out <= 4'hcd6d;
         4'h1a80 	:	val_out <= 4'hcd81;
         4'h1a81 	:	val_out <= 4'hcd81;
         4'h1a82 	:	val_out <= 4'hcd81;
         4'h1a83 	:	val_out <= 4'hcd81;
         4'h1a88 	:	val_out <= 4'hcd95;
         4'h1a89 	:	val_out <= 4'hcd95;
         4'h1a8a 	:	val_out <= 4'hcd95;
         4'h1a8b 	:	val_out <= 4'hcd95;
         4'h1a90 	:	val_out <= 4'hcda9;
         4'h1a91 	:	val_out <= 4'hcda9;
         4'h1a92 	:	val_out <= 4'hcda9;
         4'h1a93 	:	val_out <= 4'hcda9;
         4'h1a98 	:	val_out <= 4'hcdbd;
         4'h1a99 	:	val_out <= 4'hcdbd;
         4'h1a9a 	:	val_out <= 4'hcdbd;
         4'h1a9b 	:	val_out <= 4'hcdbd;
         4'h1aa0 	:	val_out <= 4'hcdd1;
         4'h1aa1 	:	val_out <= 4'hcdd1;
         4'h1aa2 	:	val_out <= 4'hcdd1;
         4'h1aa3 	:	val_out <= 4'hcdd1;
         4'h1aa8 	:	val_out <= 4'hcde5;
         4'h1aa9 	:	val_out <= 4'hcde5;
         4'h1aaa 	:	val_out <= 4'hcde5;
         4'h1aab 	:	val_out <= 4'hcde5;
         4'h1ab0 	:	val_out <= 4'hcdf9;
         4'h1ab1 	:	val_out <= 4'hcdf9;
         4'h1ab2 	:	val_out <= 4'hcdf9;
         4'h1ab3 	:	val_out <= 4'hcdf9;
         4'h1ab8 	:	val_out <= 4'hce0d;
         4'h1ab9 	:	val_out <= 4'hce0d;
         4'h1aba 	:	val_out <= 4'hce0d;
         4'h1abb 	:	val_out <= 4'hce0d;
         4'h1ac0 	:	val_out <= 4'hce21;
         4'h1ac1 	:	val_out <= 4'hce21;
         4'h1ac2 	:	val_out <= 4'hce21;
         4'h1ac3 	:	val_out <= 4'hce21;
         4'h1ac8 	:	val_out <= 4'hce34;
         4'h1ac9 	:	val_out <= 4'hce34;
         4'h1aca 	:	val_out <= 4'hce34;
         4'h1acb 	:	val_out <= 4'hce34;
         4'h1ad0 	:	val_out <= 4'hce48;
         4'h1ad1 	:	val_out <= 4'hce48;
         4'h1ad2 	:	val_out <= 4'hce48;
         4'h1ad3 	:	val_out <= 4'hce48;
         4'h1ad8 	:	val_out <= 4'hce5c;
         4'h1ad9 	:	val_out <= 4'hce5c;
         4'h1ada 	:	val_out <= 4'hce5c;
         4'h1adb 	:	val_out <= 4'hce5c;
         4'h1ae0 	:	val_out <= 4'hce70;
         4'h1ae1 	:	val_out <= 4'hce70;
         4'h1ae2 	:	val_out <= 4'hce70;
         4'h1ae3 	:	val_out <= 4'hce70;
         4'h1ae8 	:	val_out <= 4'hce84;
         4'h1ae9 	:	val_out <= 4'hce84;
         4'h1aea 	:	val_out <= 4'hce84;
         4'h1aeb 	:	val_out <= 4'hce84;
         4'h1af0 	:	val_out <= 4'hce98;
         4'h1af1 	:	val_out <= 4'hce98;
         4'h1af2 	:	val_out <= 4'hce98;
         4'h1af3 	:	val_out <= 4'hce98;
         4'h1af8 	:	val_out <= 4'hceac;
         4'h1af9 	:	val_out <= 4'hceac;
         4'h1afa 	:	val_out <= 4'hceac;
         4'h1afb 	:	val_out <= 4'hceac;
         4'h1b00 	:	val_out <= 4'hcebf;
         4'h1b01 	:	val_out <= 4'hcebf;
         4'h1b02 	:	val_out <= 4'hcebf;
         4'h1b03 	:	val_out <= 4'hcebf;
         4'h1b08 	:	val_out <= 4'hced3;
         4'h1b09 	:	val_out <= 4'hced3;
         4'h1b0a 	:	val_out <= 4'hced3;
         4'h1b0b 	:	val_out <= 4'hced3;
         4'h1b10 	:	val_out <= 4'hcee7;
         4'h1b11 	:	val_out <= 4'hcee7;
         4'h1b12 	:	val_out <= 4'hcee7;
         4'h1b13 	:	val_out <= 4'hcee7;
         4'h1b18 	:	val_out <= 4'hcefb;
         4'h1b19 	:	val_out <= 4'hcefb;
         4'h1b1a 	:	val_out <= 4'hcefb;
         4'h1b1b 	:	val_out <= 4'hcefb;
         4'h1b20 	:	val_out <= 4'hcf0f;
         4'h1b21 	:	val_out <= 4'hcf0f;
         4'h1b22 	:	val_out <= 4'hcf0f;
         4'h1b23 	:	val_out <= 4'hcf0f;
         4'h1b28 	:	val_out <= 4'hcf22;
         4'h1b29 	:	val_out <= 4'hcf22;
         4'h1b2a 	:	val_out <= 4'hcf22;
         4'h1b2b 	:	val_out <= 4'hcf22;
         4'h1b30 	:	val_out <= 4'hcf36;
         4'h1b31 	:	val_out <= 4'hcf36;
         4'h1b32 	:	val_out <= 4'hcf36;
         4'h1b33 	:	val_out <= 4'hcf36;
         4'h1b38 	:	val_out <= 4'hcf4a;
         4'h1b39 	:	val_out <= 4'hcf4a;
         4'h1b3a 	:	val_out <= 4'hcf4a;
         4'h1b3b 	:	val_out <= 4'hcf4a;
         4'h1b40 	:	val_out <= 4'hcf5e;
         4'h1b41 	:	val_out <= 4'hcf5e;
         4'h1b42 	:	val_out <= 4'hcf5e;
         4'h1b43 	:	val_out <= 4'hcf5e;
         4'h1b48 	:	val_out <= 4'hcf71;
         4'h1b49 	:	val_out <= 4'hcf71;
         4'h1b4a 	:	val_out <= 4'hcf71;
         4'h1b4b 	:	val_out <= 4'hcf71;
         4'h1b50 	:	val_out <= 4'hcf85;
         4'h1b51 	:	val_out <= 4'hcf85;
         4'h1b52 	:	val_out <= 4'hcf85;
         4'h1b53 	:	val_out <= 4'hcf85;
         4'h1b58 	:	val_out <= 4'hcf99;
         4'h1b59 	:	val_out <= 4'hcf99;
         4'h1b5a 	:	val_out <= 4'hcf99;
         4'h1b5b 	:	val_out <= 4'hcf99;
         4'h1b60 	:	val_out <= 4'hcfac;
         4'h1b61 	:	val_out <= 4'hcfac;
         4'h1b62 	:	val_out <= 4'hcfac;
         4'h1b63 	:	val_out <= 4'hcfac;
         4'h1b68 	:	val_out <= 4'hcfc0;
         4'h1b69 	:	val_out <= 4'hcfc0;
         4'h1b6a 	:	val_out <= 4'hcfc0;
         4'h1b6b 	:	val_out <= 4'hcfc0;
         4'h1b70 	:	val_out <= 4'hcfd4;
         4'h1b71 	:	val_out <= 4'hcfd4;
         4'h1b72 	:	val_out <= 4'hcfd4;
         4'h1b73 	:	val_out <= 4'hcfd4;
         4'h1b78 	:	val_out <= 4'hcfe7;
         4'h1b79 	:	val_out <= 4'hcfe7;
         4'h1b7a 	:	val_out <= 4'hcfe7;
         4'h1b7b 	:	val_out <= 4'hcfe7;
         4'h1b80 	:	val_out <= 4'hcffb;
         4'h1b81 	:	val_out <= 4'hcffb;
         4'h1b82 	:	val_out <= 4'hcffb;
         4'h1b83 	:	val_out <= 4'hcffb;
         4'h1b88 	:	val_out <= 4'hd00f;
         4'h1b89 	:	val_out <= 4'hd00f;
         4'h1b8a 	:	val_out <= 4'hd00f;
         4'h1b8b 	:	val_out <= 4'hd00f;
         4'h1b90 	:	val_out <= 4'hd022;
         4'h1b91 	:	val_out <= 4'hd022;
         4'h1b92 	:	val_out <= 4'hd022;
         4'h1b93 	:	val_out <= 4'hd022;
         4'h1b98 	:	val_out <= 4'hd036;
         4'h1b99 	:	val_out <= 4'hd036;
         4'h1b9a 	:	val_out <= 4'hd036;
         4'h1b9b 	:	val_out <= 4'hd036;
         4'h1ba0 	:	val_out <= 4'hd049;
         4'h1ba1 	:	val_out <= 4'hd049;
         4'h1ba2 	:	val_out <= 4'hd049;
         4'h1ba3 	:	val_out <= 4'hd049;
         4'h1ba8 	:	val_out <= 4'hd05d;
         4'h1ba9 	:	val_out <= 4'hd05d;
         4'h1baa 	:	val_out <= 4'hd05d;
         4'h1bab 	:	val_out <= 4'hd05d;
         4'h1bb0 	:	val_out <= 4'hd070;
         4'h1bb1 	:	val_out <= 4'hd070;
         4'h1bb2 	:	val_out <= 4'hd070;
         4'h1bb3 	:	val_out <= 4'hd070;
         4'h1bb8 	:	val_out <= 4'hd084;
         4'h1bb9 	:	val_out <= 4'hd084;
         4'h1bba 	:	val_out <= 4'hd084;
         4'h1bbb 	:	val_out <= 4'hd084;
         4'h1bc0 	:	val_out <= 4'hd097;
         4'h1bc1 	:	val_out <= 4'hd097;
         4'h1bc2 	:	val_out <= 4'hd097;
         4'h1bc3 	:	val_out <= 4'hd097;
         4'h1bc8 	:	val_out <= 4'hd0ab;
         4'h1bc9 	:	val_out <= 4'hd0ab;
         4'h1bca 	:	val_out <= 4'hd0ab;
         4'h1bcb 	:	val_out <= 4'hd0ab;
         4'h1bd0 	:	val_out <= 4'hd0bf;
         4'h1bd1 	:	val_out <= 4'hd0bf;
         4'h1bd2 	:	val_out <= 4'hd0bf;
         4'h1bd3 	:	val_out <= 4'hd0bf;
         4'h1bd8 	:	val_out <= 4'hd0d2;
         4'h1bd9 	:	val_out <= 4'hd0d2;
         4'h1bda 	:	val_out <= 4'hd0d2;
         4'h1bdb 	:	val_out <= 4'hd0d2;
         4'h1be0 	:	val_out <= 4'hd0e5;
         4'h1be1 	:	val_out <= 4'hd0e5;
         4'h1be2 	:	val_out <= 4'hd0e5;
         4'h1be3 	:	val_out <= 4'hd0e5;
         4'h1be8 	:	val_out <= 4'hd0f9;
         4'h1be9 	:	val_out <= 4'hd0f9;
         4'h1bea 	:	val_out <= 4'hd0f9;
         4'h1beb 	:	val_out <= 4'hd0f9;
         4'h1bf0 	:	val_out <= 4'hd10c;
         4'h1bf1 	:	val_out <= 4'hd10c;
         4'h1bf2 	:	val_out <= 4'hd10c;
         4'h1bf3 	:	val_out <= 4'hd10c;
         4'h1bf8 	:	val_out <= 4'hd120;
         4'h1bf9 	:	val_out <= 4'hd120;
         4'h1bfa 	:	val_out <= 4'hd120;
         4'h1bfb 	:	val_out <= 4'hd120;
         4'h1c00 	:	val_out <= 4'hd133;
         4'h1c01 	:	val_out <= 4'hd133;
         4'h1c02 	:	val_out <= 4'hd133;
         4'h1c03 	:	val_out <= 4'hd133;
         4'h1c08 	:	val_out <= 4'hd147;
         4'h1c09 	:	val_out <= 4'hd147;
         4'h1c0a 	:	val_out <= 4'hd147;
         4'h1c0b 	:	val_out <= 4'hd147;
         4'h1c10 	:	val_out <= 4'hd15a;
         4'h1c11 	:	val_out <= 4'hd15a;
         4'h1c12 	:	val_out <= 4'hd15a;
         4'h1c13 	:	val_out <= 4'hd15a;
         4'h1c18 	:	val_out <= 4'hd16e;
         4'h1c19 	:	val_out <= 4'hd16e;
         4'h1c1a 	:	val_out <= 4'hd16e;
         4'h1c1b 	:	val_out <= 4'hd16e;
         4'h1c20 	:	val_out <= 4'hd181;
         4'h1c21 	:	val_out <= 4'hd181;
         4'h1c22 	:	val_out <= 4'hd181;
         4'h1c23 	:	val_out <= 4'hd181;
         4'h1c28 	:	val_out <= 4'hd194;
         4'h1c29 	:	val_out <= 4'hd194;
         4'h1c2a 	:	val_out <= 4'hd194;
         4'h1c2b 	:	val_out <= 4'hd194;
         4'h1c30 	:	val_out <= 4'hd1a8;
         4'h1c31 	:	val_out <= 4'hd1a8;
         4'h1c32 	:	val_out <= 4'hd1a8;
         4'h1c33 	:	val_out <= 4'hd1a8;
         4'h1c38 	:	val_out <= 4'hd1bb;
         4'h1c39 	:	val_out <= 4'hd1bb;
         4'h1c3a 	:	val_out <= 4'hd1bb;
         4'h1c3b 	:	val_out <= 4'hd1bb;
         4'h1c40 	:	val_out <= 4'hd1ce;
         4'h1c41 	:	val_out <= 4'hd1ce;
         4'h1c42 	:	val_out <= 4'hd1ce;
         4'h1c43 	:	val_out <= 4'hd1ce;
         4'h1c48 	:	val_out <= 4'hd1e2;
         4'h1c49 	:	val_out <= 4'hd1e2;
         4'h1c4a 	:	val_out <= 4'hd1e2;
         4'h1c4b 	:	val_out <= 4'hd1e2;
         4'h1c50 	:	val_out <= 4'hd1f5;
         4'h1c51 	:	val_out <= 4'hd1f5;
         4'h1c52 	:	val_out <= 4'hd1f5;
         4'h1c53 	:	val_out <= 4'hd1f5;
         4'h1c58 	:	val_out <= 4'hd208;
         4'h1c59 	:	val_out <= 4'hd208;
         4'h1c5a 	:	val_out <= 4'hd208;
         4'h1c5b 	:	val_out <= 4'hd208;
         4'h1c60 	:	val_out <= 4'hd21c;
         4'h1c61 	:	val_out <= 4'hd21c;
         4'h1c62 	:	val_out <= 4'hd21c;
         4'h1c63 	:	val_out <= 4'hd21c;
         4'h1c68 	:	val_out <= 4'hd22f;
         4'h1c69 	:	val_out <= 4'hd22f;
         4'h1c6a 	:	val_out <= 4'hd22f;
         4'h1c6b 	:	val_out <= 4'hd22f;
         4'h1c70 	:	val_out <= 4'hd242;
         4'h1c71 	:	val_out <= 4'hd242;
         4'h1c72 	:	val_out <= 4'hd242;
         4'h1c73 	:	val_out <= 4'hd242;
         4'h1c78 	:	val_out <= 4'hd255;
         4'h1c79 	:	val_out <= 4'hd255;
         4'h1c7a 	:	val_out <= 4'hd255;
         4'h1c7b 	:	val_out <= 4'hd255;
         4'h1c80 	:	val_out <= 4'hd269;
         4'h1c81 	:	val_out <= 4'hd269;
         4'h1c82 	:	val_out <= 4'hd269;
         4'h1c83 	:	val_out <= 4'hd269;
         4'h1c88 	:	val_out <= 4'hd27c;
         4'h1c89 	:	val_out <= 4'hd27c;
         4'h1c8a 	:	val_out <= 4'hd27c;
         4'h1c8b 	:	val_out <= 4'hd27c;
         4'h1c90 	:	val_out <= 4'hd28f;
         4'h1c91 	:	val_out <= 4'hd28f;
         4'h1c92 	:	val_out <= 4'hd28f;
         4'h1c93 	:	val_out <= 4'hd28f;
         4'h1c98 	:	val_out <= 4'hd2a2;
         4'h1c99 	:	val_out <= 4'hd2a2;
         4'h1c9a 	:	val_out <= 4'hd2a2;
         4'h1c9b 	:	val_out <= 4'hd2a2;
         4'h1ca0 	:	val_out <= 4'hd2b5;
         4'h1ca1 	:	val_out <= 4'hd2b5;
         4'h1ca2 	:	val_out <= 4'hd2b5;
         4'h1ca3 	:	val_out <= 4'hd2b5;
         4'h1ca8 	:	val_out <= 4'hd2c9;
         4'h1ca9 	:	val_out <= 4'hd2c9;
         4'h1caa 	:	val_out <= 4'hd2c9;
         4'h1cab 	:	val_out <= 4'hd2c9;
         4'h1cb0 	:	val_out <= 4'hd2dc;
         4'h1cb1 	:	val_out <= 4'hd2dc;
         4'h1cb2 	:	val_out <= 4'hd2dc;
         4'h1cb3 	:	val_out <= 4'hd2dc;
         4'h1cb8 	:	val_out <= 4'hd2ef;
         4'h1cb9 	:	val_out <= 4'hd2ef;
         4'h1cba 	:	val_out <= 4'hd2ef;
         4'h1cbb 	:	val_out <= 4'hd2ef;
         4'h1cc0 	:	val_out <= 4'hd302;
         4'h1cc1 	:	val_out <= 4'hd302;
         4'h1cc2 	:	val_out <= 4'hd302;
         4'h1cc3 	:	val_out <= 4'hd302;
         4'h1cc8 	:	val_out <= 4'hd315;
         4'h1cc9 	:	val_out <= 4'hd315;
         4'h1cca 	:	val_out <= 4'hd315;
         4'h1ccb 	:	val_out <= 4'hd315;
         4'h1cd0 	:	val_out <= 4'hd328;
         4'h1cd1 	:	val_out <= 4'hd328;
         4'h1cd2 	:	val_out <= 4'hd328;
         4'h1cd3 	:	val_out <= 4'hd328;
         4'h1cd8 	:	val_out <= 4'hd33b;
         4'h1cd9 	:	val_out <= 4'hd33b;
         4'h1cda 	:	val_out <= 4'hd33b;
         4'h1cdb 	:	val_out <= 4'hd33b;
         4'h1ce0 	:	val_out <= 4'hd34e;
         4'h1ce1 	:	val_out <= 4'hd34e;
         4'h1ce2 	:	val_out <= 4'hd34e;
         4'h1ce3 	:	val_out <= 4'hd34e;
         4'h1ce8 	:	val_out <= 4'hd362;
         4'h1ce9 	:	val_out <= 4'hd362;
         4'h1cea 	:	val_out <= 4'hd362;
         4'h1ceb 	:	val_out <= 4'hd362;
         4'h1cf0 	:	val_out <= 4'hd375;
         4'h1cf1 	:	val_out <= 4'hd375;
         4'h1cf2 	:	val_out <= 4'hd375;
         4'h1cf3 	:	val_out <= 4'hd375;
         4'h1cf8 	:	val_out <= 4'hd388;
         4'h1cf9 	:	val_out <= 4'hd388;
         4'h1cfa 	:	val_out <= 4'hd388;
         4'h1cfb 	:	val_out <= 4'hd388;
         4'h1d00 	:	val_out <= 4'hd39b;
         4'h1d01 	:	val_out <= 4'hd39b;
         4'h1d02 	:	val_out <= 4'hd39b;
         4'h1d03 	:	val_out <= 4'hd39b;
         4'h1d08 	:	val_out <= 4'hd3ae;
         4'h1d09 	:	val_out <= 4'hd3ae;
         4'h1d0a 	:	val_out <= 4'hd3ae;
         4'h1d0b 	:	val_out <= 4'hd3ae;
         4'h1d10 	:	val_out <= 4'hd3c1;
         4'h1d11 	:	val_out <= 4'hd3c1;
         4'h1d12 	:	val_out <= 4'hd3c1;
         4'h1d13 	:	val_out <= 4'hd3c1;
         4'h1d18 	:	val_out <= 4'hd3d4;
         4'h1d19 	:	val_out <= 4'hd3d4;
         4'h1d1a 	:	val_out <= 4'hd3d4;
         4'h1d1b 	:	val_out <= 4'hd3d4;
         4'h1d20 	:	val_out <= 4'hd3e7;
         4'h1d21 	:	val_out <= 4'hd3e7;
         4'h1d22 	:	val_out <= 4'hd3e7;
         4'h1d23 	:	val_out <= 4'hd3e7;
         4'h1d28 	:	val_out <= 4'hd3fa;
         4'h1d29 	:	val_out <= 4'hd3fa;
         4'h1d2a 	:	val_out <= 4'hd3fa;
         4'h1d2b 	:	val_out <= 4'hd3fa;
         4'h1d30 	:	val_out <= 4'hd40d;
         4'h1d31 	:	val_out <= 4'hd40d;
         4'h1d32 	:	val_out <= 4'hd40d;
         4'h1d33 	:	val_out <= 4'hd40d;
         4'h1d38 	:	val_out <= 4'hd420;
         4'h1d39 	:	val_out <= 4'hd420;
         4'h1d3a 	:	val_out <= 4'hd420;
         4'h1d3b 	:	val_out <= 4'hd420;
         4'h1d40 	:	val_out <= 4'hd433;
         4'h1d41 	:	val_out <= 4'hd433;
         4'h1d42 	:	val_out <= 4'hd433;
         4'h1d43 	:	val_out <= 4'hd433;
         4'h1d48 	:	val_out <= 4'hd445;
         4'h1d49 	:	val_out <= 4'hd445;
         4'h1d4a 	:	val_out <= 4'hd445;
         4'h1d4b 	:	val_out <= 4'hd445;
         4'h1d50 	:	val_out <= 4'hd458;
         4'h1d51 	:	val_out <= 4'hd458;
         4'h1d52 	:	val_out <= 4'hd458;
         4'h1d53 	:	val_out <= 4'hd458;
         4'h1d58 	:	val_out <= 4'hd46b;
         4'h1d59 	:	val_out <= 4'hd46b;
         4'h1d5a 	:	val_out <= 4'hd46b;
         4'h1d5b 	:	val_out <= 4'hd46b;
         4'h1d60 	:	val_out <= 4'hd47e;
         4'h1d61 	:	val_out <= 4'hd47e;
         4'h1d62 	:	val_out <= 4'hd47e;
         4'h1d63 	:	val_out <= 4'hd47e;
         4'h1d68 	:	val_out <= 4'hd491;
         4'h1d69 	:	val_out <= 4'hd491;
         4'h1d6a 	:	val_out <= 4'hd491;
         4'h1d6b 	:	val_out <= 4'hd491;
         4'h1d70 	:	val_out <= 4'hd4a4;
         4'h1d71 	:	val_out <= 4'hd4a4;
         4'h1d72 	:	val_out <= 4'hd4a4;
         4'h1d73 	:	val_out <= 4'hd4a4;
         4'h1d78 	:	val_out <= 4'hd4b7;
         4'h1d79 	:	val_out <= 4'hd4b7;
         4'h1d7a 	:	val_out <= 4'hd4b7;
         4'h1d7b 	:	val_out <= 4'hd4b7;
         4'h1d80 	:	val_out <= 4'hd4ca;
         4'h1d81 	:	val_out <= 4'hd4ca;
         4'h1d82 	:	val_out <= 4'hd4ca;
         4'h1d83 	:	val_out <= 4'hd4ca;
         4'h1d88 	:	val_out <= 4'hd4dc;
         4'h1d89 	:	val_out <= 4'hd4dc;
         4'h1d8a 	:	val_out <= 4'hd4dc;
         4'h1d8b 	:	val_out <= 4'hd4dc;
         4'h1d90 	:	val_out <= 4'hd4ef;
         4'h1d91 	:	val_out <= 4'hd4ef;
         4'h1d92 	:	val_out <= 4'hd4ef;
         4'h1d93 	:	val_out <= 4'hd4ef;
         4'h1d98 	:	val_out <= 4'hd502;
         4'h1d99 	:	val_out <= 4'hd502;
         4'h1d9a 	:	val_out <= 4'hd502;
         4'h1d9b 	:	val_out <= 4'hd502;
         4'h1da0 	:	val_out <= 4'hd515;
         4'h1da1 	:	val_out <= 4'hd515;
         4'h1da2 	:	val_out <= 4'hd515;
         4'h1da3 	:	val_out <= 4'hd515;
         4'h1da8 	:	val_out <= 4'hd528;
         4'h1da9 	:	val_out <= 4'hd528;
         4'h1daa 	:	val_out <= 4'hd528;
         4'h1dab 	:	val_out <= 4'hd528;
         4'h1db0 	:	val_out <= 4'hd53a;
         4'h1db1 	:	val_out <= 4'hd53a;
         4'h1db2 	:	val_out <= 4'hd53a;
         4'h1db3 	:	val_out <= 4'hd53a;
         4'h1db8 	:	val_out <= 4'hd54d;
         4'h1db9 	:	val_out <= 4'hd54d;
         4'h1dba 	:	val_out <= 4'hd54d;
         4'h1dbb 	:	val_out <= 4'hd54d;
         4'h1dc0 	:	val_out <= 4'hd560;
         4'h1dc1 	:	val_out <= 4'hd560;
         4'h1dc2 	:	val_out <= 4'hd560;
         4'h1dc3 	:	val_out <= 4'hd560;
         4'h1dc8 	:	val_out <= 4'hd572;
         4'h1dc9 	:	val_out <= 4'hd572;
         4'h1dca 	:	val_out <= 4'hd572;
         4'h1dcb 	:	val_out <= 4'hd572;
         4'h1dd0 	:	val_out <= 4'hd585;
         4'h1dd1 	:	val_out <= 4'hd585;
         4'h1dd2 	:	val_out <= 4'hd585;
         4'h1dd3 	:	val_out <= 4'hd585;
         4'h1dd8 	:	val_out <= 4'hd598;
         4'h1dd9 	:	val_out <= 4'hd598;
         4'h1dda 	:	val_out <= 4'hd598;
         4'h1ddb 	:	val_out <= 4'hd598;
         4'h1de0 	:	val_out <= 4'hd5ab;
         4'h1de1 	:	val_out <= 4'hd5ab;
         4'h1de2 	:	val_out <= 4'hd5ab;
         4'h1de3 	:	val_out <= 4'hd5ab;
         4'h1de8 	:	val_out <= 4'hd5bd;
         4'h1de9 	:	val_out <= 4'hd5bd;
         4'h1dea 	:	val_out <= 4'hd5bd;
         4'h1deb 	:	val_out <= 4'hd5bd;
         4'h1df0 	:	val_out <= 4'hd5d0;
         4'h1df1 	:	val_out <= 4'hd5d0;
         4'h1df2 	:	val_out <= 4'hd5d0;
         4'h1df3 	:	val_out <= 4'hd5d0;
         4'h1df8 	:	val_out <= 4'hd5e3;
         4'h1df9 	:	val_out <= 4'hd5e3;
         4'h1dfa 	:	val_out <= 4'hd5e3;
         4'h1dfb 	:	val_out <= 4'hd5e3;
         4'h1e00 	:	val_out <= 4'hd5f5;
         4'h1e01 	:	val_out <= 4'hd5f5;
         4'h1e02 	:	val_out <= 4'hd5f5;
         4'h1e03 	:	val_out <= 4'hd5f5;
         4'h1e08 	:	val_out <= 4'hd608;
         4'h1e09 	:	val_out <= 4'hd608;
         4'h1e0a 	:	val_out <= 4'hd608;
         4'h1e0b 	:	val_out <= 4'hd608;
         4'h1e10 	:	val_out <= 4'hd61a;
         4'h1e11 	:	val_out <= 4'hd61a;
         4'h1e12 	:	val_out <= 4'hd61a;
         4'h1e13 	:	val_out <= 4'hd61a;
         4'h1e18 	:	val_out <= 4'hd62d;
         4'h1e19 	:	val_out <= 4'hd62d;
         4'h1e1a 	:	val_out <= 4'hd62d;
         4'h1e1b 	:	val_out <= 4'hd62d;
         4'h1e20 	:	val_out <= 4'hd640;
         4'h1e21 	:	val_out <= 4'hd640;
         4'h1e22 	:	val_out <= 4'hd640;
         4'h1e23 	:	val_out <= 4'hd640;
         4'h1e28 	:	val_out <= 4'hd652;
         4'h1e29 	:	val_out <= 4'hd652;
         4'h1e2a 	:	val_out <= 4'hd652;
         4'h1e2b 	:	val_out <= 4'hd652;
         4'h1e30 	:	val_out <= 4'hd665;
         4'h1e31 	:	val_out <= 4'hd665;
         4'h1e32 	:	val_out <= 4'hd665;
         4'h1e33 	:	val_out <= 4'hd665;
         4'h1e38 	:	val_out <= 4'hd677;
         4'h1e39 	:	val_out <= 4'hd677;
         4'h1e3a 	:	val_out <= 4'hd677;
         4'h1e3b 	:	val_out <= 4'hd677;
         4'h1e40 	:	val_out <= 4'hd68a;
         4'h1e41 	:	val_out <= 4'hd68a;
         4'h1e42 	:	val_out <= 4'hd68a;
         4'h1e43 	:	val_out <= 4'hd68a;
         4'h1e48 	:	val_out <= 4'hd69c;
         4'h1e49 	:	val_out <= 4'hd69c;
         4'h1e4a 	:	val_out <= 4'hd69c;
         4'h1e4b 	:	val_out <= 4'hd69c;
         4'h1e50 	:	val_out <= 4'hd6af;
         4'h1e51 	:	val_out <= 4'hd6af;
         4'h1e52 	:	val_out <= 4'hd6af;
         4'h1e53 	:	val_out <= 4'hd6af;
         4'h1e58 	:	val_out <= 4'hd6c1;
         4'h1e59 	:	val_out <= 4'hd6c1;
         4'h1e5a 	:	val_out <= 4'hd6c1;
         4'h1e5b 	:	val_out <= 4'hd6c1;
         4'h1e60 	:	val_out <= 4'hd6d4;
         4'h1e61 	:	val_out <= 4'hd6d4;
         4'h1e62 	:	val_out <= 4'hd6d4;
         4'h1e63 	:	val_out <= 4'hd6d4;
         4'h1e68 	:	val_out <= 4'hd6e6;
         4'h1e69 	:	val_out <= 4'hd6e6;
         4'h1e6a 	:	val_out <= 4'hd6e6;
         4'h1e6b 	:	val_out <= 4'hd6e6;
         4'h1e70 	:	val_out <= 4'hd6f9;
         4'h1e71 	:	val_out <= 4'hd6f9;
         4'h1e72 	:	val_out <= 4'hd6f9;
         4'h1e73 	:	val_out <= 4'hd6f9;
         4'h1e78 	:	val_out <= 4'hd70b;
         4'h1e79 	:	val_out <= 4'hd70b;
         4'h1e7a 	:	val_out <= 4'hd70b;
         4'h1e7b 	:	val_out <= 4'hd70b;
         4'h1e80 	:	val_out <= 4'hd71d;
         4'h1e81 	:	val_out <= 4'hd71d;
         4'h1e82 	:	val_out <= 4'hd71d;
         4'h1e83 	:	val_out <= 4'hd71d;
         4'h1e88 	:	val_out <= 4'hd730;
         4'h1e89 	:	val_out <= 4'hd730;
         4'h1e8a 	:	val_out <= 4'hd730;
         4'h1e8b 	:	val_out <= 4'hd730;
         4'h1e90 	:	val_out <= 4'hd742;
         4'h1e91 	:	val_out <= 4'hd742;
         4'h1e92 	:	val_out <= 4'hd742;
         4'h1e93 	:	val_out <= 4'hd742;
         4'h1e98 	:	val_out <= 4'hd755;
         4'h1e99 	:	val_out <= 4'hd755;
         4'h1e9a 	:	val_out <= 4'hd755;
         4'h1e9b 	:	val_out <= 4'hd755;
         4'h1ea0 	:	val_out <= 4'hd767;
         4'h1ea1 	:	val_out <= 4'hd767;
         4'h1ea2 	:	val_out <= 4'hd767;
         4'h1ea3 	:	val_out <= 4'hd767;
         4'h1ea8 	:	val_out <= 4'hd779;
         4'h1ea9 	:	val_out <= 4'hd779;
         4'h1eaa 	:	val_out <= 4'hd779;
         4'h1eab 	:	val_out <= 4'hd779;
         4'h1eb0 	:	val_out <= 4'hd78c;
         4'h1eb1 	:	val_out <= 4'hd78c;
         4'h1eb2 	:	val_out <= 4'hd78c;
         4'h1eb3 	:	val_out <= 4'hd78c;
         4'h1eb8 	:	val_out <= 4'hd79e;
         4'h1eb9 	:	val_out <= 4'hd79e;
         4'h1eba 	:	val_out <= 4'hd79e;
         4'h1ebb 	:	val_out <= 4'hd79e;
         4'h1ec0 	:	val_out <= 4'hd7b0;
         4'h1ec1 	:	val_out <= 4'hd7b0;
         4'h1ec2 	:	val_out <= 4'hd7b0;
         4'h1ec3 	:	val_out <= 4'hd7b0;
         4'h1ec8 	:	val_out <= 4'hd7c3;
         4'h1ec9 	:	val_out <= 4'hd7c3;
         4'h1eca 	:	val_out <= 4'hd7c3;
         4'h1ecb 	:	val_out <= 4'hd7c3;
         4'h1ed0 	:	val_out <= 4'hd7d5;
         4'h1ed1 	:	val_out <= 4'hd7d5;
         4'h1ed2 	:	val_out <= 4'hd7d5;
         4'h1ed3 	:	val_out <= 4'hd7d5;
         4'h1ed8 	:	val_out <= 4'hd7e7;
         4'h1ed9 	:	val_out <= 4'hd7e7;
         4'h1eda 	:	val_out <= 4'hd7e7;
         4'h1edb 	:	val_out <= 4'hd7e7;
         4'h1ee0 	:	val_out <= 4'hd7f9;
         4'h1ee1 	:	val_out <= 4'hd7f9;
         4'h1ee2 	:	val_out <= 4'hd7f9;
         4'h1ee3 	:	val_out <= 4'hd7f9;
         4'h1ee8 	:	val_out <= 4'hd80c;
         4'h1ee9 	:	val_out <= 4'hd80c;
         4'h1eea 	:	val_out <= 4'hd80c;
         4'h1eeb 	:	val_out <= 4'hd80c;
         4'h1ef0 	:	val_out <= 4'hd81e;
         4'h1ef1 	:	val_out <= 4'hd81e;
         4'h1ef2 	:	val_out <= 4'hd81e;
         4'h1ef3 	:	val_out <= 4'hd81e;
         4'h1ef8 	:	val_out <= 4'hd830;
         4'h1ef9 	:	val_out <= 4'hd830;
         4'h1efa 	:	val_out <= 4'hd830;
         4'h1efb 	:	val_out <= 4'hd830;
         4'h1f00 	:	val_out <= 4'hd842;
         4'h1f01 	:	val_out <= 4'hd842;
         4'h1f02 	:	val_out <= 4'hd842;
         4'h1f03 	:	val_out <= 4'hd842;
         4'h1f08 	:	val_out <= 4'hd855;
         4'h1f09 	:	val_out <= 4'hd855;
         4'h1f0a 	:	val_out <= 4'hd855;
         4'h1f0b 	:	val_out <= 4'hd855;
         4'h1f10 	:	val_out <= 4'hd867;
         4'h1f11 	:	val_out <= 4'hd867;
         4'h1f12 	:	val_out <= 4'hd867;
         4'h1f13 	:	val_out <= 4'hd867;
         4'h1f18 	:	val_out <= 4'hd879;
         4'h1f19 	:	val_out <= 4'hd879;
         4'h1f1a 	:	val_out <= 4'hd879;
         4'h1f1b 	:	val_out <= 4'hd879;
         4'h1f20 	:	val_out <= 4'hd88b;
         4'h1f21 	:	val_out <= 4'hd88b;
         4'h1f22 	:	val_out <= 4'hd88b;
         4'h1f23 	:	val_out <= 4'hd88b;
         4'h1f28 	:	val_out <= 4'hd89d;
         4'h1f29 	:	val_out <= 4'hd89d;
         4'h1f2a 	:	val_out <= 4'hd89d;
         4'h1f2b 	:	val_out <= 4'hd89d;
         4'h1f30 	:	val_out <= 4'hd8af;
         4'h1f31 	:	val_out <= 4'hd8af;
         4'h1f32 	:	val_out <= 4'hd8af;
         4'h1f33 	:	val_out <= 4'hd8af;
         4'h1f38 	:	val_out <= 4'hd8c1;
         4'h1f39 	:	val_out <= 4'hd8c1;
         4'h1f3a 	:	val_out <= 4'hd8c1;
         4'h1f3b 	:	val_out <= 4'hd8c1;
         4'h1f40 	:	val_out <= 4'hd8d4;
         4'h1f41 	:	val_out <= 4'hd8d4;
         4'h1f42 	:	val_out <= 4'hd8d4;
         4'h1f43 	:	val_out <= 4'hd8d4;
         4'h1f48 	:	val_out <= 4'hd8e6;
         4'h1f49 	:	val_out <= 4'hd8e6;
         4'h1f4a 	:	val_out <= 4'hd8e6;
         4'h1f4b 	:	val_out <= 4'hd8e6;
         4'h1f50 	:	val_out <= 4'hd8f8;
         4'h1f51 	:	val_out <= 4'hd8f8;
         4'h1f52 	:	val_out <= 4'hd8f8;
         4'h1f53 	:	val_out <= 4'hd8f8;
         4'h1f58 	:	val_out <= 4'hd90a;
         4'h1f59 	:	val_out <= 4'hd90a;
         4'h1f5a 	:	val_out <= 4'hd90a;
         4'h1f5b 	:	val_out <= 4'hd90a;
         4'h1f60 	:	val_out <= 4'hd91c;
         4'h1f61 	:	val_out <= 4'hd91c;
         4'h1f62 	:	val_out <= 4'hd91c;
         4'h1f63 	:	val_out <= 4'hd91c;
         4'h1f68 	:	val_out <= 4'hd92e;
         4'h1f69 	:	val_out <= 4'hd92e;
         4'h1f6a 	:	val_out <= 4'hd92e;
         4'h1f6b 	:	val_out <= 4'hd92e;
         4'h1f70 	:	val_out <= 4'hd940;
         4'h1f71 	:	val_out <= 4'hd940;
         4'h1f72 	:	val_out <= 4'hd940;
         4'h1f73 	:	val_out <= 4'hd940;
         4'h1f78 	:	val_out <= 4'hd952;
         4'h1f79 	:	val_out <= 4'hd952;
         4'h1f7a 	:	val_out <= 4'hd952;
         4'h1f7b 	:	val_out <= 4'hd952;
         4'h1f80 	:	val_out <= 4'hd964;
         4'h1f81 	:	val_out <= 4'hd964;
         4'h1f82 	:	val_out <= 4'hd964;
         4'h1f83 	:	val_out <= 4'hd964;
         4'h1f88 	:	val_out <= 4'hd976;
         4'h1f89 	:	val_out <= 4'hd976;
         4'h1f8a 	:	val_out <= 4'hd976;
         4'h1f8b 	:	val_out <= 4'hd976;
         4'h1f90 	:	val_out <= 4'hd988;
         4'h1f91 	:	val_out <= 4'hd988;
         4'h1f92 	:	val_out <= 4'hd988;
         4'h1f93 	:	val_out <= 4'hd988;
         4'h1f98 	:	val_out <= 4'hd99a;
         4'h1f99 	:	val_out <= 4'hd99a;
         4'h1f9a 	:	val_out <= 4'hd99a;
         4'h1f9b 	:	val_out <= 4'hd99a;
         4'h1fa0 	:	val_out <= 4'hd9ac;
         4'h1fa1 	:	val_out <= 4'hd9ac;
         4'h1fa2 	:	val_out <= 4'hd9ac;
         4'h1fa3 	:	val_out <= 4'hd9ac;
         4'h1fa8 	:	val_out <= 4'hd9be;
         4'h1fa9 	:	val_out <= 4'hd9be;
         4'h1faa 	:	val_out <= 4'hd9be;
         4'h1fab 	:	val_out <= 4'hd9be;
         4'h1fb0 	:	val_out <= 4'hd9d0;
         4'h1fb1 	:	val_out <= 4'hd9d0;
         4'h1fb2 	:	val_out <= 4'hd9d0;
         4'h1fb3 	:	val_out <= 4'hd9d0;
         4'h1fb8 	:	val_out <= 4'hd9e1;
         4'h1fb9 	:	val_out <= 4'hd9e1;
         4'h1fba 	:	val_out <= 4'hd9e1;
         4'h1fbb 	:	val_out <= 4'hd9e1;
         4'h1fc0 	:	val_out <= 4'hd9f3;
         4'h1fc1 	:	val_out <= 4'hd9f3;
         4'h1fc2 	:	val_out <= 4'hd9f3;
         4'h1fc3 	:	val_out <= 4'hd9f3;
         4'h1fc8 	:	val_out <= 4'hda05;
         4'h1fc9 	:	val_out <= 4'hda05;
         4'h1fca 	:	val_out <= 4'hda05;
         4'h1fcb 	:	val_out <= 4'hda05;
         4'h1fd0 	:	val_out <= 4'hda17;
         4'h1fd1 	:	val_out <= 4'hda17;
         4'h1fd2 	:	val_out <= 4'hda17;
         4'h1fd3 	:	val_out <= 4'hda17;
         4'h1fd8 	:	val_out <= 4'hda29;
         4'h1fd9 	:	val_out <= 4'hda29;
         4'h1fda 	:	val_out <= 4'hda29;
         4'h1fdb 	:	val_out <= 4'hda29;
         4'h1fe0 	:	val_out <= 4'hda3b;
         4'h1fe1 	:	val_out <= 4'hda3b;
         4'h1fe2 	:	val_out <= 4'hda3b;
         4'h1fe3 	:	val_out <= 4'hda3b;
         4'h1fe8 	:	val_out <= 4'hda4d;
         4'h1fe9 	:	val_out <= 4'hda4d;
         4'h1fea 	:	val_out <= 4'hda4d;
         4'h1feb 	:	val_out <= 4'hda4d;
         4'h1ff0 	:	val_out <= 4'hda5e;
         4'h1ff1 	:	val_out <= 4'hda5e;
         4'h1ff2 	:	val_out <= 4'hda5e;
         4'h1ff3 	:	val_out <= 4'hda5e;
         4'h1ff8 	:	val_out <= 4'hda70;
         4'h1ff9 	:	val_out <= 4'hda70;
         4'h1ffa 	:	val_out <= 4'hda70;
         4'h1ffb 	:	val_out <= 4'hda70;
         4'h2000 	:	val_out <= 4'hda82;
         4'h2001 	:	val_out <= 4'hda82;
         4'h2002 	:	val_out <= 4'hda82;
         4'h2003 	:	val_out <= 4'hda82;
         4'h2008 	:	val_out <= 4'hda94;
         4'h2009 	:	val_out <= 4'hda94;
         4'h200a 	:	val_out <= 4'hda94;
         4'h200b 	:	val_out <= 4'hda94;
         4'h2010 	:	val_out <= 4'hdaa5;
         4'h2011 	:	val_out <= 4'hdaa5;
         4'h2012 	:	val_out <= 4'hdaa5;
         4'h2013 	:	val_out <= 4'hdaa5;
         4'h2018 	:	val_out <= 4'hdab7;
         4'h2019 	:	val_out <= 4'hdab7;
         4'h201a 	:	val_out <= 4'hdab7;
         4'h201b 	:	val_out <= 4'hdab7;
         4'h2020 	:	val_out <= 4'hdac9;
         4'h2021 	:	val_out <= 4'hdac9;
         4'h2022 	:	val_out <= 4'hdac9;
         4'h2023 	:	val_out <= 4'hdac9;
         4'h2028 	:	val_out <= 4'hdadb;
         4'h2029 	:	val_out <= 4'hdadb;
         4'h202a 	:	val_out <= 4'hdadb;
         4'h202b 	:	val_out <= 4'hdadb;
         4'h2030 	:	val_out <= 4'hdaec;
         4'h2031 	:	val_out <= 4'hdaec;
         4'h2032 	:	val_out <= 4'hdaec;
         4'h2033 	:	val_out <= 4'hdaec;
         4'h2038 	:	val_out <= 4'hdafe;
         4'h2039 	:	val_out <= 4'hdafe;
         4'h203a 	:	val_out <= 4'hdafe;
         4'h203b 	:	val_out <= 4'hdafe;
         4'h2040 	:	val_out <= 4'hdb10;
         4'h2041 	:	val_out <= 4'hdb10;
         4'h2042 	:	val_out <= 4'hdb10;
         4'h2043 	:	val_out <= 4'hdb10;
         4'h2048 	:	val_out <= 4'hdb21;
         4'h2049 	:	val_out <= 4'hdb21;
         4'h204a 	:	val_out <= 4'hdb21;
         4'h204b 	:	val_out <= 4'hdb21;
         4'h2050 	:	val_out <= 4'hdb33;
         4'h2051 	:	val_out <= 4'hdb33;
         4'h2052 	:	val_out <= 4'hdb33;
         4'h2053 	:	val_out <= 4'hdb33;
         4'h2058 	:	val_out <= 4'hdb45;
         4'h2059 	:	val_out <= 4'hdb45;
         4'h205a 	:	val_out <= 4'hdb45;
         4'h205b 	:	val_out <= 4'hdb45;
         4'h2060 	:	val_out <= 4'hdb56;
         4'h2061 	:	val_out <= 4'hdb56;
         4'h2062 	:	val_out <= 4'hdb56;
         4'h2063 	:	val_out <= 4'hdb56;
         4'h2068 	:	val_out <= 4'hdb68;
         4'h2069 	:	val_out <= 4'hdb68;
         4'h206a 	:	val_out <= 4'hdb68;
         4'h206b 	:	val_out <= 4'hdb68;
         4'h2070 	:	val_out <= 4'hdb79;
         4'h2071 	:	val_out <= 4'hdb79;
         4'h2072 	:	val_out <= 4'hdb79;
         4'h2073 	:	val_out <= 4'hdb79;
         4'h2078 	:	val_out <= 4'hdb8b;
         4'h2079 	:	val_out <= 4'hdb8b;
         4'h207a 	:	val_out <= 4'hdb8b;
         4'h207b 	:	val_out <= 4'hdb8b;
         4'h2080 	:	val_out <= 4'hdb9d;
         4'h2081 	:	val_out <= 4'hdb9d;
         4'h2082 	:	val_out <= 4'hdb9d;
         4'h2083 	:	val_out <= 4'hdb9d;
         4'h2088 	:	val_out <= 4'hdbae;
         4'h2089 	:	val_out <= 4'hdbae;
         4'h208a 	:	val_out <= 4'hdbae;
         4'h208b 	:	val_out <= 4'hdbae;
         4'h2090 	:	val_out <= 4'hdbc0;
         4'h2091 	:	val_out <= 4'hdbc0;
         4'h2092 	:	val_out <= 4'hdbc0;
         4'h2093 	:	val_out <= 4'hdbc0;
         4'h2098 	:	val_out <= 4'hdbd1;
         4'h2099 	:	val_out <= 4'hdbd1;
         4'h209a 	:	val_out <= 4'hdbd1;
         4'h209b 	:	val_out <= 4'hdbd1;
         4'h20a0 	:	val_out <= 4'hdbe3;
         4'h20a1 	:	val_out <= 4'hdbe3;
         4'h20a2 	:	val_out <= 4'hdbe3;
         4'h20a3 	:	val_out <= 4'hdbe3;
         4'h20a8 	:	val_out <= 4'hdbf4;
         4'h20a9 	:	val_out <= 4'hdbf4;
         4'h20aa 	:	val_out <= 4'hdbf4;
         4'h20ab 	:	val_out <= 4'hdbf4;
         4'h20b0 	:	val_out <= 4'hdc06;
         4'h20b1 	:	val_out <= 4'hdc06;
         4'h20b2 	:	val_out <= 4'hdc06;
         4'h20b3 	:	val_out <= 4'hdc06;
         4'h20b8 	:	val_out <= 4'hdc17;
         4'h20b9 	:	val_out <= 4'hdc17;
         4'h20ba 	:	val_out <= 4'hdc17;
         4'h20bb 	:	val_out <= 4'hdc17;
         4'h20c0 	:	val_out <= 4'hdc29;
         4'h20c1 	:	val_out <= 4'hdc29;
         4'h20c2 	:	val_out <= 4'hdc29;
         4'h20c3 	:	val_out <= 4'hdc29;
         4'h20c8 	:	val_out <= 4'hdc3a;
         4'h20c9 	:	val_out <= 4'hdc3a;
         4'h20ca 	:	val_out <= 4'hdc3a;
         4'h20cb 	:	val_out <= 4'hdc3a;
         4'h20d0 	:	val_out <= 4'hdc4b;
         4'h20d1 	:	val_out <= 4'hdc4b;
         4'h20d2 	:	val_out <= 4'hdc4b;
         4'h20d3 	:	val_out <= 4'hdc4b;
         4'h20d8 	:	val_out <= 4'hdc5d;
         4'h20d9 	:	val_out <= 4'hdc5d;
         4'h20da 	:	val_out <= 4'hdc5d;
         4'h20db 	:	val_out <= 4'hdc5d;
         4'h20e0 	:	val_out <= 4'hdc6e;
         4'h20e1 	:	val_out <= 4'hdc6e;
         4'h20e2 	:	val_out <= 4'hdc6e;
         4'h20e3 	:	val_out <= 4'hdc6e;
         4'h20e8 	:	val_out <= 4'hdc80;
         4'h20e9 	:	val_out <= 4'hdc80;
         4'h20ea 	:	val_out <= 4'hdc80;
         4'h20eb 	:	val_out <= 4'hdc80;
         4'h20f0 	:	val_out <= 4'hdc91;
         4'h20f1 	:	val_out <= 4'hdc91;
         4'h20f2 	:	val_out <= 4'hdc91;
         4'h20f3 	:	val_out <= 4'hdc91;
         4'h20f8 	:	val_out <= 4'hdca2;
         4'h20f9 	:	val_out <= 4'hdca2;
         4'h20fa 	:	val_out <= 4'hdca2;
         4'h20fb 	:	val_out <= 4'hdca2;
         4'h2100 	:	val_out <= 4'hdcb4;
         4'h2101 	:	val_out <= 4'hdcb4;
         4'h2102 	:	val_out <= 4'hdcb4;
         4'h2103 	:	val_out <= 4'hdcb4;
         4'h2108 	:	val_out <= 4'hdcc5;
         4'h2109 	:	val_out <= 4'hdcc5;
         4'h210a 	:	val_out <= 4'hdcc5;
         4'h210b 	:	val_out <= 4'hdcc5;
         4'h2110 	:	val_out <= 4'hdcd6;
         4'h2111 	:	val_out <= 4'hdcd6;
         4'h2112 	:	val_out <= 4'hdcd6;
         4'h2113 	:	val_out <= 4'hdcd6;
         4'h2118 	:	val_out <= 4'hdce8;
         4'h2119 	:	val_out <= 4'hdce8;
         4'h211a 	:	val_out <= 4'hdce8;
         4'h211b 	:	val_out <= 4'hdce8;
         4'h2120 	:	val_out <= 4'hdcf9;
         4'h2121 	:	val_out <= 4'hdcf9;
         4'h2122 	:	val_out <= 4'hdcf9;
         4'h2123 	:	val_out <= 4'hdcf9;
         4'h2128 	:	val_out <= 4'hdd0a;
         4'h2129 	:	val_out <= 4'hdd0a;
         4'h212a 	:	val_out <= 4'hdd0a;
         4'h212b 	:	val_out <= 4'hdd0a;
         4'h2130 	:	val_out <= 4'hdd1b;
         4'h2131 	:	val_out <= 4'hdd1b;
         4'h2132 	:	val_out <= 4'hdd1b;
         4'h2133 	:	val_out <= 4'hdd1b;
         4'h2138 	:	val_out <= 4'hdd2d;
         4'h2139 	:	val_out <= 4'hdd2d;
         4'h213a 	:	val_out <= 4'hdd2d;
         4'h213b 	:	val_out <= 4'hdd2d;
         4'h2140 	:	val_out <= 4'hdd3e;
         4'h2141 	:	val_out <= 4'hdd3e;
         4'h2142 	:	val_out <= 4'hdd3e;
         4'h2143 	:	val_out <= 4'hdd3e;
         4'h2148 	:	val_out <= 4'hdd4f;
         4'h2149 	:	val_out <= 4'hdd4f;
         4'h214a 	:	val_out <= 4'hdd4f;
         4'h214b 	:	val_out <= 4'hdd4f;
         4'h2150 	:	val_out <= 4'hdd60;
         4'h2151 	:	val_out <= 4'hdd60;
         4'h2152 	:	val_out <= 4'hdd60;
         4'h2153 	:	val_out <= 4'hdd60;
         4'h2158 	:	val_out <= 4'hdd71;
         4'h2159 	:	val_out <= 4'hdd71;
         4'h215a 	:	val_out <= 4'hdd71;
         4'h215b 	:	val_out <= 4'hdd71;
         4'h2160 	:	val_out <= 4'hdd83;
         4'h2161 	:	val_out <= 4'hdd83;
         4'h2162 	:	val_out <= 4'hdd83;
         4'h2163 	:	val_out <= 4'hdd83;
         4'h2168 	:	val_out <= 4'hdd94;
         4'h2169 	:	val_out <= 4'hdd94;
         4'h216a 	:	val_out <= 4'hdd94;
         4'h216b 	:	val_out <= 4'hdd94;
         4'h2170 	:	val_out <= 4'hdda5;
         4'h2171 	:	val_out <= 4'hdda5;
         4'h2172 	:	val_out <= 4'hdda5;
         4'h2173 	:	val_out <= 4'hdda5;
         4'h2178 	:	val_out <= 4'hddb6;
         4'h2179 	:	val_out <= 4'hddb6;
         4'h217a 	:	val_out <= 4'hddb6;
         4'h217b 	:	val_out <= 4'hddb6;
         4'h2180 	:	val_out <= 4'hddc7;
         4'h2181 	:	val_out <= 4'hddc7;
         4'h2182 	:	val_out <= 4'hddc7;
         4'h2183 	:	val_out <= 4'hddc7;
         4'h2188 	:	val_out <= 4'hddd8;
         4'h2189 	:	val_out <= 4'hddd8;
         4'h218a 	:	val_out <= 4'hddd8;
         4'h218b 	:	val_out <= 4'hddd8;
         4'h2190 	:	val_out <= 4'hdde9;
         4'h2191 	:	val_out <= 4'hdde9;
         4'h2192 	:	val_out <= 4'hdde9;
         4'h2193 	:	val_out <= 4'hdde9;
         4'h2198 	:	val_out <= 4'hddfa;
         4'h2199 	:	val_out <= 4'hddfa;
         4'h219a 	:	val_out <= 4'hddfa;
         4'h219b 	:	val_out <= 4'hddfa;
         4'h21a0 	:	val_out <= 4'hde0b;
         4'h21a1 	:	val_out <= 4'hde0b;
         4'h21a2 	:	val_out <= 4'hde0b;
         4'h21a3 	:	val_out <= 4'hde0b;
         4'h21a8 	:	val_out <= 4'hde1c;
         4'h21a9 	:	val_out <= 4'hde1c;
         4'h21aa 	:	val_out <= 4'hde1c;
         4'h21ab 	:	val_out <= 4'hde1c;
         4'h21b0 	:	val_out <= 4'hde2d;
         4'h21b1 	:	val_out <= 4'hde2d;
         4'h21b2 	:	val_out <= 4'hde2d;
         4'h21b3 	:	val_out <= 4'hde2d;
         4'h21b8 	:	val_out <= 4'hde3f;
         4'h21b9 	:	val_out <= 4'hde3f;
         4'h21ba 	:	val_out <= 4'hde3f;
         4'h21bb 	:	val_out <= 4'hde3f;
         4'h21c0 	:	val_out <= 4'hde50;
         4'h21c1 	:	val_out <= 4'hde50;
         4'h21c2 	:	val_out <= 4'hde50;
         4'h21c3 	:	val_out <= 4'hde50;
         4'h21c8 	:	val_out <= 4'hde60;
         4'h21c9 	:	val_out <= 4'hde60;
         4'h21ca 	:	val_out <= 4'hde60;
         4'h21cb 	:	val_out <= 4'hde60;
         4'h21d0 	:	val_out <= 4'hde71;
         4'h21d1 	:	val_out <= 4'hde71;
         4'h21d2 	:	val_out <= 4'hde71;
         4'h21d3 	:	val_out <= 4'hde71;
         4'h21d8 	:	val_out <= 4'hde82;
         4'h21d9 	:	val_out <= 4'hde82;
         4'h21da 	:	val_out <= 4'hde82;
         4'h21db 	:	val_out <= 4'hde82;
         4'h21e0 	:	val_out <= 4'hde93;
         4'h21e1 	:	val_out <= 4'hde93;
         4'h21e2 	:	val_out <= 4'hde93;
         4'h21e3 	:	val_out <= 4'hde93;
         4'h21e8 	:	val_out <= 4'hdea4;
         4'h21e9 	:	val_out <= 4'hdea4;
         4'h21ea 	:	val_out <= 4'hdea4;
         4'h21eb 	:	val_out <= 4'hdea4;
         4'h21f0 	:	val_out <= 4'hdeb5;
         4'h21f1 	:	val_out <= 4'hdeb5;
         4'h21f2 	:	val_out <= 4'hdeb5;
         4'h21f3 	:	val_out <= 4'hdeb5;
         4'h21f8 	:	val_out <= 4'hdec6;
         4'h21f9 	:	val_out <= 4'hdec6;
         4'h21fa 	:	val_out <= 4'hdec6;
         4'h21fb 	:	val_out <= 4'hdec6;
         4'h2200 	:	val_out <= 4'hded7;
         4'h2201 	:	val_out <= 4'hded7;
         4'h2202 	:	val_out <= 4'hded7;
         4'h2203 	:	val_out <= 4'hded7;
         4'h2208 	:	val_out <= 4'hdee8;
         4'h2209 	:	val_out <= 4'hdee8;
         4'h220a 	:	val_out <= 4'hdee8;
         4'h220b 	:	val_out <= 4'hdee8;
         4'h2210 	:	val_out <= 4'hdef9;
         4'h2211 	:	val_out <= 4'hdef9;
         4'h2212 	:	val_out <= 4'hdef9;
         4'h2213 	:	val_out <= 4'hdef9;
         4'h2218 	:	val_out <= 4'hdf0a;
         4'h2219 	:	val_out <= 4'hdf0a;
         4'h221a 	:	val_out <= 4'hdf0a;
         4'h221b 	:	val_out <= 4'hdf0a;
         4'h2220 	:	val_out <= 4'hdf1a;
         4'h2221 	:	val_out <= 4'hdf1a;
         4'h2222 	:	val_out <= 4'hdf1a;
         4'h2223 	:	val_out <= 4'hdf1a;
         4'h2228 	:	val_out <= 4'hdf2b;
         4'h2229 	:	val_out <= 4'hdf2b;
         4'h222a 	:	val_out <= 4'hdf2b;
         4'h222b 	:	val_out <= 4'hdf2b;
         4'h2230 	:	val_out <= 4'hdf3c;
         4'h2231 	:	val_out <= 4'hdf3c;
         4'h2232 	:	val_out <= 4'hdf3c;
         4'h2233 	:	val_out <= 4'hdf3c;
         4'h2238 	:	val_out <= 4'hdf4d;
         4'h2239 	:	val_out <= 4'hdf4d;
         4'h223a 	:	val_out <= 4'hdf4d;
         4'h223b 	:	val_out <= 4'hdf4d;
         4'h2240 	:	val_out <= 4'hdf5e;
         4'h2241 	:	val_out <= 4'hdf5e;
         4'h2242 	:	val_out <= 4'hdf5e;
         4'h2243 	:	val_out <= 4'hdf5e;
         4'h2248 	:	val_out <= 4'hdf6e;
         4'h2249 	:	val_out <= 4'hdf6e;
         4'h224a 	:	val_out <= 4'hdf6e;
         4'h224b 	:	val_out <= 4'hdf6e;
         4'h2250 	:	val_out <= 4'hdf7f;
         4'h2251 	:	val_out <= 4'hdf7f;
         4'h2252 	:	val_out <= 4'hdf7f;
         4'h2253 	:	val_out <= 4'hdf7f;
         4'h2258 	:	val_out <= 4'hdf90;
         4'h2259 	:	val_out <= 4'hdf90;
         4'h225a 	:	val_out <= 4'hdf90;
         4'h225b 	:	val_out <= 4'hdf90;
         4'h2260 	:	val_out <= 4'hdfa0;
         4'h2261 	:	val_out <= 4'hdfa0;
         4'h2262 	:	val_out <= 4'hdfa0;
         4'h2263 	:	val_out <= 4'hdfa0;
         4'h2268 	:	val_out <= 4'hdfb1;
         4'h2269 	:	val_out <= 4'hdfb1;
         4'h226a 	:	val_out <= 4'hdfb1;
         4'h226b 	:	val_out <= 4'hdfb1;
         4'h2270 	:	val_out <= 4'hdfc2;
         4'h2271 	:	val_out <= 4'hdfc2;
         4'h2272 	:	val_out <= 4'hdfc2;
         4'h2273 	:	val_out <= 4'hdfc2;
         4'h2278 	:	val_out <= 4'hdfd3;
         4'h2279 	:	val_out <= 4'hdfd3;
         4'h227a 	:	val_out <= 4'hdfd3;
         4'h227b 	:	val_out <= 4'hdfd3;
         4'h2280 	:	val_out <= 4'hdfe3;
         4'h2281 	:	val_out <= 4'hdfe3;
         4'h2282 	:	val_out <= 4'hdfe3;
         4'h2283 	:	val_out <= 4'hdfe3;
         4'h2288 	:	val_out <= 4'hdff4;
         4'h2289 	:	val_out <= 4'hdff4;
         4'h228a 	:	val_out <= 4'hdff4;
         4'h228b 	:	val_out <= 4'hdff4;
         4'h2290 	:	val_out <= 4'he004;
         4'h2291 	:	val_out <= 4'he004;
         4'h2292 	:	val_out <= 4'he004;
         4'h2293 	:	val_out <= 4'he004;
         4'h2298 	:	val_out <= 4'he015;
         4'h2299 	:	val_out <= 4'he015;
         4'h229a 	:	val_out <= 4'he015;
         4'h229b 	:	val_out <= 4'he015;
         4'h22a0 	:	val_out <= 4'he026;
         4'h22a1 	:	val_out <= 4'he026;
         4'h22a2 	:	val_out <= 4'he026;
         4'h22a3 	:	val_out <= 4'he026;
         4'h22a8 	:	val_out <= 4'he036;
         4'h22a9 	:	val_out <= 4'he036;
         4'h22aa 	:	val_out <= 4'he036;
         4'h22ab 	:	val_out <= 4'he036;
         4'h22b0 	:	val_out <= 4'he047;
         4'h22b1 	:	val_out <= 4'he047;
         4'h22b2 	:	val_out <= 4'he047;
         4'h22b3 	:	val_out <= 4'he047;
         4'h22b8 	:	val_out <= 4'he057;
         4'h22b9 	:	val_out <= 4'he057;
         4'h22ba 	:	val_out <= 4'he057;
         4'h22bb 	:	val_out <= 4'he057;
         4'h22c0 	:	val_out <= 4'he068;
         4'h22c1 	:	val_out <= 4'he068;
         4'h22c2 	:	val_out <= 4'he068;
         4'h22c3 	:	val_out <= 4'he068;
         4'h22c8 	:	val_out <= 4'he078;
         4'h22c9 	:	val_out <= 4'he078;
         4'h22ca 	:	val_out <= 4'he078;
         4'h22cb 	:	val_out <= 4'he078;
         4'h22d0 	:	val_out <= 4'he089;
         4'h22d1 	:	val_out <= 4'he089;
         4'h22d2 	:	val_out <= 4'he089;
         4'h22d3 	:	val_out <= 4'he089;
         4'h22d8 	:	val_out <= 4'he099;
         4'h22d9 	:	val_out <= 4'he099;
         4'h22da 	:	val_out <= 4'he099;
         4'h22db 	:	val_out <= 4'he099;
         4'h22e0 	:	val_out <= 4'he0aa;
         4'h22e1 	:	val_out <= 4'he0aa;
         4'h22e2 	:	val_out <= 4'he0aa;
         4'h22e3 	:	val_out <= 4'he0aa;
         4'h22e8 	:	val_out <= 4'he0ba;
         4'h22e9 	:	val_out <= 4'he0ba;
         4'h22ea 	:	val_out <= 4'he0ba;
         4'h22eb 	:	val_out <= 4'he0ba;
         4'h22f0 	:	val_out <= 4'he0cb;
         4'h22f1 	:	val_out <= 4'he0cb;
         4'h22f2 	:	val_out <= 4'he0cb;
         4'h22f3 	:	val_out <= 4'he0cb;
         4'h22f8 	:	val_out <= 4'he0db;
         4'h22f9 	:	val_out <= 4'he0db;
         4'h22fa 	:	val_out <= 4'he0db;
         4'h22fb 	:	val_out <= 4'he0db;
         4'h2300 	:	val_out <= 4'he0ec;
         4'h2301 	:	val_out <= 4'he0ec;
         4'h2302 	:	val_out <= 4'he0ec;
         4'h2303 	:	val_out <= 4'he0ec;
         4'h2308 	:	val_out <= 4'he0fc;
         4'h2309 	:	val_out <= 4'he0fc;
         4'h230a 	:	val_out <= 4'he0fc;
         4'h230b 	:	val_out <= 4'he0fc;
         4'h2310 	:	val_out <= 4'he10d;
         4'h2311 	:	val_out <= 4'he10d;
         4'h2312 	:	val_out <= 4'he10d;
         4'h2313 	:	val_out <= 4'he10d;
         4'h2318 	:	val_out <= 4'he11d;
         4'h2319 	:	val_out <= 4'he11d;
         4'h231a 	:	val_out <= 4'he11d;
         4'h231b 	:	val_out <= 4'he11d;
         4'h2320 	:	val_out <= 4'he12d;
         4'h2321 	:	val_out <= 4'he12d;
         4'h2322 	:	val_out <= 4'he12d;
         4'h2323 	:	val_out <= 4'he12d;
         4'h2328 	:	val_out <= 4'he13e;
         4'h2329 	:	val_out <= 4'he13e;
         4'h232a 	:	val_out <= 4'he13e;
         4'h232b 	:	val_out <= 4'he13e;
         4'h2330 	:	val_out <= 4'he14e;
         4'h2331 	:	val_out <= 4'he14e;
         4'h2332 	:	val_out <= 4'he14e;
         4'h2333 	:	val_out <= 4'he14e;
         4'h2338 	:	val_out <= 4'he15e;
         4'h2339 	:	val_out <= 4'he15e;
         4'h233a 	:	val_out <= 4'he15e;
         4'h233b 	:	val_out <= 4'he15e;
         4'h2340 	:	val_out <= 4'he16f;
         4'h2341 	:	val_out <= 4'he16f;
         4'h2342 	:	val_out <= 4'he16f;
         4'h2343 	:	val_out <= 4'he16f;
         4'h2348 	:	val_out <= 4'he17f;
         4'h2349 	:	val_out <= 4'he17f;
         4'h234a 	:	val_out <= 4'he17f;
         4'h234b 	:	val_out <= 4'he17f;
         4'h2350 	:	val_out <= 4'he18f;
         4'h2351 	:	val_out <= 4'he18f;
         4'h2352 	:	val_out <= 4'he18f;
         4'h2353 	:	val_out <= 4'he18f;
         4'h2358 	:	val_out <= 4'he19f;
         4'h2359 	:	val_out <= 4'he19f;
         4'h235a 	:	val_out <= 4'he19f;
         4'h235b 	:	val_out <= 4'he19f;
         4'h2360 	:	val_out <= 4'he1b0;
         4'h2361 	:	val_out <= 4'he1b0;
         4'h2362 	:	val_out <= 4'he1b0;
         4'h2363 	:	val_out <= 4'he1b0;
         4'h2368 	:	val_out <= 4'he1c0;
         4'h2369 	:	val_out <= 4'he1c0;
         4'h236a 	:	val_out <= 4'he1c0;
         4'h236b 	:	val_out <= 4'he1c0;
         4'h2370 	:	val_out <= 4'he1d0;
         4'h2371 	:	val_out <= 4'he1d0;
         4'h2372 	:	val_out <= 4'he1d0;
         4'h2373 	:	val_out <= 4'he1d0;
         4'h2378 	:	val_out <= 4'he1e0;
         4'h2379 	:	val_out <= 4'he1e0;
         4'h237a 	:	val_out <= 4'he1e0;
         4'h237b 	:	val_out <= 4'he1e0;
         4'h2380 	:	val_out <= 4'he1f1;
         4'h2381 	:	val_out <= 4'he1f1;
         4'h2382 	:	val_out <= 4'he1f1;
         4'h2383 	:	val_out <= 4'he1f1;
         4'h2388 	:	val_out <= 4'he201;
         4'h2389 	:	val_out <= 4'he201;
         4'h238a 	:	val_out <= 4'he201;
         4'h238b 	:	val_out <= 4'he201;
         4'h2390 	:	val_out <= 4'he211;
         4'h2391 	:	val_out <= 4'he211;
         4'h2392 	:	val_out <= 4'he211;
         4'h2393 	:	val_out <= 4'he211;
         4'h2398 	:	val_out <= 4'he221;
         4'h2399 	:	val_out <= 4'he221;
         4'h239a 	:	val_out <= 4'he221;
         4'h239b 	:	val_out <= 4'he221;
         4'h23a0 	:	val_out <= 4'he231;
         4'h23a1 	:	val_out <= 4'he231;
         4'h23a2 	:	val_out <= 4'he231;
         4'h23a3 	:	val_out <= 4'he231;
         4'h23a8 	:	val_out <= 4'he241;
         4'h23a9 	:	val_out <= 4'he241;
         4'h23aa 	:	val_out <= 4'he241;
         4'h23ab 	:	val_out <= 4'he241;
         4'h23b0 	:	val_out <= 4'he251;
         4'h23b1 	:	val_out <= 4'he251;
         4'h23b2 	:	val_out <= 4'he251;
         4'h23b3 	:	val_out <= 4'he251;
         4'h23b8 	:	val_out <= 4'he261;
         4'h23b9 	:	val_out <= 4'he261;
         4'h23ba 	:	val_out <= 4'he261;
         4'h23bb 	:	val_out <= 4'he261;
         4'h23c0 	:	val_out <= 4'he271;
         4'h23c1 	:	val_out <= 4'he271;
         4'h23c2 	:	val_out <= 4'he271;
         4'h23c3 	:	val_out <= 4'he271;
         4'h23c8 	:	val_out <= 4'he282;
         4'h23c9 	:	val_out <= 4'he282;
         4'h23ca 	:	val_out <= 4'he282;
         4'h23cb 	:	val_out <= 4'he282;
         4'h23d0 	:	val_out <= 4'he292;
         4'h23d1 	:	val_out <= 4'he292;
         4'h23d2 	:	val_out <= 4'he292;
         4'h23d3 	:	val_out <= 4'he292;
         4'h23d8 	:	val_out <= 4'he2a2;
         4'h23d9 	:	val_out <= 4'he2a2;
         4'h23da 	:	val_out <= 4'he2a2;
         4'h23db 	:	val_out <= 4'he2a2;
         4'h23e0 	:	val_out <= 4'he2b2;
         4'h23e1 	:	val_out <= 4'he2b2;
         4'h23e2 	:	val_out <= 4'he2b2;
         4'h23e3 	:	val_out <= 4'he2b2;
         4'h23e8 	:	val_out <= 4'he2c2;
         4'h23e9 	:	val_out <= 4'he2c2;
         4'h23ea 	:	val_out <= 4'he2c2;
         4'h23eb 	:	val_out <= 4'he2c2;
         4'h23f0 	:	val_out <= 4'he2d2;
         4'h23f1 	:	val_out <= 4'he2d2;
         4'h23f2 	:	val_out <= 4'he2d2;
         4'h23f3 	:	val_out <= 4'he2d2;
         4'h23f8 	:	val_out <= 4'he2e2;
         4'h23f9 	:	val_out <= 4'he2e2;
         4'h23fa 	:	val_out <= 4'he2e2;
         4'h23fb 	:	val_out <= 4'he2e2;
         4'h2400 	:	val_out <= 4'he2f2;
         4'h2401 	:	val_out <= 4'he2f2;
         4'h2402 	:	val_out <= 4'he2f2;
         4'h2403 	:	val_out <= 4'he2f2;
         4'h2408 	:	val_out <= 4'he301;
         4'h2409 	:	val_out <= 4'he301;
         4'h240a 	:	val_out <= 4'he301;
         4'h240b 	:	val_out <= 4'he301;
         4'h2410 	:	val_out <= 4'he311;
         4'h2411 	:	val_out <= 4'he311;
         4'h2412 	:	val_out <= 4'he311;
         4'h2413 	:	val_out <= 4'he311;
         4'h2418 	:	val_out <= 4'he321;
         4'h2419 	:	val_out <= 4'he321;
         4'h241a 	:	val_out <= 4'he321;
         4'h241b 	:	val_out <= 4'he321;
         4'h2420 	:	val_out <= 4'he331;
         4'h2421 	:	val_out <= 4'he331;
         4'h2422 	:	val_out <= 4'he331;
         4'h2423 	:	val_out <= 4'he331;
         4'h2428 	:	val_out <= 4'he341;
         4'h2429 	:	val_out <= 4'he341;
         4'h242a 	:	val_out <= 4'he341;
         4'h242b 	:	val_out <= 4'he341;
         4'h2430 	:	val_out <= 4'he351;
         4'h2431 	:	val_out <= 4'he351;
         4'h2432 	:	val_out <= 4'he351;
         4'h2433 	:	val_out <= 4'he351;
         4'h2438 	:	val_out <= 4'he361;
         4'h2439 	:	val_out <= 4'he361;
         4'h243a 	:	val_out <= 4'he361;
         4'h243b 	:	val_out <= 4'he361;
         4'h2440 	:	val_out <= 4'he371;
         4'h2441 	:	val_out <= 4'he371;
         4'h2442 	:	val_out <= 4'he371;
         4'h2443 	:	val_out <= 4'he371;
         4'h2448 	:	val_out <= 4'he380;
         4'h2449 	:	val_out <= 4'he380;
         4'h244a 	:	val_out <= 4'he380;
         4'h244b 	:	val_out <= 4'he380;
         4'h2450 	:	val_out <= 4'he390;
         4'h2451 	:	val_out <= 4'he390;
         4'h2452 	:	val_out <= 4'he390;
         4'h2453 	:	val_out <= 4'he390;
         4'h2458 	:	val_out <= 4'he3a0;
         4'h2459 	:	val_out <= 4'he3a0;
         4'h245a 	:	val_out <= 4'he3a0;
         4'h245b 	:	val_out <= 4'he3a0;
         4'h2460 	:	val_out <= 4'he3b0;
         4'h2461 	:	val_out <= 4'he3b0;
         4'h2462 	:	val_out <= 4'he3b0;
         4'h2463 	:	val_out <= 4'he3b0;
         4'h2468 	:	val_out <= 4'he3c0;
         4'h2469 	:	val_out <= 4'he3c0;
         4'h246a 	:	val_out <= 4'he3c0;
         4'h246b 	:	val_out <= 4'he3c0;
         4'h2470 	:	val_out <= 4'he3cf;
         4'h2471 	:	val_out <= 4'he3cf;
         4'h2472 	:	val_out <= 4'he3cf;
         4'h2473 	:	val_out <= 4'he3cf;
         4'h2478 	:	val_out <= 4'he3df;
         4'h2479 	:	val_out <= 4'he3df;
         4'h247a 	:	val_out <= 4'he3df;
         4'h247b 	:	val_out <= 4'he3df;
         4'h2480 	:	val_out <= 4'he3ef;
         4'h2481 	:	val_out <= 4'he3ef;
         4'h2482 	:	val_out <= 4'he3ef;
         4'h2483 	:	val_out <= 4'he3ef;
         4'h2488 	:	val_out <= 4'he3fe;
         4'h2489 	:	val_out <= 4'he3fe;
         4'h248a 	:	val_out <= 4'he3fe;
         4'h248b 	:	val_out <= 4'he3fe;
         4'h2490 	:	val_out <= 4'he40e;
         4'h2491 	:	val_out <= 4'he40e;
         4'h2492 	:	val_out <= 4'he40e;
         4'h2493 	:	val_out <= 4'he40e;
         4'h2498 	:	val_out <= 4'he41e;
         4'h2499 	:	val_out <= 4'he41e;
         4'h249a 	:	val_out <= 4'he41e;
         4'h249b 	:	val_out <= 4'he41e;
         4'h24a0 	:	val_out <= 4'he42d;
         4'h24a1 	:	val_out <= 4'he42d;
         4'h24a2 	:	val_out <= 4'he42d;
         4'h24a3 	:	val_out <= 4'he42d;
         4'h24a8 	:	val_out <= 4'he43d;
         4'h24a9 	:	val_out <= 4'he43d;
         4'h24aa 	:	val_out <= 4'he43d;
         4'h24ab 	:	val_out <= 4'he43d;
         4'h24b0 	:	val_out <= 4'he44d;
         4'h24b1 	:	val_out <= 4'he44d;
         4'h24b2 	:	val_out <= 4'he44d;
         4'h24b3 	:	val_out <= 4'he44d;
         4'h24b8 	:	val_out <= 4'he45c;
         4'h24b9 	:	val_out <= 4'he45c;
         4'h24ba 	:	val_out <= 4'he45c;
         4'h24bb 	:	val_out <= 4'he45c;
         4'h24c0 	:	val_out <= 4'he46c;
         4'h24c1 	:	val_out <= 4'he46c;
         4'h24c2 	:	val_out <= 4'he46c;
         4'h24c3 	:	val_out <= 4'he46c;
         4'h24c8 	:	val_out <= 4'he47b;
         4'h24c9 	:	val_out <= 4'he47b;
         4'h24ca 	:	val_out <= 4'he47b;
         4'h24cb 	:	val_out <= 4'he47b;
         4'h24d0 	:	val_out <= 4'he48b;
         4'h24d1 	:	val_out <= 4'he48b;
         4'h24d2 	:	val_out <= 4'he48b;
         4'h24d3 	:	val_out <= 4'he48b;
         4'h24d8 	:	val_out <= 4'he49b;
         4'h24d9 	:	val_out <= 4'he49b;
         4'h24da 	:	val_out <= 4'he49b;
         4'h24db 	:	val_out <= 4'he49b;
         4'h24e0 	:	val_out <= 4'he4aa;
         4'h24e1 	:	val_out <= 4'he4aa;
         4'h24e2 	:	val_out <= 4'he4aa;
         4'h24e3 	:	val_out <= 4'he4aa;
         4'h24e8 	:	val_out <= 4'he4ba;
         4'h24e9 	:	val_out <= 4'he4ba;
         4'h24ea 	:	val_out <= 4'he4ba;
         4'h24eb 	:	val_out <= 4'he4ba;
         4'h24f0 	:	val_out <= 4'he4c9;
         4'h24f1 	:	val_out <= 4'he4c9;
         4'h24f2 	:	val_out <= 4'he4c9;
         4'h24f3 	:	val_out <= 4'he4c9;
         4'h24f8 	:	val_out <= 4'he4d9;
         4'h24f9 	:	val_out <= 4'he4d9;
         4'h24fa 	:	val_out <= 4'he4d9;
         4'h24fb 	:	val_out <= 4'he4d9;
         4'h2500 	:	val_out <= 4'he4e8;
         4'h2501 	:	val_out <= 4'he4e8;
         4'h2502 	:	val_out <= 4'he4e8;
         4'h2503 	:	val_out <= 4'he4e8;
         4'h2508 	:	val_out <= 4'he4f7;
         4'h2509 	:	val_out <= 4'he4f7;
         4'h250a 	:	val_out <= 4'he4f7;
         4'h250b 	:	val_out <= 4'he4f7;
         4'h2510 	:	val_out <= 4'he507;
         4'h2511 	:	val_out <= 4'he507;
         4'h2512 	:	val_out <= 4'he507;
         4'h2513 	:	val_out <= 4'he507;
         4'h2518 	:	val_out <= 4'he516;
         4'h2519 	:	val_out <= 4'he516;
         4'h251a 	:	val_out <= 4'he516;
         4'h251b 	:	val_out <= 4'he516;
         4'h2520 	:	val_out <= 4'he526;
         4'h2521 	:	val_out <= 4'he526;
         4'h2522 	:	val_out <= 4'he526;
         4'h2523 	:	val_out <= 4'he526;
         4'h2528 	:	val_out <= 4'he535;
         4'h2529 	:	val_out <= 4'he535;
         4'h252a 	:	val_out <= 4'he535;
         4'h252b 	:	val_out <= 4'he535;
         4'h2530 	:	val_out <= 4'he545;
         4'h2531 	:	val_out <= 4'he545;
         4'h2532 	:	val_out <= 4'he545;
         4'h2533 	:	val_out <= 4'he545;
         4'h2538 	:	val_out <= 4'he554;
         4'h2539 	:	val_out <= 4'he554;
         4'h253a 	:	val_out <= 4'he554;
         4'h253b 	:	val_out <= 4'he554;
         4'h2540 	:	val_out <= 4'he563;
         4'h2541 	:	val_out <= 4'he563;
         4'h2542 	:	val_out <= 4'he563;
         4'h2543 	:	val_out <= 4'he563;
         4'h2548 	:	val_out <= 4'he573;
         4'h2549 	:	val_out <= 4'he573;
         4'h254a 	:	val_out <= 4'he573;
         4'h254b 	:	val_out <= 4'he573;
         4'h2550 	:	val_out <= 4'he582;
         4'h2551 	:	val_out <= 4'he582;
         4'h2552 	:	val_out <= 4'he582;
         4'h2553 	:	val_out <= 4'he582;
         4'h2558 	:	val_out <= 4'he591;
         4'h2559 	:	val_out <= 4'he591;
         4'h255a 	:	val_out <= 4'he591;
         4'h255b 	:	val_out <= 4'he591;
         4'h2560 	:	val_out <= 4'he5a0;
         4'h2561 	:	val_out <= 4'he5a0;
         4'h2562 	:	val_out <= 4'he5a0;
         4'h2563 	:	val_out <= 4'he5a0;
         4'h2568 	:	val_out <= 4'he5b0;
         4'h2569 	:	val_out <= 4'he5b0;
         4'h256a 	:	val_out <= 4'he5b0;
         4'h256b 	:	val_out <= 4'he5b0;
         4'h2570 	:	val_out <= 4'he5bf;
         4'h2571 	:	val_out <= 4'he5bf;
         4'h2572 	:	val_out <= 4'he5bf;
         4'h2573 	:	val_out <= 4'he5bf;
         4'h2578 	:	val_out <= 4'he5ce;
         4'h2579 	:	val_out <= 4'he5ce;
         4'h257a 	:	val_out <= 4'he5ce;
         4'h257b 	:	val_out <= 4'he5ce;
         4'h2580 	:	val_out <= 4'he5dd;
         4'h2581 	:	val_out <= 4'he5dd;
         4'h2582 	:	val_out <= 4'he5dd;
         4'h2583 	:	val_out <= 4'he5dd;
         4'h2588 	:	val_out <= 4'he5ed;
         4'h2589 	:	val_out <= 4'he5ed;
         4'h258a 	:	val_out <= 4'he5ed;
         4'h258b 	:	val_out <= 4'he5ed;
         4'h2590 	:	val_out <= 4'he5fc;
         4'h2591 	:	val_out <= 4'he5fc;
         4'h2592 	:	val_out <= 4'he5fc;
         4'h2593 	:	val_out <= 4'he5fc;
         4'h2598 	:	val_out <= 4'he60b;
         4'h2599 	:	val_out <= 4'he60b;
         4'h259a 	:	val_out <= 4'he60b;
         4'h259b 	:	val_out <= 4'he60b;
         4'h25a0 	:	val_out <= 4'he61a;
         4'h25a1 	:	val_out <= 4'he61a;
         4'h25a2 	:	val_out <= 4'he61a;
         4'h25a3 	:	val_out <= 4'he61a;
         4'h25a8 	:	val_out <= 4'he629;
         4'h25a9 	:	val_out <= 4'he629;
         4'h25aa 	:	val_out <= 4'he629;
         4'h25ab 	:	val_out <= 4'he629;
         4'h25b0 	:	val_out <= 4'he639;
         4'h25b1 	:	val_out <= 4'he639;
         4'h25b2 	:	val_out <= 4'he639;
         4'h25b3 	:	val_out <= 4'he639;
         4'h25b8 	:	val_out <= 4'he648;
         4'h25b9 	:	val_out <= 4'he648;
         4'h25ba 	:	val_out <= 4'he648;
         4'h25bb 	:	val_out <= 4'he648;
         4'h25c0 	:	val_out <= 4'he657;
         4'h25c1 	:	val_out <= 4'he657;
         4'h25c2 	:	val_out <= 4'he657;
         4'h25c3 	:	val_out <= 4'he657;
         4'h25c8 	:	val_out <= 4'he666;
         4'h25c9 	:	val_out <= 4'he666;
         4'h25ca 	:	val_out <= 4'he666;
         4'h25cb 	:	val_out <= 4'he666;
         4'h25d0 	:	val_out <= 4'he675;
         4'h25d1 	:	val_out <= 4'he675;
         4'h25d2 	:	val_out <= 4'he675;
         4'h25d3 	:	val_out <= 4'he675;
         4'h25d8 	:	val_out <= 4'he684;
         4'h25d9 	:	val_out <= 4'he684;
         4'h25da 	:	val_out <= 4'he684;
         4'h25db 	:	val_out <= 4'he684;
         4'h25e0 	:	val_out <= 4'he693;
         4'h25e1 	:	val_out <= 4'he693;
         4'h25e2 	:	val_out <= 4'he693;
         4'h25e3 	:	val_out <= 4'he693;
         4'h25e8 	:	val_out <= 4'he6a2;
         4'h25e9 	:	val_out <= 4'he6a2;
         4'h25ea 	:	val_out <= 4'he6a2;
         4'h25eb 	:	val_out <= 4'he6a2;
         4'h25f0 	:	val_out <= 4'he6b1;
         4'h25f1 	:	val_out <= 4'he6b1;
         4'h25f2 	:	val_out <= 4'he6b1;
         4'h25f3 	:	val_out <= 4'he6b1;
         4'h25f8 	:	val_out <= 4'he6c0;
         4'h25f9 	:	val_out <= 4'he6c0;
         4'h25fa 	:	val_out <= 4'he6c0;
         4'h25fb 	:	val_out <= 4'he6c0;
         4'h2600 	:	val_out <= 4'he6cf;
         4'h2601 	:	val_out <= 4'he6cf;
         4'h2602 	:	val_out <= 4'he6cf;
         4'h2603 	:	val_out <= 4'he6cf;
         4'h2608 	:	val_out <= 4'he6de;
         4'h2609 	:	val_out <= 4'he6de;
         4'h260a 	:	val_out <= 4'he6de;
         4'h260b 	:	val_out <= 4'he6de;
         4'h2610 	:	val_out <= 4'he6ed;
         4'h2611 	:	val_out <= 4'he6ed;
         4'h2612 	:	val_out <= 4'he6ed;
         4'h2613 	:	val_out <= 4'he6ed;
         4'h2618 	:	val_out <= 4'he6fc;
         4'h2619 	:	val_out <= 4'he6fc;
         4'h261a 	:	val_out <= 4'he6fc;
         4'h261b 	:	val_out <= 4'he6fc;
         4'h2620 	:	val_out <= 4'he70b;
         4'h2621 	:	val_out <= 4'he70b;
         4'h2622 	:	val_out <= 4'he70b;
         4'h2623 	:	val_out <= 4'he70b;
         4'h2628 	:	val_out <= 4'he71a;
         4'h2629 	:	val_out <= 4'he71a;
         4'h262a 	:	val_out <= 4'he71a;
         4'h262b 	:	val_out <= 4'he71a;
         4'h2630 	:	val_out <= 4'he729;
         4'h2631 	:	val_out <= 4'he729;
         4'h2632 	:	val_out <= 4'he729;
         4'h2633 	:	val_out <= 4'he729;
         4'h2638 	:	val_out <= 4'he737;
         4'h2639 	:	val_out <= 4'he737;
         4'h263a 	:	val_out <= 4'he737;
         4'h263b 	:	val_out <= 4'he737;
         4'h2640 	:	val_out <= 4'he746;
         4'h2641 	:	val_out <= 4'he746;
         4'h2642 	:	val_out <= 4'he746;
         4'h2643 	:	val_out <= 4'he746;
         4'h2648 	:	val_out <= 4'he755;
         4'h2649 	:	val_out <= 4'he755;
         4'h264a 	:	val_out <= 4'he755;
         4'h264b 	:	val_out <= 4'he755;
         4'h2650 	:	val_out <= 4'he764;
         4'h2651 	:	val_out <= 4'he764;
         4'h2652 	:	val_out <= 4'he764;
         4'h2653 	:	val_out <= 4'he764;
         4'h2658 	:	val_out <= 4'he773;
         4'h2659 	:	val_out <= 4'he773;
         4'h265a 	:	val_out <= 4'he773;
         4'h265b 	:	val_out <= 4'he773;
         4'h2660 	:	val_out <= 4'he782;
         4'h2661 	:	val_out <= 4'he782;
         4'h2662 	:	val_out <= 4'he782;
         4'h2663 	:	val_out <= 4'he782;
         4'h2668 	:	val_out <= 4'he790;
         4'h2669 	:	val_out <= 4'he790;
         4'h266a 	:	val_out <= 4'he790;
         4'h266b 	:	val_out <= 4'he790;
         4'h2670 	:	val_out <= 4'he79f;
         4'h2671 	:	val_out <= 4'he79f;
         4'h2672 	:	val_out <= 4'he79f;
         4'h2673 	:	val_out <= 4'he79f;
         4'h2678 	:	val_out <= 4'he7ae;
         4'h2679 	:	val_out <= 4'he7ae;
         4'h267a 	:	val_out <= 4'he7ae;
         4'h267b 	:	val_out <= 4'he7ae;
         4'h2680 	:	val_out <= 4'he7bd;
         4'h2681 	:	val_out <= 4'he7bd;
         4'h2682 	:	val_out <= 4'he7bd;
         4'h2683 	:	val_out <= 4'he7bd;
         4'h2688 	:	val_out <= 4'he7cb;
         4'h2689 	:	val_out <= 4'he7cb;
         4'h268a 	:	val_out <= 4'he7cb;
         4'h268b 	:	val_out <= 4'he7cb;
         4'h2690 	:	val_out <= 4'he7da;
         4'h2691 	:	val_out <= 4'he7da;
         4'h2692 	:	val_out <= 4'he7da;
         4'h2693 	:	val_out <= 4'he7da;
         4'h2698 	:	val_out <= 4'he7e9;
         4'h2699 	:	val_out <= 4'he7e9;
         4'h269a 	:	val_out <= 4'he7e9;
         4'h269b 	:	val_out <= 4'he7e9;
         4'h26a0 	:	val_out <= 4'he7f7;
         4'h26a1 	:	val_out <= 4'he7f7;
         4'h26a2 	:	val_out <= 4'he7f7;
         4'h26a3 	:	val_out <= 4'he7f7;
         4'h26a8 	:	val_out <= 4'he806;
         4'h26a9 	:	val_out <= 4'he806;
         4'h26aa 	:	val_out <= 4'he806;
         4'h26ab 	:	val_out <= 4'he806;
         4'h26b0 	:	val_out <= 4'he815;
         4'h26b1 	:	val_out <= 4'he815;
         4'h26b2 	:	val_out <= 4'he815;
         4'h26b3 	:	val_out <= 4'he815;
         4'h26b8 	:	val_out <= 4'he823;
         4'h26b9 	:	val_out <= 4'he823;
         4'h26ba 	:	val_out <= 4'he823;
         4'h26bb 	:	val_out <= 4'he823;
         4'h26c0 	:	val_out <= 4'he832;
         4'h26c1 	:	val_out <= 4'he832;
         4'h26c2 	:	val_out <= 4'he832;
         4'h26c3 	:	val_out <= 4'he832;
         4'h26c8 	:	val_out <= 4'he840;
         4'h26c9 	:	val_out <= 4'he840;
         4'h26ca 	:	val_out <= 4'he840;
         4'h26cb 	:	val_out <= 4'he840;
         4'h26d0 	:	val_out <= 4'he84f;
         4'h26d1 	:	val_out <= 4'he84f;
         4'h26d2 	:	val_out <= 4'he84f;
         4'h26d3 	:	val_out <= 4'he84f;
         4'h26d8 	:	val_out <= 4'he85e;
         4'h26d9 	:	val_out <= 4'he85e;
         4'h26da 	:	val_out <= 4'he85e;
         4'h26db 	:	val_out <= 4'he85e;
         4'h26e0 	:	val_out <= 4'he86c;
         4'h26e1 	:	val_out <= 4'he86c;
         4'h26e2 	:	val_out <= 4'he86c;
         4'h26e3 	:	val_out <= 4'he86c;
         4'h26e8 	:	val_out <= 4'he87b;
         4'h26e9 	:	val_out <= 4'he87b;
         4'h26ea 	:	val_out <= 4'he87b;
         4'h26eb 	:	val_out <= 4'he87b;
         4'h26f0 	:	val_out <= 4'he889;
         4'h26f1 	:	val_out <= 4'he889;
         4'h26f2 	:	val_out <= 4'he889;
         4'h26f3 	:	val_out <= 4'he889;
         4'h26f8 	:	val_out <= 4'he898;
         4'h26f9 	:	val_out <= 4'he898;
         4'h26fa 	:	val_out <= 4'he898;
         4'h26fb 	:	val_out <= 4'he898;
         4'h2700 	:	val_out <= 4'he8a6;
         4'h2701 	:	val_out <= 4'he8a6;
         4'h2702 	:	val_out <= 4'he8a6;
         4'h2703 	:	val_out <= 4'he8a6;
         4'h2708 	:	val_out <= 4'he8b5;
         4'h2709 	:	val_out <= 4'he8b5;
         4'h270a 	:	val_out <= 4'he8b5;
         4'h270b 	:	val_out <= 4'he8b5;
         4'h2710 	:	val_out <= 4'he8c3;
         4'h2711 	:	val_out <= 4'he8c3;
         4'h2712 	:	val_out <= 4'he8c3;
         4'h2713 	:	val_out <= 4'he8c3;
         4'h2718 	:	val_out <= 4'he8d1;
         4'h2719 	:	val_out <= 4'he8d1;
         4'h271a 	:	val_out <= 4'he8d1;
         4'h271b 	:	val_out <= 4'he8d1;
         4'h2720 	:	val_out <= 4'he8e0;
         4'h2721 	:	val_out <= 4'he8e0;
         4'h2722 	:	val_out <= 4'he8e0;
         4'h2723 	:	val_out <= 4'he8e0;
         4'h2728 	:	val_out <= 4'he8ee;
         4'h2729 	:	val_out <= 4'he8ee;
         4'h272a 	:	val_out <= 4'he8ee;
         4'h272b 	:	val_out <= 4'he8ee;
         4'h2730 	:	val_out <= 4'he8fd;
         4'h2731 	:	val_out <= 4'he8fd;
         4'h2732 	:	val_out <= 4'he8fd;
         4'h2733 	:	val_out <= 4'he8fd;
         4'h2738 	:	val_out <= 4'he90b;
         4'h2739 	:	val_out <= 4'he90b;
         4'h273a 	:	val_out <= 4'he90b;
         4'h273b 	:	val_out <= 4'he90b;
         4'h2740 	:	val_out <= 4'he919;
         4'h2741 	:	val_out <= 4'he919;
         4'h2742 	:	val_out <= 4'he919;
         4'h2743 	:	val_out <= 4'he919;
         4'h2748 	:	val_out <= 4'he928;
         4'h2749 	:	val_out <= 4'he928;
         4'h274a 	:	val_out <= 4'he928;
         4'h274b 	:	val_out <= 4'he928;
         4'h2750 	:	val_out <= 4'he936;
         4'h2751 	:	val_out <= 4'he936;
         4'h2752 	:	val_out <= 4'he936;
         4'h2753 	:	val_out <= 4'he936;
         4'h2758 	:	val_out <= 4'he944;
         4'h2759 	:	val_out <= 4'he944;
         4'h275a 	:	val_out <= 4'he944;
         4'h275b 	:	val_out <= 4'he944;
         4'h2760 	:	val_out <= 4'he953;
         4'h2761 	:	val_out <= 4'he953;
         4'h2762 	:	val_out <= 4'he953;
         4'h2763 	:	val_out <= 4'he953;
         4'h2768 	:	val_out <= 4'he961;
         4'h2769 	:	val_out <= 4'he961;
         4'h276a 	:	val_out <= 4'he961;
         4'h276b 	:	val_out <= 4'he961;
         4'h2770 	:	val_out <= 4'he96f;
         4'h2771 	:	val_out <= 4'he96f;
         4'h2772 	:	val_out <= 4'he96f;
         4'h2773 	:	val_out <= 4'he96f;
         4'h2778 	:	val_out <= 4'he97d;
         4'h2779 	:	val_out <= 4'he97d;
         4'h277a 	:	val_out <= 4'he97d;
         4'h277b 	:	val_out <= 4'he97d;
         4'h2780 	:	val_out <= 4'he98c;
         4'h2781 	:	val_out <= 4'he98c;
         4'h2782 	:	val_out <= 4'he98c;
         4'h2783 	:	val_out <= 4'he98c;
         4'h2788 	:	val_out <= 4'he99a;
         4'h2789 	:	val_out <= 4'he99a;
         4'h278a 	:	val_out <= 4'he99a;
         4'h278b 	:	val_out <= 4'he99a;
         4'h2790 	:	val_out <= 4'he9a8;
         4'h2791 	:	val_out <= 4'he9a8;
         4'h2792 	:	val_out <= 4'he9a8;
         4'h2793 	:	val_out <= 4'he9a8;
         4'h2798 	:	val_out <= 4'he9b6;
         4'h2799 	:	val_out <= 4'he9b6;
         4'h279a 	:	val_out <= 4'he9b6;
         4'h279b 	:	val_out <= 4'he9b6;
         4'h27a0 	:	val_out <= 4'he9c4;
         4'h27a1 	:	val_out <= 4'he9c4;
         4'h27a2 	:	val_out <= 4'he9c4;
         4'h27a3 	:	val_out <= 4'he9c4;
         4'h27a8 	:	val_out <= 4'he9d3;
         4'h27a9 	:	val_out <= 4'he9d3;
         4'h27aa 	:	val_out <= 4'he9d3;
         4'h27ab 	:	val_out <= 4'he9d3;
         4'h27b0 	:	val_out <= 4'he9e1;
         4'h27b1 	:	val_out <= 4'he9e1;
         4'h27b2 	:	val_out <= 4'he9e1;
         4'h27b3 	:	val_out <= 4'he9e1;
         4'h27b8 	:	val_out <= 4'he9ef;
         4'h27b9 	:	val_out <= 4'he9ef;
         4'h27ba 	:	val_out <= 4'he9ef;
         4'h27bb 	:	val_out <= 4'he9ef;
         4'h27c0 	:	val_out <= 4'he9fd;
         4'h27c1 	:	val_out <= 4'he9fd;
         4'h27c2 	:	val_out <= 4'he9fd;
         4'h27c3 	:	val_out <= 4'he9fd;
         4'h27c8 	:	val_out <= 4'hea0b;
         4'h27c9 	:	val_out <= 4'hea0b;
         4'h27ca 	:	val_out <= 4'hea0b;
         4'h27cb 	:	val_out <= 4'hea0b;
         4'h27d0 	:	val_out <= 4'hea19;
         4'h27d1 	:	val_out <= 4'hea19;
         4'h27d2 	:	val_out <= 4'hea19;
         4'h27d3 	:	val_out <= 4'hea19;
         4'h27d8 	:	val_out <= 4'hea27;
         4'h27d9 	:	val_out <= 4'hea27;
         4'h27da 	:	val_out <= 4'hea27;
         4'h27db 	:	val_out <= 4'hea27;
         4'h27e0 	:	val_out <= 4'hea35;
         4'h27e1 	:	val_out <= 4'hea35;
         4'h27e2 	:	val_out <= 4'hea35;
         4'h27e3 	:	val_out <= 4'hea35;
         4'h27e8 	:	val_out <= 4'hea43;
         4'h27e9 	:	val_out <= 4'hea43;
         4'h27ea 	:	val_out <= 4'hea43;
         4'h27eb 	:	val_out <= 4'hea43;
         4'h27f0 	:	val_out <= 4'hea51;
         4'h27f1 	:	val_out <= 4'hea51;
         4'h27f2 	:	val_out <= 4'hea51;
         4'h27f3 	:	val_out <= 4'hea51;
         4'h27f8 	:	val_out <= 4'hea5f;
         4'h27f9 	:	val_out <= 4'hea5f;
         4'h27fa 	:	val_out <= 4'hea5f;
         4'h27fb 	:	val_out <= 4'hea5f;
         4'h2800 	:	val_out <= 4'hea6d;
         4'h2801 	:	val_out <= 4'hea6d;
         4'h2802 	:	val_out <= 4'hea6d;
         4'h2803 	:	val_out <= 4'hea6d;
         4'h2808 	:	val_out <= 4'hea7b;
         4'h2809 	:	val_out <= 4'hea7b;
         4'h280a 	:	val_out <= 4'hea7b;
         4'h280b 	:	val_out <= 4'hea7b;
         4'h2810 	:	val_out <= 4'hea89;
         4'h2811 	:	val_out <= 4'hea89;
         4'h2812 	:	val_out <= 4'hea89;
         4'h2813 	:	val_out <= 4'hea89;
         4'h2818 	:	val_out <= 4'hea97;
         4'h2819 	:	val_out <= 4'hea97;
         4'h281a 	:	val_out <= 4'hea97;
         4'h281b 	:	val_out <= 4'hea97;
         4'h2820 	:	val_out <= 4'heaa5;
         4'h2821 	:	val_out <= 4'heaa5;
         4'h2822 	:	val_out <= 4'heaa5;
         4'h2823 	:	val_out <= 4'heaa5;
         4'h2828 	:	val_out <= 4'heab3;
         4'h2829 	:	val_out <= 4'heab3;
         4'h282a 	:	val_out <= 4'heab3;
         4'h282b 	:	val_out <= 4'heab3;
         4'h2830 	:	val_out <= 4'heac1;
         4'h2831 	:	val_out <= 4'heac1;
         4'h2832 	:	val_out <= 4'heac1;
         4'h2833 	:	val_out <= 4'heac1;
         4'h2838 	:	val_out <= 4'heace;
         4'h2839 	:	val_out <= 4'heace;
         4'h283a 	:	val_out <= 4'heace;
         4'h283b 	:	val_out <= 4'heace;
         4'h2840 	:	val_out <= 4'headc;
         4'h2841 	:	val_out <= 4'headc;
         4'h2842 	:	val_out <= 4'headc;
         4'h2843 	:	val_out <= 4'headc;
         4'h2848 	:	val_out <= 4'heaea;
         4'h2849 	:	val_out <= 4'heaea;
         4'h284a 	:	val_out <= 4'heaea;
         4'h284b 	:	val_out <= 4'heaea;
         4'h2850 	:	val_out <= 4'heaf8;
         4'h2851 	:	val_out <= 4'heaf8;
         4'h2852 	:	val_out <= 4'heaf8;
         4'h2853 	:	val_out <= 4'heaf8;
         4'h2858 	:	val_out <= 4'heb06;
         4'h2859 	:	val_out <= 4'heb06;
         4'h285a 	:	val_out <= 4'heb06;
         4'h285b 	:	val_out <= 4'heb06;
         4'h2860 	:	val_out <= 4'heb13;
         4'h2861 	:	val_out <= 4'heb13;
         4'h2862 	:	val_out <= 4'heb13;
         4'h2863 	:	val_out <= 4'heb13;
         4'h2868 	:	val_out <= 4'heb21;
         4'h2869 	:	val_out <= 4'heb21;
         4'h286a 	:	val_out <= 4'heb21;
         4'h286b 	:	val_out <= 4'heb21;
         4'h2870 	:	val_out <= 4'heb2f;
         4'h2871 	:	val_out <= 4'heb2f;
         4'h2872 	:	val_out <= 4'heb2f;
         4'h2873 	:	val_out <= 4'heb2f;
         4'h2878 	:	val_out <= 4'heb3d;
         4'h2879 	:	val_out <= 4'heb3d;
         4'h287a 	:	val_out <= 4'heb3d;
         4'h287b 	:	val_out <= 4'heb3d;
         4'h2880 	:	val_out <= 4'heb4a;
         4'h2881 	:	val_out <= 4'heb4a;
         4'h2882 	:	val_out <= 4'heb4a;
         4'h2883 	:	val_out <= 4'heb4a;
         4'h2888 	:	val_out <= 4'heb58;
         4'h2889 	:	val_out <= 4'heb58;
         4'h288a 	:	val_out <= 4'heb58;
         4'h288b 	:	val_out <= 4'heb58;
         4'h2890 	:	val_out <= 4'heb66;
         4'h2891 	:	val_out <= 4'heb66;
         4'h2892 	:	val_out <= 4'heb66;
         4'h2893 	:	val_out <= 4'heb66;
         4'h2898 	:	val_out <= 4'heb73;
         4'h2899 	:	val_out <= 4'heb73;
         4'h289a 	:	val_out <= 4'heb73;
         4'h289b 	:	val_out <= 4'heb73;
         4'h28a0 	:	val_out <= 4'heb81;
         4'h28a1 	:	val_out <= 4'heb81;
         4'h28a2 	:	val_out <= 4'heb81;
         4'h28a3 	:	val_out <= 4'heb81;
         4'h28a8 	:	val_out <= 4'heb8f;
         4'h28a9 	:	val_out <= 4'heb8f;
         4'h28aa 	:	val_out <= 4'heb8f;
         4'h28ab 	:	val_out <= 4'heb8f;
         4'h28b0 	:	val_out <= 4'heb9c;
         4'h28b1 	:	val_out <= 4'heb9c;
         4'h28b2 	:	val_out <= 4'heb9c;
         4'h28b3 	:	val_out <= 4'heb9c;
         4'h28b8 	:	val_out <= 4'hebaa;
         4'h28b9 	:	val_out <= 4'hebaa;
         4'h28ba 	:	val_out <= 4'hebaa;
         4'h28bb 	:	val_out <= 4'hebaa;
         4'h28c0 	:	val_out <= 4'hebb8;
         4'h28c1 	:	val_out <= 4'hebb8;
         4'h28c2 	:	val_out <= 4'hebb8;
         4'h28c3 	:	val_out <= 4'hebb8;
         4'h28c8 	:	val_out <= 4'hebc5;
         4'h28c9 	:	val_out <= 4'hebc5;
         4'h28ca 	:	val_out <= 4'hebc5;
         4'h28cb 	:	val_out <= 4'hebc5;
         4'h28d0 	:	val_out <= 4'hebd3;
         4'h28d1 	:	val_out <= 4'hebd3;
         4'h28d2 	:	val_out <= 4'hebd3;
         4'h28d3 	:	val_out <= 4'hebd3;
         4'h28d8 	:	val_out <= 4'hebe0;
         4'h28d9 	:	val_out <= 4'hebe0;
         4'h28da 	:	val_out <= 4'hebe0;
         4'h28db 	:	val_out <= 4'hebe0;
         4'h28e0 	:	val_out <= 4'hebee;
         4'h28e1 	:	val_out <= 4'hebee;
         4'h28e2 	:	val_out <= 4'hebee;
         4'h28e3 	:	val_out <= 4'hebee;
         4'h28e8 	:	val_out <= 4'hebfb;
         4'h28e9 	:	val_out <= 4'hebfb;
         4'h28ea 	:	val_out <= 4'hebfb;
         4'h28eb 	:	val_out <= 4'hebfb;
         4'h28f0 	:	val_out <= 4'hec09;
         4'h28f1 	:	val_out <= 4'hec09;
         4'h28f2 	:	val_out <= 4'hec09;
         4'h28f3 	:	val_out <= 4'hec09;
         4'h28f8 	:	val_out <= 4'hec16;
         4'h28f9 	:	val_out <= 4'hec16;
         4'h28fa 	:	val_out <= 4'hec16;
         4'h28fb 	:	val_out <= 4'hec16;
         4'h2900 	:	val_out <= 4'hec24;
         4'h2901 	:	val_out <= 4'hec24;
         4'h2902 	:	val_out <= 4'hec24;
         4'h2903 	:	val_out <= 4'hec24;
         4'h2908 	:	val_out <= 4'hec31;
         4'h2909 	:	val_out <= 4'hec31;
         4'h290a 	:	val_out <= 4'hec31;
         4'h290b 	:	val_out <= 4'hec31;
         4'h2910 	:	val_out <= 4'hec3f;
         4'h2911 	:	val_out <= 4'hec3f;
         4'h2912 	:	val_out <= 4'hec3f;
         4'h2913 	:	val_out <= 4'hec3f;
         4'h2918 	:	val_out <= 4'hec4c;
         4'h2919 	:	val_out <= 4'hec4c;
         4'h291a 	:	val_out <= 4'hec4c;
         4'h291b 	:	val_out <= 4'hec4c;
         4'h2920 	:	val_out <= 4'hec59;
         4'h2921 	:	val_out <= 4'hec59;
         4'h2922 	:	val_out <= 4'hec59;
         4'h2923 	:	val_out <= 4'hec59;
         4'h2928 	:	val_out <= 4'hec67;
         4'h2929 	:	val_out <= 4'hec67;
         4'h292a 	:	val_out <= 4'hec67;
         4'h292b 	:	val_out <= 4'hec67;
         4'h2930 	:	val_out <= 4'hec74;
         4'h2931 	:	val_out <= 4'hec74;
         4'h2932 	:	val_out <= 4'hec74;
         4'h2933 	:	val_out <= 4'hec74;
         4'h2938 	:	val_out <= 4'hec81;
         4'h2939 	:	val_out <= 4'hec81;
         4'h293a 	:	val_out <= 4'hec81;
         4'h293b 	:	val_out <= 4'hec81;
         4'h2940 	:	val_out <= 4'hec8f;
         4'h2941 	:	val_out <= 4'hec8f;
         4'h2942 	:	val_out <= 4'hec8f;
         4'h2943 	:	val_out <= 4'hec8f;
         4'h2948 	:	val_out <= 4'hec9c;
         4'h2949 	:	val_out <= 4'hec9c;
         4'h294a 	:	val_out <= 4'hec9c;
         4'h294b 	:	val_out <= 4'hec9c;
         4'h2950 	:	val_out <= 4'heca9;
         4'h2951 	:	val_out <= 4'heca9;
         4'h2952 	:	val_out <= 4'heca9;
         4'h2953 	:	val_out <= 4'heca9;
         4'h2958 	:	val_out <= 4'hecb7;
         4'h2959 	:	val_out <= 4'hecb7;
         4'h295a 	:	val_out <= 4'hecb7;
         4'h295b 	:	val_out <= 4'hecb7;
         4'h2960 	:	val_out <= 4'hecc4;
         4'h2961 	:	val_out <= 4'hecc4;
         4'h2962 	:	val_out <= 4'hecc4;
         4'h2963 	:	val_out <= 4'hecc4;
         4'h2968 	:	val_out <= 4'hecd1;
         4'h2969 	:	val_out <= 4'hecd1;
         4'h296a 	:	val_out <= 4'hecd1;
         4'h296b 	:	val_out <= 4'hecd1;
         4'h2970 	:	val_out <= 4'hecde;
         4'h2971 	:	val_out <= 4'hecde;
         4'h2972 	:	val_out <= 4'hecde;
         4'h2973 	:	val_out <= 4'hecde;
         4'h2978 	:	val_out <= 4'hecec;
         4'h2979 	:	val_out <= 4'hecec;
         4'h297a 	:	val_out <= 4'hecec;
         4'h297b 	:	val_out <= 4'hecec;
         4'h2980 	:	val_out <= 4'hecf9;
         4'h2981 	:	val_out <= 4'hecf9;
         4'h2982 	:	val_out <= 4'hecf9;
         4'h2983 	:	val_out <= 4'hecf9;
         4'h2988 	:	val_out <= 4'hed06;
         4'h2989 	:	val_out <= 4'hed06;
         4'h298a 	:	val_out <= 4'hed06;
         4'h298b 	:	val_out <= 4'hed06;
         4'h2990 	:	val_out <= 4'hed13;
         4'h2991 	:	val_out <= 4'hed13;
         4'h2992 	:	val_out <= 4'hed13;
         4'h2993 	:	val_out <= 4'hed13;
         4'h2998 	:	val_out <= 4'hed20;
         4'h2999 	:	val_out <= 4'hed20;
         4'h299a 	:	val_out <= 4'hed20;
         4'h299b 	:	val_out <= 4'hed20;
         4'h29a0 	:	val_out <= 4'hed2d;
         4'h29a1 	:	val_out <= 4'hed2d;
         4'h29a2 	:	val_out <= 4'hed2d;
         4'h29a3 	:	val_out <= 4'hed2d;
         4'h29a8 	:	val_out <= 4'hed3a;
         4'h29a9 	:	val_out <= 4'hed3a;
         4'h29aa 	:	val_out <= 4'hed3a;
         4'h29ab 	:	val_out <= 4'hed3a;
         4'h29b0 	:	val_out <= 4'hed48;
         4'h29b1 	:	val_out <= 4'hed48;
         4'h29b2 	:	val_out <= 4'hed48;
         4'h29b3 	:	val_out <= 4'hed48;
         4'h29b8 	:	val_out <= 4'hed55;
         4'h29b9 	:	val_out <= 4'hed55;
         4'h29ba 	:	val_out <= 4'hed55;
         4'h29bb 	:	val_out <= 4'hed55;
         4'h29c0 	:	val_out <= 4'hed62;
         4'h29c1 	:	val_out <= 4'hed62;
         4'h29c2 	:	val_out <= 4'hed62;
         4'h29c3 	:	val_out <= 4'hed62;
         4'h29c8 	:	val_out <= 4'hed6f;
         4'h29c9 	:	val_out <= 4'hed6f;
         4'h29ca 	:	val_out <= 4'hed6f;
         4'h29cb 	:	val_out <= 4'hed6f;
         4'h29d0 	:	val_out <= 4'hed7c;
         4'h29d1 	:	val_out <= 4'hed7c;
         4'h29d2 	:	val_out <= 4'hed7c;
         4'h29d3 	:	val_out <= 4'hed7c;
         4'h29d8 	:	val_out <= 4'hed89;
         4'h29d9 	:	val_out <= 4'hed89;
         4'h29da 	:	val_out <= 4'hed89;
         4'h29db 	:	val_out <= 4'hed89;
         4'h29e0 	:	val_out <= 4'hed96;
         4'h29e1 	:	val_out <= 4'hed96;
         4'h29e2 	:	val_out <= 4'hed96;
         4'h29e3 	:	val_out <= 4'hed96;
         4'h29e8 	:	val_out <= 4'heda3;
         4'h29e9 	:	val_out <= 4'heda3;
         4'h29ea 	:	val_out <= 4'heda3;
         4'h29eb 	:	val_out <= 4'heda3;
         4'h29f0 	:	val_out <= 4'hedb0;
         4'h29f1 	:	val_out <= 4'hedb0;
         4'h29f2 	:	val_out <= 4'hedb0;
         4'h29f3 	:	val_out <= 4'hedb0;
         4'h29f8 	:	val_out <= 4'hedbd;
         4'h29f9 	:	val_out <= 4'hedbd;
         4'h29fa 	:	val_out <= 4'hedbd;
         4'h29fb 	:	val_out <= 4'hedbd;
         4'h2a00 	:	val_out <= 4'hedca;
         4'h2a01 	:	val_out <= 4'hedca;
         4'h2a02 	:	val_out <= 4'hedca;
         4'h2a03 	:	val_out <= 4'hedca;
         4'h2a08 	:	val_out <= 4'hedd6;
         4'h2a09 	:	val_out <= 4'hedd6;
         4'h2a0a 	:	val_out <= 4'hedd6;
         4'h2a0b 	:	val_out <= 4'hedd6;
         4'h2a10 	:	val_out <= 4'hede3;
         4'h2a11 	:	val_out <= 4'hede3;
         4'h2a12 	:	val_out <= 4'hede3;
         4'h2a13 	:	val_out <= 4'hede3;
         4'h2a18 	:	val_out <= 4'hedf0;
         4'h2a19 	:	val_out <= 4'hedf0;
         4'h2a1a 	:	val_out <= 4'hedf0;
         4'h2a1b 	:	val_out <= 4'hedf0;
         4'h2a20 	:	val_out <= 4'hedfd;
         4'h2a21 	:	val_out <= 4'hedfd;
         4'h2a22 	:	val_out <= 4'hedfd;
         4'h2a23 	:	val_out <= 4'hedfd;
         4'h2a28 	:	val_out <= 4'hee0a;
         4'h2a29 	:	val_out <= 4'hee0a;
         4'h2a2a 	:	val_out <= 4'hee0a;
         4'h2a2b 	:	val_out <= 4'hee0a;
         4'h2a30 	:	val_out <= 4'hee17;
         4'h2a31 	:	val_out <= 4'hee17;
         4'h2a32 	:	val_out <= 4'hee17;
         4'h2a33 	:	val_out <= 4'hee17;
         4'h2a38 	:	val_out <= 4'hee24;
         4'h2a39 	:	val_out <= 4'hee24;
         4'h2a3a 	:	val_out <= 4'hee24;
         4'h2a3b 	:	val_out <= 4'hee24;
         4'h2a40 	:	val_out <= 4'hee30;
         4'h2a41 	:	val_out <= 4'hee30;
         4'h2a42 	:	val_out <= 4'hee30;
         4'h2a43 	:	val_out <= 4'hee30;
         4'h2a48 	:	val_out <= 4'hee3d;
         4'h2a49 	:	val_out <= 4'hee3d;
         4'h2a4a 	:	val_out <= 4'hee3d;
         4'h2a4b 	:	val_out <= 4'hee3d;
         4'h2a50 	:	val_out <= 4'hee4a;
         4'h2a51 	:	val_out <= 4'hee4a;
         4'h2a52 	:	val_out <= 4'hee4a;
         4'h2a53 	:	val_out <= 4'hee4a;
         4'h2a58 	:	val_out <= 4'hee57;
         4'h2a59 	:	val_out <= 4'hee57;
         4'h2a5a 	:	val_out <= 4'hee57;
         4'h2a5b 	:	val_out <= 4'hee57;
         4'h2a60 	:	val_out <= 4'hee63;
         4'h2a61 	:	val_out <= 4'hee63;
         4'h2a62 	:	val_out <= 4'hee63;
         4'h2a63 	:	val_out <= 4'hee63;
         4'h2a68 	:	val_out <= 4'hee70;
         4'h2a69 	:	val_out <= 4'hee70;
         4'h2a6a 	:	val_out <= 4'hee70;
         4'h2a6b 	:	val_out <= 4'hee70;
         4'h2a70 	:	val_out <= 4'hee7d;
         4'h2a71 	:	val_out <= 4'hee7d;
         4'h2a72 	:	val_out <= 4'hee7d;
         4'h2a73 	:	val_out <= 4'hee7d;
         4'h2a78 	:	val_out <= 4'hee89;
         4'h2a79 	:	val_out <= 4'hee89;
         4'h2a7a 	:	val_out <= 4'hee89;
         4'h2a7b 	:	val_out <= 4'hee89;
         4'h2a80 	:	val_out <= 4'hee96;
         4'h2a81 	:	val_out <= 4'hee96;
         4'h2a82 	:	val_out <= 4'hee96;
         4'h2a83 	:	val_out <= 4'hee96;
         4'h2a88 	:	val_out <= 4'heea3;
         4'h2a89 	:	val_out <= 4'heea3;
         4'h2a8a 	:	val_out <= 4'heea3;
         4'h2a8b 	:	val_out <= 4'heea3;
         4'h2a90 	:	val_out <= 4'heeaf;
         4'h2a91 	:	val_out <= 4'heeaf;
         4'h2a92 	:	val_out <= 4'heeaf;
         4'h2a93 	:	val_out <= 4'heeaf;
         4'h2a98 	:	val_out <= 4'heebc;
         4'h2a99 	:	val_out <= 4'heebc;
         4'h2a9a 	:	val_out <= 4'heebc;
         4'h2a9b 	:	val_out <= 4'heebc;
         4'h2aa0 	:	val_out <= 4'heec9;
         4'h2aa1 	:	val_out <= 4'heec9;
         4'h2aa2 	:	val_out <= 4'heec9;
         4'h2aa3 	:	val_out <= 4'heec9;
         4'h2aa8 	:	val_out <= 4'heed5;
         4'h2aa9 	:	val_out <= 4'heed5;
         4'h2aaa 	:	val_out <= 4'heed5;
         4'h2aab 	:	val_out <= 4'heed5;
         4'h2ab0 	:	val_out <= 4'heee2;
         4'h2ab1 	:	val_out <= 4'heee2;
         4'h2ab2 	:	val_out <= 4'heee2;
         4'h2ab3 	:	val_out <= 4'heee2;
         4'h2ab8 	:	val_out <= 4'heeee;
         4'h2ab9 	:	val_out <= 4'heeee;
         4'h2aba 	:	val_out <= 4'heeee;
         4'h2abb 	:	val_out <= 4'heeee;
         4'h2ac0 	:	val_out <= 4'heefb;
         4'h2ac1 	:	val_out <= 4'heefb;
         4'h2ac2 	:	val_out <= 4'heefb;
         4'h2ac3 	:	val_out <= 4'heefb;
         4'h2ac8 	:	val_out <= 4'hef07;
         4'h2ac9 	:	val_out <= 4'hef07;
         4'h2aca 	:	val_out <= 4'hef07;
         4'h2acb 	:	val_out <= 4'hef07;
         4'h2ad0 	:	val_out <= 4'hef14;
         4'h2ad1 	:	val_out <= 4'hef14;
         4'h2ad2 	:	val_out <= 4'hef14;
         4'h2ad3 	:	val_out <= 4'hef14;
         4'h2ad8 	:	val_out <= 4'hef20;
         4'h2ad9 	:	val_out <= 4'hef20;
         4'h2ada 	:	val_out <= 4'hef20;
         4'h2adb 	:	val_out <= 4'hef20;
         4'h2ae0 	:	val_out <= 4'hef2d;
         4'h2ae1 	:	val_out <= 4'hef2d;
         4'h2ae2 	:	val_out <= 4'hef2d;
         4'h2ae3 	:	val_out <= 4'hef2d;
         4'h2ae8 	:	val_out <= 4'hef39;
         4'h2ae9 	:	val_out <= 4'hef39;
         4'h2aea 	:	val_out <= 4'hef39;
         4'h2aeb 	:	val_out <= 4'hef39;
         4'h2af0 	:	val_out <= 4'hef46;
         4'h2af1 	:	val_out <= 4'hef46;
         4'h2af2 	:	val_out <= 4'hef46;
         4'h2af3 	:	val_out <= 4'hef46;
         4'h2af8 	:	val_out <= 4'hef52;
         4'h2af9 	:	val_out <= 4'hef52;
         4'h2afa 	:	val_out <= 4'hef52;
         4'h2afb 	:	val_out <= 4'hef52;
         4'h2b00 	:	val_out <= 4'hef5f;
         4'h2b01 	:	val_out <= 4'hef5f;
         4'h2b02 	:	val_out <= 4'hef5f;
         4'h2b03 	:	val_out <= 4'hef5f;
         4'h2b08 	:	val_out <= 4'hef6b;
         4'h2b09 	:	val_out <= 4'hef6b;
         4'h2b0a 	:	val_out <= 4'hef6b;
         4'h2b0b 	:	val_out <= 4'hef6b;
         4'h2b10 	:	val_out <= 4'hef77;
         4'h2b11 	:	val_out <= 4'hef77;
         4'h2b12 	:	val_out <= 4'hef77;
         4'h2b13 	:	val_out <= 4'hef77;
         4'h2b18 	:	val_out <= 4'hef84;
         4'h2b19 	:	val_out <= 4'hef84;
         4'h2b1a 	:	val_out <= 4'hef84;
         4'h2b1b 	:	val_out <= 4'hef84;
         4'h2b20 	:	val_out <= 4'hef90;
         4'h2b21 	:	val_out <= 4'hef90;
         4'h2b22 	:	val_out <= 4'hef90;
         4'h2b23 	:	val_out <= 4'hef90;
         4'h2b28 	:	val_out <= 4'hef9c;
         4'h2b29 	:	val_out <= 4'hef9c;
         4'h2b2a 	:	val_out <= 4'hef9c;
         4'h2b2b 	:	val_out <= 4'hef9c;
         4'h2b30 	:	val_out <= 4'hefa9;
         4'h2b31 	:	val_out <= 4'hefa9;
         4'h2b32 	:	val_out <= 4'hefa9;
         4'h2b33 	:	val_out <= 4'hefa9;
         4'h2b38 	:	val_out <= 4'hefb5;
         4'h2b39 	:	val_out <= 4'hefb5;
         4'h2b3a 	:	val_out <= 4'hefb5;
         4'h2b3b 	:	val_out <= 4'hefb5;
         4'h2b40 	:	val_out <= 4'hefc1;
         4'h2b41 	:	val_out <= 4'hefc1;
         4'h2b42 	:	val_out <= 4'hefc1;
         4'h2b43 	:	val_out <= 4'hefc1;
         4'h2b48 	:	val_out <= 4'hefcd;
         4'h2b49 	:	val_out <= 4'hefcd;
         4'h2b4a 	:	val_out <= 4'hefcd;
         4'h2b4b 	:	val_out <= 4'hefcd;
         4'h2b50 	:	val_out <= 4'hefda;
         4'h2b51 	:	val_out <= 4'hefda;
         4'h2b52 	:	val_out <= 4'hefda;
         4'h2b53 	:	val_out <= 4'hefda;
         4'h2b58 	:	val_out <= 4'hefe6;
         4'h2b59 	:	val_out <= 4'hefe6;
         4'h2b5a 	:	val_out <= 4'hefe6;
         4'h2b5b 	:	val_out <= 4'hefe6;
         4'h2b60 	:	val_out <= 4'heff2;
         4'h2b61 	:	val_out <= 4'heff2;
         4'h2b62 	:	val_out <= 4'heff2;
         4'h2b63 	:	val_out <= 4'heff2;
         4'h2b68 	:	val_out <= 4'heffe;
         4'h2b69 	:	val_out <= 4'heffe;
         4'h2b6a 	:	val_out <= 4'heffe;
         4'h2b6b 	:	val_out <= 4'heffe;
         4'h2b70 	:	val_out <= 4'hf00a;
         4'h2b71 	:	val_out <= 4'hf00a;
         4'h2b72 	:	val_out <= 4'hf00a;
         4'h2b73 	:	val_out <= 4'hf00a;
         4'h2b78 	:	val_out <= 4'hf016;
         4'h2b79 	:	val_out <= 4'hf016;
         4'h2b7a 	:	val_out <= 4'hf016;
         4'h2b7b 	:	val_out <= 4'hf016;
         4'h2b80 	:	val_out <= 4'hf023;
         4'h2b81 	:	val_out <= 4'hf023;
         4'h2b82 	:	val_out <= 4'hf023;
         4'h2b83 	:	val_out <= 4'hf023;
         4'h2b88 	:	val_out <= 4'hf02f;
         4'h2b89 	:	val_out <= 4'hf02f;
         4'h2b8a 	:	val_out <= 4'hf02f;
         4'h2b8b 	:	val_out <= 4'hf02f;
         4'h2b90 	:	val_out <= 4'hf03b;
         4'h2b91 	:	val_out <= 4'hf03b;
         4'h2b92 	:	val_out <= 4'hf03b;
         4'h2b93 	:	val_out <= 4'hf03b;
         4'h2b98 	:	val_out <= 4'hf047;
         4'h2b99 	:	val_out <= 4'hf047;
         4'h2b9a 	:	val_out <= 4'hf047;
         4'h2b9b 	:	val_out <= 4'hf047;
         4'h2ba0 	:	val_out <= 4'hf053;
         4'h2ba1 	:	val_out <= 4'hf053;
         4'h2ba2 	:	val_out <= 4'hf053;
         4'h2ba3 	:	val_out <= 4'hf053;
         4'h2ba8 	:	val_out <= 4'hf05f;
         4'h2ba9 	:	val_out <= 4'hf05f;
         4'h2baa 	:	val_out <= 4'hf05f;
         4'h2bab 	:	val_out <= 4'hf05f;
         4'h2bb0 	:	val_out <= 4'hf06b;
         4'h2bb1 	:	val_out <= 4'hf06b;
         4'h2bb2 	:	val_out <= 4'hf06b;
         4'h2bb3 	:	val_out <= 4'hf06b;
         4'h2bb8 	:	val_out <= 4'hf077;
         4'h2bb9 	:	val_out <= 4'hf077;
         4'h2bba 	:	val_out <= 4'hf077;
         4'h2bbb 	:	val_out <= 4'hf077;
         4'h2bc0 	:	val_out <= 4'hf083;
         4'h2bc1 	:	val_out <= 4'hf083;
         4'h2bc2 	:	val_out <= 4'hf083;
         4'h2bc3 	:	val_out <= 4'hf083;
         4'h2bc8 	:	val_out <= 4'hf08f;
         4'h2bc9 	:	val_out <= 4'hf08f;
         4'h2bca 	:	val_out <= 4'hf08f;
         4'h2bcb 	:	val_out <= 4'hf08f;
         4'h2bd0 	:	val_out <= 4'hf09b;
         4'h2bd1 	:	val_out <= 4'hf09b;
         4'h2bd2 	:	val_out <= 4'hf09b;
         4'h2bd3 	:	val_out <= 4'hf09b;
         4'h2bd8 	:	val_out <= 4'hf0a7;
         4'h2bd9 	:	val_out <= 4'hf0a7;
         4'h2bda 	:	val_out <= 4'hf0a7;
         4'h2bdb 	:	val_out <= 4'hf0a7;
         4'h2be0 	:	val_out <= 4'hf0b3;
         4'h2be1 	:	val_out <= 4'hf0b3;
         4'h2be2 	:	val_out <= 4'hf0b3;
         4'h2be3 	:	val_out <= 4'hf0b3;
         4'h2be8 	:	val_out <= 4'hf0bf;
         4'h2be9 	:	val_out <= 4'hf0bf;
         4'h2bea 	:	val_out <= 4'hf0bf;
         4'h2beb 	:	val_out <= 4'hf0bf;
         4'h2bf0 	:	val_out <= 4'hf0cb;
         4'h2bf1 	:	val_out <= 4'hf0cb;
         4'h2bf2 	:	val_out <= 4'hf0cb;
         4'h2bf3 	:	val_out <= 4'hf0cb;
         4'h2bf8 	:	val_out <= 4'hf0d6;
         4'h2bf9 	:	val_out <= 4'hf0d6;
         4'h2bfa 	:	val_out <= 4'hf0d6;
         4'h2bfb 	:	val_out <= 4'hf0d6;
         4'h2c00 	:	val_out <= 4'hf0e2;
         4'h2c01 	:	val_out <= 4'hf0e2;
         4'h2c02 	:	val_out <= 4'hf0e2;
         4'h2c03 	:	val_out <= 4'hf0e2;
         4'h2c08 	:	val_out <= 4'hf0ee;
         4'h2c09 	:	val_out <= 4'hf0ee;
         4'h2c0a 	:	val_out <= 4'hf0ee;
         4'h2c0b 	:	val_out <= 4'hf0ee;
         4'h2c10 	:	val_out <= 4'hf0fa;
         4'h2c11 	:	val_out <= 4'hf0fa;
         4'h2c12 	:	val_out <= 4'hf0fa;
         4'h2c13 	:	val_out <= 4'hf0fa;
         4'h2c18 	:	val_out <= 4'hf106;
         4'h2c19 	:	val_out <= 4'hf106;
         4'h2c1a 	:	val_out <= 4'hf106;
         4'h2c1b 	:	val_out <= 4'hf106;
         4'h2c20 	:	val_out <= 4'hf112;
         4'h2c21 	:	val_out <= 4'hf112;
         4'h2c22 	:	val_out <= 4'hf112;
         4'h2c23 	:	val_out <= 4'hf112;
         4'h2c28 	:	val_out <= 4'hf11d;
         4'h2c29 	:	val_out <= 4'hf11d;
         4'h2c2a 	:	val_out <= 4'hf11d;
         4'h2c2b 	:	val_out <= 4'hf11d;
         4'h2c30 	:	val_out <= 4'hf129;
         4'h2c31 	:	val_out <= 4'hf129;
         4'h2c32 	:	val_out <= 4'hf129;
         4'h2c33 	:	val_out <= 4'hf129;
         4'h2c38 	:	val_out <= 4'hf135;
         4'h2c39 	:	val_out <= 4'hf135;
         4'h2c3a 	:	val_out <= 4'hf135;
         4'h2c3b 	:	val_out <= 4'hf135;
         4'h2c40 	:	val_out <= 4'hf141;
         4'h2c41 	:	val_out <= 4'hf141;
         4'h2c42 	:	val_out <= 4'hf141;
         4'h2c43 	:	val_out <= 4'hf141;
         4'h2c48 	:	val_out <= 4'hf14c;
         4'h2c49 	:	val_out <= 4'hf14c;
         4'h2c4a 	:	val_out <= 4'hf14c;
         4'h2c4b 	:	val_out <= 4'hf14c;
         4'h2c50 	:	val_out <= 4'hf158;
         4'h2c51 	:	val_out <= 4'hf158;
         4'h2c52 	:	val_out <= 4'hf158;
         4'h2c53 	:	val_out <= 4'hf158;
         4'h2c58 	:	val_out <= 4'hf164;
         4'h2c59 	:	val_out <= 4'hf164;
         4'h2c5a 	:	val_out <= 4'hf164;
         4'h2c5b 	:	val_out <= 4'hf164;
         4'h2c60 	:	val_out <= 4'hf16f;
         4'h2c61 	:	val_out <= 4'hf16f;
         4'h2c62 	:	val_out <= 4'hf16f;
         4'h2c63 	:	val_out <= 4'hf16f;
         4'h2c68 	:	val_out <= 4'hf17b;
         4'h2c69 	:	val_out <= 4'hf17b;
         4'h2c6a 	:	val_out <= 4'hf17b;
         4'h2c6b 	:	val_out <= 4'hf17b;
         4'h2c70 	:	val_out <= 4'hf186;
         4'h2c71 	:	val_out <= 4'hf186;
         4'h2c72 	:	val_out <= 4'hf186;
         4'h2c73 	:	val_out <= 4'hf186;
         4'h2c78 	:	val_out <= 4'hf192;
         4'h2c79 	:	val_out <= 4'hf192;
         4'h2c7a 	:	val_out <= 4'hf192;
         4'h2c7b 	:	val_out <= 4'hf192;
         4'h2c80 	:	val_out <= 4'hf19e;
         4'h2c81 	:	val_out <= 4'hf19e;
         4'h2c82 	:	val_out <= 4'hf19e;
         4'h2c83 	:	val_out <= 4'hf19e;
         4'h2c88 	:	val_out <= 4'hf1a9;
         4'h2c89 	:	val_out <= 4'hf1a9;
         4'h2c8a 	:	val_out <= 4'hf1a9;
         4'h2c8b 	:	val_out <= 4'hf1a9;
         4'h2c90 	:	val_out <= 4'hf1b5;
         4'h2c91 	:	val_out <= 4'hf1b5;
         4'h2c92 	:	val_out <= 4'hf1b5;
         4'h2c93 	:	val_out <= 4'hf1b5;
         4'h2c98 	:	val_out <= 4'hf1c0;
         4'h2c99 	:	val_out <= 4'hf1c0;
         4'h2c9a 	:	val_out <= 4'hf1c0;
         4'h2c9b 	:	val_out <= 4'hf1c0;
         4'h2ca0 	:	val_out <= 4'hf1cc;
         4'h2ca1 	:	val_out <= 4'hf1cc;
         4'h2ca2 	:	val_out <= 4'hf1cc;
         4'h2ca3 	:	val_out <= 4'hf1cc;
         4'h2ca8 	:	val_out <= 4'hf1d7;
         4'h2ca9 	:	val_out <= 4'hf1d7;
         4'h2caa 	:	val_out <= 4'hf1d7;
         4'h2cab 	:	val_out <= 4'hf1d7;
         4'h2cb0 	:	val_out <= 4'hf1e3;
         4'h2cb1 	:	val_out <= 4'hf1e3;
         4'h2cb2 	:	val_out <= 4'hf1e3;
         4'h2cb3 	:	val_out <= 4'hf1e3;
         4'h2cb8 	:	val_out <= 4'hf1ee;
         4'h2cb9 	:	val_out <= 4'hf1ee;
         4'h2cba 	:	val_out <= 4'hf1ee;
         4'h2cbb 	:	val_out <= 4'hf1ee;
         4'h2cc0 	:	val_out <= 4'hf1fa;
         4'h2cc1 	:	val_out <= 4'hf1fa;
         4'h2cc2 	:	val_out <= 4'hf1fa;
         4'h2cc3 	:	val_out <= 4'hf1fa;
         4'h2cc8 	:	val_out <= 4'hf205;
         4'h2cc9 	:	val_out <= 4'hf205;
         4'h2cca 	:	val_out <= 4'hf205;
         4'h2ccb 	:	val_out <= 4'hf205;
         4'h2cd0 	:	val_out <= 4'hf211;
         4'h2cd1 	:	val_out <= 4'hf211;
         4'h2cd2 	:	val_out <= 4'hf211;
         4'h2cd3 	:	val_out <= 4'hf211;
         4'h2cd8 	:	val_out <= 4'hf21c;
         4'h2cd9 	:	val_out <= 4'hf21c;
         4'h2cda 	:	val_out <= 4'hf21c;
         4'h2cdb 	:	val_out <= 4'hf21c;
         4'h2ce0 	:	val_out <= 4'hf227;
         4'h2ce1 	:	val_out <= 4'hf227;
         4'h2ce2 	:	val_out <= 4'hf227;
         4'h2ce3 	:	val_out <= 4'hf227;
         4'h2ce8 	:	val_out <= 4'hf233;
         4'h2ce9 	:	val_out <= 4'hf233;
         4'h2cea 	:	val_out <= 4'hf233;
         4'h2ceb 	:	val_out <= 4'hf233;
         4'h2cf0 	:	val_out <= 4'hf23e;
         4'h2cf1 	:	val_out <= 4'hf23e;
         4'h2cf2 	:	val_out <= 4'hf23e;
         4'h2cf3 	:	val_out <= 4'hf23e;
         4'h2cf8 	:	val_out <= 4'hf249;
         4'h2cf9 	:	val_out <= 4'hf249;
         4'h2cfa 	:	val_out <= 4'hf249;
         4'h2cfb 	:	val_out <= 4'hf249;
         4'h2d00 	:	val_out <= 4'hf255;
         4'h2d01 	:	val_out <= 4'hf255;
         4'h2d02 	:	val_out <= 4'hf255;
         4'h2d03 	:	val_out <= 4'hf255;
         4'h2d08 	:	val_out <= 4'hf260;
         4'h2d09 	:	val_out <= 4'hf260;
         4'h2d0a 	:	val_out <= 4'hf260;
         4'h2d0b 	:	val_out <= 4'hf260;
         4'h2d10 	:	val_out <= 4'hf26b;
         4'h2d11 	:	val_out <= 4'hf26b;
         4'h2d12 	:	val_out <= 4'hf26b;
         4'h2d13 	:	val_out <= 4'hf26b;
         4'h2d18 	:	val_out <= 4'hf276;
         4'h2d19 	:	val_out <= 4'hf276;
         4'h2d1a 	:	val_out <= 4'hf276;
         4'h2d1b 	:	val_out <= 4'hf276;
         4'h2d20 	:	val_out <= 4'hf282;
         4'h2d21 	:	val_out <= 4'hf282;
         4'h2d22 	:	val_out <= 4'hf282;
         4'h2d23 	:	val_out <= 4'hf282;
         4'h2d28 	:	val_out <= 4'hf28d;
         4'h2d29 	:	val_out <= 4'hf28d;
         4'h2d2a 	:	val_out <= 4'hf28d;
         4'h2d2b 	:	val_out <= 4'hf28d;
         4'h2d30 	:	val_out <= 4'hf298;
         4'h2d31 	:	val_out <= 4'hf298;
         4'h2d32 	:	val_out <= 4'hf298;
         4'h2d33 	:	val_out <= 4'hf298;
         4'h2d38 	:	val_out <= 4'hf2a3;
         4'h2d39 	:	val_out <= 4'hf2a3;
         4'h2d3a 	:	val_out <= 4'hf2a3;
         4'h2d3b 	:	val_out <= 4'hf2a3;
         4'h2d40 	:	val_out <= 4'hf2af;
         4'h2d41 	:	val_out <= 4'hf2af;
         4'h2d42 	:	val_out <= 4'hf2af;
         4'h2d43 	:	val_out <= 4'hf2af;
         4'h2d48 	:	val_out <= 4'hf2ba;
         4'h2d49 	:	val_out <= 4'hf2ba;
         4'h2d4a 	:	val_out <= 4'hf2ba;
         4'h2d4b 	:	val_out <= 4'hf2ba;
         4'h2d50 	:	val_out <= 4'hf2c5;
         4'h2d51 	:	val_out <= 4'hf2c5;
         4'h2d52 	:	val_out <= 4'hf2c5;
         4'h2d53 	:	val_out <= 4'hf2c5;
         4'h2d58 	:	val_out <= 4'hf2d0;
         4'h2d59 	:	val_out <= 4'hf2d0;
         4'h2d5a 	:	val_out <= 4'hf2d0;
         4'h2d5b 	:	val_out <= 4'hf2d0;
         4'h2d60 	:	val_out <= 4'hf2db;
         4'h2d61 	:	val_out <= 4'hf2db;
         4'h2d62 	:	val_out <= 4'hf2db;
         4'h2d63 	:	val_out <= 4'hf2db;
         4'h2d68 	:	val_out <= 4'hf2e6;
         4'h2d69 	:	val_out <= 4'hf2e6;
         4'h2d6a 	:	val_out <= 4'hf2e6;
         4'h2d6b 	:	val_out <= 4'hf2e6;
         4'h2d70 	:	val_out <= 4'hf2f1;
         4'h2d71 	:	val_out <= 4'hf2f1;
         4'h2d72 	:	val_out <= 4'hf2f1;
         4'h2d73 	:	val_out <= 4'hf2f1;
         4'h2d78 	:	val_out <= 4'hf2fc;
         4'h2d79 	:	val_out <= 4'hf2fc;
         4'h2d7a 	:	val_out <= 4'hf2fc;
         4'h2d7b 	:	val_out <= 4'hf2fc;
         4'h2d80 	:	val_out <= 4'hf307;
         4'h2d81 	:	val_out <= 4'hf307;
         4'h2d82 	:	val_out <= 4'hf307;
         4'h2d83 	:	val_out <= 4'hf307;
         4'h2d88 	:	val_out <= 4'hf312;
         4'h2d89 	:	val_out <= 4'hf312;
         4'h2d8a 	:	val_out <= 4'hf312;
         4'h2d8b 	:	val_out <= 4'hf312;
         4'h2d90 	:	val_out <= 4'hf31d;
         4'h2d91 	:	val_out <= 4'hf31d;
         4'h2d92 	:	val_out <= 4'hf31d;
         4'h2d93 	:	val_out <= 4'hf31d;
         4'h2d98 	:	val_out <= 4'hf328;
         4'h2d99 	:	val_out <= 4'hf328;
         4'h2d9a 	:	val_out <= 4'hf328;
         4'h2d9b 	:	val_out <= 4'hf328;
         4'h2da0 	:	val_out <= 4'hf333;
         4'h2da1 	:	val_out <= 4'hf333;
         4'h2da2 	:	val_out <= 4'hf333;
         4'h2da3 	:	val_out <= 4'hf333;
         4'h2da8 	:	val_out <= 4'hf33e;
         4'h2da9 	:	val_out <= 4'hf33e;
         4'h2daa 	:	val_out <= 4'hf33e;
         4'h2dab 	:	val_out <= 4'hf33e;
         4'h2db0 	:	val_out <= 4'hf349;
         4'h2db1 	:	val_out <= 4'hf349;
         4'h2db2 	:	val_out <= 4'hf349;
         4'h2db3 	:	val_out <= 4'hf349;
         4'h2db8 	:	val_out <= 4'hf354;
         4'h2db9 	:	val_out <= 4'hf354;
         4'h2dba 	:	val_out <= 4'hf354;
         4'h2dbb 	:	val_out <= 4'hf354;
         4'h2dc0 	:	val_out <= 4'hf35f;
         4'h2dc1 	:	val_out <= 4'hf35f;
         4'h2dc2 	:	val_out <= 4'hf35f;
         4'h2dc3 	:	val_out <= 4'hf35f;
         4'h2dc8 	:	val_out <= 4'hf36a;
         4'h2dc9 	:	val_out <= 4'hf36a;
         4'h2dca 	:	val_out <= 4'hf36a;
         4'h2dcb 	:	val_out <= 4'hf36a;
         4'h2dd0 	:	val_out <= 4'hf375;
         4'h2dd1 	:	val_out <= 4'hf375;
         4'h2dd2 	:	val_out <= 4'hf375;
         4'h2dd3 	:	val_out <= 4'hf375;
         4'h2dd8 	:	val_out <= 4'hf37f;
         4'h2dd9 	:	val_out <= 4'hf37f;
         4'h2dda 	:	val_out <= 4'hf37f;
         4'h2ddb 	:	val_out <= 4'hf37f;
         4'h2de0 	:	val_out <= 4'hf38a;
         4'h2de1 	:	val_out <= 4'hf38a;
         4'h2de2 	:	val_out <= 4'hf38a;
         4'h2de3 	:	val_out <= 4'hf38a;
         4'h2de8 	:	val_out <= 4'hf395;
         4'h2de9 	:	val_out <= 4'hf395;
         4'h2dea 	:	val_out <= 4'hf395;
         4'h2deb 	:	val_out <= 4'hf395;
         4'h2df0 	:	val_out <= 4'hf3a0;
         4'h2df1 	:	val_out <= 4'hf3a0;
         4'h2df2 	:	val_out <= 4'hf3a0;
         4'h2df3 	:	val_out <= 4'hf3a0;
         4'h2df8 	:	val_out <= 4'hf3ab;
         4'h2df9 	:	val_out <= 4'hf3ab;
         4'h2dfa 	:	val_out <= 4'hf3ab;
         4'h2dfb 	:	val_out <= 4'hf3ab;
         4'h2e00 	:	val_out <= 4'hf3b5;
         4'h2e01 	:	val_out <= 4'hf3b5;
         4'h2e02 	:	val_out <= 4'hf3b5;
         4'h2e03 	:	val_out <= 4'hf3b5;
         4'h2e08 	:	val_out <= 4'hf3c0;
         4'h2e09 	:	val_out <= 4'hf3c0;
         4'h2e0a 	:	val_out <= 4'hf3c0;
         4'h2e0b 	:	val_out <= 4'hf3c0;
         4'h2e10 	:	val_out <= 4'hf3cb;
         4'h2e11 	:	val_out <= 4'hf3cb;
         4'h2e12 	:	val_out <= 4'hf3cb;
         4'h2e13 	:	val_out <= 4'hf3cb;
         4'h2e18 	:	val_out <= 4'hf3d6;
         4'h2e19 	:	val_out <= 4'hf3d6;
         4'h2e1a 	:	val_out <= 4'hf3d6;
         4'h2e1b 	:	val_out <= 4'hf3d6;
         4'h2e20 	:	val_out <= 4'hf3e0;
         4'h2e21 	:	val_out <= 4'hf3e0;
         4'h2e22 	:	val_out <= 4'hf3e0;
         4'h2e23 	:	val_out <= 4'hf3e0;
         4'h2e28 	:	val_out <= 4'hf3eb;
         4'h2e29 	:	val_out <= 4'hf3eb;
         4'h2e2a 	:	val_out <= 4'hf3eb;
         4'h2e2b 	:	val_out <= 4'hf3eb;
         4'h2e30 	:	val_out <= 4'hf3f6;
         4'h2e31 	:	val_out <= 4'hf3f6;
         4'h2e32 	:	val_out <= 4'hf3f6;
         4'h2e33 	:	val_out <= 4'hf3f6;
         4'h2e38 	:	val_out <= 4'hf400;
         4'h2e39 	:	val_out <= 4'hf400;
         4'h2e3a 	:	val_out <= 4'hf400;
         4'h2e3b 	:	val_out <= 4'hf400;
         4'h2e40 	:	val_out <= 4'hf40b;
         4'h2e41 	:	val_out <= 4'hf40b;
         4'h2e42 	:	val_out <= 4'hf40b;
         4'h2e43 	:	val_out <= 4'hf40b;
         4'h2e48 	:	val_out <= 4'hf415;
         4'h2e49 	:	val_out <= 4'hf415;
         4'h2e4a 	:	val_out <= 4'hf415;
         4'h2e4b 	:	val_out <= 4'hf415;
         4'h2e50 	:	val_out <= 4'hf420;
         4'h2e51 	:	val_out <= 4'hf420;
         4'h2e52 	:	val_out <= 4'hf420;
         4'h2e53 	:	val_out <= 4'hf420;
         4'h2e58 	:	val_out <= 4'hf42b;
         4'h2e59 	:	val_out <= 4'hf42b;
         4'h2e5a 	:	val_out <= 4'hf42b;
         4'h2e5b 	:	val_out <= 4'hf42b;
         4'h2e60 	:	val_out <= 4'hf435;
         4'h2e61 	:	val_out <= 4'hf435;
         4'h2e62 	:	val_out <= 4'hf435;
         4'h2e63 	:	val_out <= 4'hf435;
         4'h2e68 	:	val_out <= 4'hf440;
         4'h2e69 	:	val_out <= 4'hf440;
         4'h2e6a 	:	val_out <= 4'hf440;
         4'h2e6b 	:	val_out <= 4'hf440;
         4'h2e70 	:	val_out <= 4'hf44a;
         4'h2e71 	:	val_out <= 4'hf44a;
         4'h2e72 	:	val_out <= 4'hf44a;
         4'h2e73 	:	val_out <= 4'hf44a;
         4'h2e78 	:	val_out <= 4'hf455;
         4'h2e79 	:	val_out <= 4'hf455;
         4'h2e7a 	:	val_out <= 4'hf455;
         4'h2e7b 	:	val_out <= 4'hf455;
         4'h2e80 	:	val_out <= 4'hf45f;
         4'h2e81 	:	val_out <= 4'hf45f;
         4'h2e82 	:	val_out <= 4'hf45f;
         4'h2e83 	:	val_out <= 4'hf45f;
         4'h2e88 	:	val_out <= 4'hf46a;
         4'h2e89 	:	val_out <= 4'hf46a;
         4'h2e8a 	:	val_out <= 4'hf46a;
         4'h2e8b 	:	val_out <= 4'hf46a;
         4'h2e90 	:	val_out <= 4'hf474;
         4'h2e91 	:	val_out <= 4'hf474;
         4'h2e92 	:	val_out <= 4'hf474;
         4'h2e93 	:	val_out <= 4'hf474;
         4'h2e98 	:	val_out <= 4'hf47e;
         4'h2e99 	:	val_out <= 4'hf47e;
         4'h2e9a 	:	val_out <= 4'hf47e;
         4'h2e9b 	:	val_out <= 4'hf47e;
         4'h2ea0 	:	val_out <= 4'hf489;
         4'h2ea1 	:	val_out <= 4'hf489;
         4'h2ea2 	:	val_out <= 4'hf489;
         4'h2ea3 	:	val_out <= 4'hf489;
         4'h2ea8 	:	val_out <= 4'hf493;
         4'h2ea9 	:	val_out <= 4'hf493;
         4'h2eaa 	:	val_out <= 4'hf493;
         4'h2eab 	:	val_out <= 4'hf493;
         4'h2eb0 	:	val_out <= 4'hf49e;
         4'h2eb1 	:	val_out <= 4'hf49e;
         4'h2eb2 	:	val_out <= 4'hf49e;
         4'h2eb3 	:	val_out <= 4'hf49e;
         4'h2eb8 	:	val_out <= 4'hf4a8;
         4'h2eb9 	:	val_out <= 4'hf4a8;
         4'h2eba 	:	val_out <= 4'hf4a8;
         4'h2ebb 	:	val_out <= 4'hf4a8;
         4'h2ec0 	:	val_out <= 4'hf4b2;
         4'h2ec1 	:	val_out <= 4'hf4b2;
         4'h2ec2 	:	val_out <= 4'hf4b2;
         4'h2ec3 	:	val_out <= 4'hf4b2;
         4'h2ec8 	:	val_out <= 4'hf4bd;
         4'h2ec9 	:	val_out <= 4'hf4bd;
         4'h2eca 	:	val_out <= 4'hf4bd;
         4'h2ecb 	:	val_out <= 4'hf4bd;
         4'h2ed0 	:	val_out <= 4'hf4c7;
         4'h2ed1 	:	val_out <= 4'hf4c7;
         4'h2ed2 	:	val_out <= 4'hf4c7;
         4'h2ed3 	:	val_out <= 4'hf4c7;
         4'h2ed8 	:	val_out <= 4'hf4d1;
         4'h2ed9 	:	val_out <= 4'hf4d1;
         4'h2eda 	:	val_out <= 4'hf4d1;
         4'h2edb 	:	val_out <= 4'hf4d1;
         4'h2ee0 	:	val_out <= 4'hf4db;
         4'h2ee1 	:	val_out <= 4'hf4db;
         4'h2ee2 	:	val_out <= 4'hf4db;
         4'h2ee3 	:	val_out <= 4'hf4db;
         4'h2ee8 	:	val_out <= 4'hf4e6;
         4'h2ee9 	:	val_out <= 4'hf4e6;
         4'h2eea 	:	val_out <= 4'hf4e6;
         4'h2eeb 	:	val_out <= 4'hf4e6;
         4'h2ef0 	:	val_out <= 4'hf4f0;
         4'h2ef1 	:	val_out <= 4'hf4f0;
         4'h2ef2 	:	val_out <= 4'hf4f0;
         4'h2ef3 	:	val_out <= 4'hf4f0;
         4'h2ef8 	:	val_out <= 4'hf4fa;
         4'h2ef9 	:	val_out <= 4'hf4fa;
         4'h2efa 	:	val_out <= 4'hf4fa;
         4'h2efb 	:	val_out <= 4'hf4fa;
         4'h2f00 	:	val_out <= 4'hf504;
         4'h2f01 	:	val_out <= 4'hf504;
         4'h2f02 	:	val_out <= 4'hf504;
         4'h2f03 	:	val_out <= 4'hf504;
         4'h2f08 	:	val_out <= 4'hf50f;
         4'h2f09 	:	val_out <= 4'hf50f;
         4'h2f0a 	:	val_out <= 4'hf50f;
         4'h2f0b 	:	val_out <= 4'hf50f;
         4'h2f10 	:	val_out <= 4'hf519;
         4'h2f11 	:	val_out <= 4'hf519;
         4'h2f12 	:	val_out <= 4'hf519;
         4'h2f13 	:	val_out <= 4'hf519;
         4'h2f18 	:	val_out <= 4'hf523;
         4'h2f19 	:	val_out <= 4'hf523;
         4'h2f1a 	:	val_out <= 4'hf523;
         4'h2f1b 	:	val_out <= 4'hf523;
         4'h2f20 	:	val_out <= 4'hf52d;
         4'h2f21 	:	val_out <= 4'hf52d;
         4'h2f22 	:	val_out <= 4'hf52d;
         4'h2f23 	:	val_out <= 4'hf52d;
         4'h2f28 	:	val_out <= 4'hf537;
         4'h2f29 	:	val_out <= 4'hf537;
         4'h2f2a 	:	val_out <= 4'hf537;
         4'h2f2b 	:	val_out <= 4'hf537;
         4'h2f30 	:	val_out <= 4'hf541;
         4'h2f31 	:	val_out <= 4'hf541;
         4'h2f32 	:	val_out <= 4'hf541;
         4'h2f33 	:	val_out <= 4'hf541;
         4'h2f38 	:	val_out <= 4'hf54b;
         4'h2f39 	:	val_out <= 4'hf54b;
         4'h2f3a 	:	val_out <= 4'hf54b;
         4'h2f3b 	:	val_out <= 4'hf54b;
         4'h2f40 	:	val_out <= 4'hf555;
         4'h2f41 	:	val_out <= 4'hf555;
         4'h2f42 	:	val_out <= 4'hf555;
         4'h2f43 	:	val_out <= 4'hf555;
         4'h2f48 	:	val_out <= 4'hf55f;
         4'h2f49 	:	val_out <= 4'hf55f;
         4'h2f4a 	:	val_out <= 4'hf55f;
         4'h2f4b 	:	val_out <= 4'hf55f;
         4'h2f50 	:	val_out <= 4'hf569;
         4'h2f51 	:	val_out <= 4'hf569;
         4'h2f52 	:	val_out <= 4'hf569;
         4'h2f53 	:	val_out <= 4'hf569;
         4'h2f58 	:	val_out <= 4'hf573;
         4'h2f59 	:	val_out <= 4'hf573;
         4'h2f5a 	:	val_out <= 4'hf573;
         4'h2f5b 	:	val_out <= 4'hf573;
         4'h2f60 	:	val_out <= 4'hf57d;
         4'h2f61 	:	val_out <= 4'hf57d;
         4'h2f62 	:	val_out <= 4'hf57d;
         4'h2f63 	:	val_out <= 4'hf57d;
         4'h2f68 	:	val_out <= 4'hf587;
         4'h2f69 	:	val_out <= 4'hf587;
         4'h2f6a 	:	val_out <= 4'hf587;
         4'h2f6b 	:	val_out <= 4'hf587;
         4'h2f70 	:	val_out <= 4'hf591;
         4'h2f71 	:	val_out <= 4'hf591;
         4'h2f72 	:	val_out <= 4'hf591;
         4'h2f73 	:	val_out <= 4'hf591;
         4'h2f78 	:	val_out <= 4'hf59b;
         4'h2f79 	:	val_out <= 4'hf59b;
         4'h2f7a 	:	val_out <= 4'hf59b;
         4'h2f7b 	:	val_out <= 4'hf59b;
         4'h2f80 	:	val_out <= 4'hf5a5;
         4'h2f81 	:	val_out <= 4'hf5a5;
         4'h2f82 	:	val_out <= 4'hf5a5;
         4'h2f83 	:	val_out <= 4'hf5a5;
         4'h2f88 	:	val_out <= 4'hf5af;
         4'h2f89 	:	val_out <= 4'hf5af;
         4'h2f8a 	:	val_out <= 4'hf5af;
         4'h2f8b 	:	val_out <= 4'hf5af;
         4'h2f90 	:	val_out <= 4'hf5b9;
         4'h2f91 	:	val_out <= 4'hf5b9;
         4'h2f92 	:	val_out <= 4'hf5b9;
         4'h2f93 	:	val_out <= 4'hf5b9;
         4'h2f98 	:	val_out <= 4'hf5c3;
         4'h2f99 	:	val_out <= 4'hf5c3;
         4'h2f9a 	:	val_out <= 4'hf5c3;
         4'h2f9b 	:	val_out <= 4'hf5c3;
         4'h2fa0 	:	val_out <= 4'hf5cc;
         4'h2fa1 	:	val_out <= 4'hf5cc;
         4'h2fa2 	:	val_out <= 4'hf5cc;
         4'h2fa3 	:	val_out <= 4'hf5cc;
         4'h2fa8 	:	val_out <= 4'hf5d6;
         4'h2fa9 	:	val_out <= 4'hf5d6;
         4'h2faa 	:	val_out <= 4'hf5d6;
         4'h2fab 	:	val_out <= 4'hf5d6;
         4'h2fb0 	:	val_out <= 4'hf5e0;
         4'h2fb1 	:	val_out <= 4'hf5e0;
         4'h2fb2 	:	val_out <= 4'hf5e0;
         4'h2fb3 	:	val_out <= 4'hf5e0;
         4'h2fb8 	:	val_out <= 4'hf5ea;
         4'h2fb9 	:	val_out <= 4'hf5ea;
         4'h2fba 	:	val_out <= 4'hf5ea;
         4'h2fbb 	:	val_out <= 4'hf5ea;
         4'h2fc0 	:	val_out <= 4'hf5f4;
         4'h2fc1 	:	val_out <= 4'hf5f4;
         4'h2fc2 	:	val_out <= 4'hf5f4;
         4'h2fc3 	:	val_out <= 4'hf5f4;
         4'h2fc8 	:	val_out <= 4'hf5fd;
         4'h2fc9 	:	val_out <= 4'hf5fd;
         4'h2fca 	:	val_out <= 4'hf5fd;
         4'h2fcb 	:	val_out <= 4'hf5fd;
         4'h2fd0 	:	val_out <= 4'hf607;
         4'h2fd1 	:	val_out <= 4'hf607;
         4'h2fd2 	:	val_out <= 4'hf607;
         4'h2fd3 	:	val_out <= 4'hf607;
         4'h2fd8 	:	val_out <= 4'hf611;
         4'h2fd9 	:	val_out <= 4'hf611;
         4'h2fda 	:	val_out <= 4'hf611;
         4'h2fdb 	:	val_out <= 4'hf611;
         4'h2fe0 	:	val_out <= 4'hf61b;
         4'h2fe1 	:	val_out <= 4'hf61b;
         4'h2fe2 	:	val_out <= 4'hf61b;
         4'h2fe3 	:	val_out <= 4'hf61b;
         4'h2fe8 	:	val_out <= 4'hf624;
         4'h2fe9 	:	val_out <= 4'hf624;
         4'h2fea 	:	val_out <= 4'hf624;
         4'h2feb 	:	val_out <= 4'hf624;
         4'h2ff0 	:	val_out <= 4'hf62e;
         4'h2ff1 	:	val_out <= 4'hf62e;
         4'h2ff2 	:	val_out <= 4'hf62e;
         4'h2ff3 	:	val_out <= 4'hf62e;
         4'h2ff8 	:	val_out <= 4'hf638;
         4'h2ff9 	:	val_out <= 4'hf638;
         4'h2ffa 	:	val_out <= 4'hf638;
         4'h2ffb 	:	val_out <= 4'hf638;
         4'h3000 	:	val_out <= 4'hf641;
         4'h3001 	:	val_out <= 4'hf641;
         4'h3002 	:	val_out <= 4'hf641;
         4'h3003 	:	val_out <= 4'hf641;
         4'h3008 	:	val_out <= 4'hf64b;
         4'h3009 	:	val_out <= 4'hf64b;
         4'h300a 	:	val_out <= 4'hf64b;
         4'h300b 	:	val_out <= 4'hf64b;
         4'h3010 	:	val_out <= 4'hf654;
         4'h3011 	:	val_out <= 4'hf654;
         4'h3012 	:	val_out <= 4'hf654;
         4'h3013 	:	val_out <= 4'hf654;
         4'h3018 	:	val_out <= 4'hf65e;
         4'h3019 	:	val_out <= 4'hf65e;
         4'h301a 	:	val_out <= 4'hf65e;
         4'h301b 	:	val_out <= 4'hf65e;
         4'h3020 	:	val_out <= 4'hf668;
         4'h3021 	:	val_out <= 4'hf668;
         4'h3022 	:	val_out <= 4'hf668;
         4'h3023 	:	val_out <= 4'hf668;
         4'h3028 	:	val_out <= 4'hf671;
         4'h3029 	:	val_out <= 4'hf671;
         4'h302a 	:	val_out <= 4'hf671;
         4'h302b 	:	val_out <= 4'hf671;
         4'h3030 	:	val_out <= 4'hf67b;
         4'h3031 	:	val_out <= 4'hf67b;
         4'h3032 	:	val_out <= 4'hf67b;
         4'h3033 	:	val_out <= 4'hf67b;
         4'h3038 	:	val_out <= 4'hf684;
         4'h3039 	:	val_out <= 4'hf684;
         4'h303a 	:	val_out <= 4'hf684;
         4'h303b 	:	val_out <= 4'hf684;
         4'h3040 	:	val_out <= 4'hf68e;
         4'h3041 	:	val_out <= 4'hf68e;
         4'h3042 	:	val_out <= 4'hf68e;
         4'h3043 	:	val_out <= 4'hf68e;
         4'h3048 	:	val_out <= 4'hf697;
         4'h3049 	:	val_out <= 4'hf697;
         4'h304a 	:	val_out <= 4'hf697;
         4'h304b 	:	val_out <= 4'hf697;
         4'h3050 	:	val_out <= 4'hf6a0;
         4'h3051 	:	val_out <= 4'hf6a0;
         4'h3052 	:	val_out <= 4'hf6a0;
         4'h3053 	:	val_out <= 4'hf6a0;
         4'h3058 	:	val_out <= 4'hf6aa;
         4'h3059 	:	val_out <= 4'hf6aa;
         4'h305a 	:	val_out <= 4'hf6aa;
         4'h305b 	:	val_out <= 4'hf6aa;
         4'h3060 	:	val_out <= 4'hf6b3;
         4'h3061 	:	val_out <= 4'hf6b3;
         4'h3062 	:	val_out <= 4'hf6b3;
         4'h3063 	:	val_out <= 4'hf6b3;
         4'h3068 	:	val_out <= 4'hf6bd;
         4'h3069 	:	val_out <= 4'hf6bd;
         4'h306a 	:	val_out <= 4'hf6bd;
         4'h306b 	:	val_out <= 4'hf6bd;
         4'h3070 	:	val_out <= 4'hf6c6;
         4'h3071 	:	val_out <= 4'hf6c6;
         4'h3072 	:	val_out <= 4'hf6c6;
         4'h3073 	:	val_out <= 4'hf6c6;
         4'h3078 	:	val_out <= 4'hf6cf;
         4'h3079 	:	val_out <= 4'hf6cf;
         4'h307a 	:	val_out <= 4'hf6cf;
         4'h307b 	:	val_out <= 4'hf6cf;
         4'h3080 	:	val_out <= 4'hf6d9;
         4'h3081 	:	val_out <= 4'hf6d9;
         4'h3082 	:	val_out <= 4'hf6d9;
         4'h3083 	:	val_out <= 4'hf6d9;
         4'h3088 	:	val_out <= 4'hf6e2;
         4'h3089 	:	val_out <= 4'hf6e2;
         4'h308a 	:	val_out <= 4'hf6e2;
         4'h308b 	:	val_out <= 4'hf6e2;
         4'h3090 	:	val_out <= 4'hf6eb;
         4'h3091 	:	val_out <= 4'hf6eb;
         4'h3092 	:	val_out <= 4'hf6eb;
         4'h3093 	:	val_out <= 4'hf6eb;
         4'h3098 	:	val_out <= 4'hf6f5;
         4'h3099 	:	val_out <= 4'hf6f5;
         4'h309a 	:	val_out <= 4'hf6f5;
         4'h309b 	:	val_out <= 4'hf6f5;
         4'h30a0 	:	val_out <= 4'hf6fe;
         4'h30a1 	:	val_out <= 4'hf6fe;
         4'h30a2 	:	val_out <= 4'hf6fe;
         4'h30a3 	:	val_out <= 4'hf6fe;
         4'h30a8 	:	val_out <= 4'hf707;
         4'h30a9 	:	val_out <= 4'hf707;
         4'h30aa 	:	val_out <= 4'hf707;
         4'h30ab 	:	val_out <= 4'hf707;
         4'h30b0 	:	val_out <= 4'hf710;
         4'h30b1 	:	val_out <= 4'hf710;
         4'h30b2 	:	val_out <= 4'hf710;
         4'h30b3 	:	val_out <= 4'hf710;
         4'h30b8 	:	val_out <= 4'hf71a;
         4'h30b9 	:	val_out <= 4'hf71a;
         4'h30ba 	:	val_out <= 4'hf71a;
         4'h30bb 	:	val_out <= 4'hf71a;
         4'h30c0 	:	val_out <= 4'hf723;
         4'h30c1 	:	val_out <= 4'hf723;
         4'h30c2 	:	val_out <= 4'hf723;
         4'h30c3 	:	val_out <= 4'hf723;
         4'h30c8 	:	val_out <= 4'hf72c;
         4'h30c9 	:	val_out <= 4'hf72c;
         4'h30ca 	:	val_out <= 4'hf72c;
         4'h30cb 	:	val_out <= 4'hf72c;
         4'h30d0 	:	val_out <= 4'hf735;
         4'h30d1 	:	val_out <= 4'hf735;
         4'h30d2 	:	val_out <= 4'hf735;
         4'h30d3 	:	val_out <= 4'hf735;
         4'h30d8 	:	val_out <= 4'hf73e;
         4'h30d9 	:	val_out <= 4'hf73e;
         4'h30da 	:	val_out <= 4'hf73e;
         4'h30db 	:	val_out <= 4'hf73e;
         4'h30e0 	:	val_out <= 4'hf747;
         4'h30e1 	:	val_out <= 4'hf747;
         4'h30e2 	:	val_out <= 4'hf747;
         4'h30e3 	:	val_out <= 4'hf747;
         4'h30e8 	:	val_out <= 4'hf751;
         4'h30e9 	:	val_out <= 4'hf751;
         4'h30ea 	:	val_out <= 4'hf751;
         4'h30eb 	:	val_out <= 4'hf751;
         4'h30f0 	:	val_out <= 4'hf75a;
         4'h30f1 	:	val_out <= 4'hf75a;
         4'h30f2 	:	val_out <= 4'hf75a;
         4'h30f3 	:	val_out <= 4'hf75a;
         4'h30f8 	:	val_out <= 4'hf763;
         4'h30f9 	:	val_out <= 4'hf763;
         4'h30fa 	:	val_out <= 4'hf763;
         4'h30fb 	:	val_out <= 4'hf763;
         4'h3100 	:	val_out <= 4'hf76c;
         4'h3101 	:	val_out <= 4'hf76c;
         4'h3102 	:	val_out <= 4'hf76c;
         4'h3103 	:	val_out <= 4'hf76c;
         4'h3108 	:	val_out <= 4'hf775;
         4'h3109 	:	val_out <= 4'hf775;
         4'h310a 	:	val_out <= 4'hf775;
         4'h310b 	:	val_out <= 4'hf775;
         4'h3110 	:	val_out <= 4'hf77e;
         4'h3111 	:	val_out <= 4'hf77e;
         4'h3112 	:	val_out <= 4'hf77e;
         4'h3113 	:	val_out <= 4'hf77e;
         4'h3118 	:	val_out <= 4'hf787;
         4'h3119 	:	val_out <= 4'hf787;
         4'h311a 	:	val_out <= 4'hf787;
         4'h311b 	:	val_out <= 4'hf787;
         4'h3120 	:	val_out <= 4'hf790;
         4'h3121 	:	val_out <= 4'hf790;
         4'h3122 	:	val_out <= 4'hf790;
         4'h3123 	:	val_out <= 4'hf790;
         4'h3128 	:	val_out <= 4'hf799;
         4'h3129 	:	val_out <= 4'hf799;
         4'h312a 	:	val_out <= 4'hf799;
         4'h312b 	:	val_out <= 4'hf799;
         4'h3130 	:	val_out <= 4'hf7a2;
         4'h3131 	:	val_out <= 4'hf7a2;
         4'h3132 	:	val_out <= 4'hf7a2;
         4'h3133 	:	val_out <= 4'hf7a2;
         4'h3138 	:	val_out <= 4'hf7ab;
         4'h3139 	:	val_out <= 4'hf7ab;
         4'h313a 	:	val_out <= 4'hf7ab;
         4'h313b 	:	val_out <= 4'hf7ab;
         4'h3140 	:	val_out <= 4'hf7b4;
         4'h3141 	:	val_out <= 4'hf7b4;
         4'h3142 	:	val_out <= 4'hf7b4;
         4'h3143 	:	val_out <= 4'hf7b4;
         4'h3148 	:	val_out <= 4'hf7bc;
         4'h3149 	:	val_out <= 4'hf7bc;
         4'h314a 	:	val_out <= 4'hf7bc;
         4'h314b 	:	val_out <= 4'hf7bc;
         4'h3150 	:	val_out <= 4'hf7c5;
         4'h3151 	:	val_out <= 4'hf7c5;
         4'h3152 	:	val_out <= 4'hf7c5;
         4'h3153 	:	val_out <= 4'hf7c5;
         4'h3158 	:	val_out <= 4'hf7ce;
         4'h3159 	:	val_out <= 4'hf7ce;
         4'h315a 	:	val_out <= 4'hf7ce;
         4'h315b 	:	val_out <= 4'hf7ce;
         4'h3160 	:	val_out <= 4'hf7d7;
         4'h3161 	:	val_out <= 4'hf7d7;
         4'h3162 	:	val_out <= 4'hf7d7;
         4'h3163 	:	val_out <= 4'hf7d7;
         4'h3168 	:	val_out <= 4'hf7e0;
         4'h3169 	:	val_out <= 4'hf7e0;
         4'h316a 	:	val_out <= 4'hf7e0;
         4'h316b 	:	val_out <= 4'hf7e0;
         4'h3170 	:	val_out <= 4'hf7e9;
         4'h3171 	:	val_out <= 4'hf7e9;
         4'h3172 	:	val_out <= 4'hf7e9;
         4'h3173 	:	val_out <= 4'hf7e9;
         4'h3178 	:	val_out <= 4'hf7f1;
         4'h3179 	:	val_out <= 4'hf7f1;
         4'h317a 	:	val_out <= 4'hf7f1;
         4'h317b 	:	val_out <= 4'hf7f1;
         4'h3180 	:	val_out <= 4'hf7fa;
         4'h3181 	:	val_out <= 4'hf7fa;
         4'h3182 	:	val_out <= 4'hf7fa;
         4'h3183 	:	val_out <= 4'hf7fa;
         4'h3188 	:	val_out <= 4'hf803;
         4'h3189 	:	val_out <= 4'hf803;
         4'h318a 	:	val_out <= 4'hf803;
         4'h318b 	:	val_out <= 4'hf803;
         4'h3190 	:	val_out <= 4'hf80c;
         4'h3191 	:	val_out <= 4'hf80c;
         4'h3192 	:	val_out <= 4'hf80c;
         4'h3193 	:	val_out <= 4'hf80c;
         4'h3198 	:	val_out <= 4'hf814;
         4'h3199 	:	val_out <= 4'hf814;
         4'h319a 	:	val_out <= 4'hf814;
         4'h319b 	:	val_out <= 4'hf814;
         4'h31a0 	:	val_out <= 4'hf81d;
         4'h31a1 	:	val_out <= 4'hf81d;
         4'h31a2 	:	val_out <= 4'hf81d;
         4'h31a3 	:	val_out <= 4'hf81d;
         4'h31a8 	:	val_out <= 4'hf826;
         4'h31a9 	:	val_out <= 4'hf826;
         4'h31aa 	:	val_out <= 4'hf826;
         4'h31ab 	:	val_out <= 4'hf826;
         4'h31b0 	:	val_out <= 4'hf82e;
         4'h31b1 	:	val_out <= 4'hf82e;
         4'h31b2 	:	val_out <= 4'hf82e;
         4'h31b3 	:	val_out <= 4'hf82e;
         4'h31b8 	:	val_out <= 4'hf837;
         4'h31b9 	:	val_out <= 4'hf837;
         4'h31ba 	:	val_out <= 4'hf837;
         4'h31bb 	:	val_out <= 4'hf837;
         4'h31c0 	:	val_out <= 4'hf840;
         4'h31c1 	:	val_out <= 4'hf840;
         4'h31c2 	:	val_out <= 4'hf840;
         4'h31c3 	:	val_out <= 4'hf840;
         4'h31c8 	:	val_out <= 4'hf848;
         4'h31c9 	:	val_out <= 4'hf848;
         4'h31ca 	:	val_out <= 4'hf848;
         4'h31cb 	:	val_out <= 4'hf848;
         4'h31d0 	:	val_out <= 4'hf851;
         4'h31d1 	:	val_out <= 4'hf851;
         4'h31d2 	:	val_out <= 4'hf851;
         4'h31d3 	:	val_out <= 4'hf851;
         4'h31d8 	:	val_out <= 4'hf859;
         4'h31d9 	:	val_out <= 4'hf859;
         4'h31da 	:	val_out <= 4'hf859;
         4'h31db 	:	val_out <= 4'hf859;
         4'h31e0 	:	val_out <= 4'hf862;
         4'h31e1 	:	val_out <= 4'hf862;
         4'h31e2 	:	val_out <= 4'hf862;
         4'h31e3 	:	val_out <= 4'hf862;
         4'h31e8 	:	val_out <= 4'hf86b;
         4'h31e9 	:	val_out <= 4'hf86b;
         4'h31ea 	:	val_out <= 4'hf86b;
         4'h31eb 	:	val_out <= 4'hf86b;
         4'h31f0 	:	val_out <= 4'hf873;
         4'h31f1 	:	val_out <= 4'hf873;
         4'h31f2 	:	val_out <= 4'hf873;
         4'h31f3 	:	val_out <= 4'hf873;
         4'h31f8 	:	val_out <= 4'hf87c;
         4'h31f9 	:	val_out <= 4'hf87c;
         4'h31fa 	:	val_out <= 4'hf87c;
         4'h31fb 	:	val_out <= 4'hf87c;
         4'h3200 	:	val_out <= 4'hf884;
         4'h3201 	:	val_out <= 4'hf884;
         4'h3202 	:	val_out <= 4'hf884;
         4'h3203 	:	val_out <= 4'hf884;
         4'h3208 	:	val_out <= 4'hf88c;
         4'h3209 	:	val_out <= 4'hf88c;
         4'h320a 	:	val_out <= 4'hf88c;
         4'h320b 	:	val_out <= 4'hf88c;
         4'h3210 	:	val_out <= 4'hf895;
         4'h3211 	:	val_out <= 4'hf895;
         4'h3212 	:	val_out <= 4'hf895;
         4'h3213 	:	val_out <= 4'hf895;
         4'h3218 	:	val_out <= 4'hf89d;
         4'h3219 	:	val_out <= 4'hf89d;
         4'h321a 	:	val_out <= 4'hf89d;
         4'h321b 	:	val_out <= 4'hf89d;
         4'h3220 	:	val_out <= 4'hf8a6;
         4'h3221 	:	val_out <= 4'hf8a6;
         4'h3222 	:	val_out <= 4'hf8a6;
         4'h3223 	:	val_out <= 4'hf8a6;
         4'h3228 	:	val_out <= 4'hf8ae;
         4'h3229 	:	val_out <= 4'hf8ae;
         4'h322a 	:	val_out <= 4'hf8ae;
         4'h322b 	:	val_out <= 4'hf8ae;
         4'h3230 	:	val_out <= 4'hf8b6;
         4'h3231 	:	val_out <= 4'hf8b6;
         4'h3232 	:	val_out <= 4'hf8b6;
         4'h3233 	:	val_out <= 4'hf8b6;
         4'h3238 	:	val_out <= 4'hf8bf;
         4'h3239 	:	val_out <= 4'hf8bf;
         4'h323a 	:	val_out <= 4'hf8bf;
         4'h323b 	:	val_out <= 4'hf8bf;
         4'h3240 	:	val_out <= 4'hf8c7;
         4'h3241 	:	val_out <= 4'hf8c7;
         4'h3242 	:	val_out <= 4'hf8c7;
         4'h3243 	:	val_out <= 4'hf8c7;
         4'h3248 	:	val_out <= 4'hf8cf;
         4'h3249 	:	val_out <= 4'hf8cf;
         4'h324a 	:	val_out <= 4'hf8cf;
         4'h324b 	:	val_out <= 4'hf8cf;
         4'h3250 	:	val_out <= 4'hf8d8;
         4'h3251 	:	val_out <= 4'hf8d8;
         4'h3252 	:	val_out <= 4'hf8d8;
         4'h3253 	:	val_out <= 4'hf8d8;
         4'h3258 	:	val_out <= 4'hf8e0;
         4'h3259 	:	val_out <= 4'hf8e0;
         4'h325a 	:	val_out <= 4'hf8e0;
         4'h325b 	:	val_out <= 4'hf8e0;
         4'h3260 	:	val_out <= 4'hf8e8;
         4'h3261 	:	val_out <= 4'hf8e8;
         4'h3262 	:	val_out <= 4'hf8e8;
         4'h3263 	:	val_out <= 4'hf8e8;
         4'h3268 	:	val_out <= 4'hf8f1;
         4'h3269 	:	val_out <= 4'hf8f1;
         4'h326a 	:	val_out <= 4'hf8f1;
         4'h326b 	:	val_out <= 4'hf8f1;
         4'h3270 	:	val_out <= 4'hf8f9;
         4'h3271 	:	val_out <= 4'hf8f9;
         4'h3272 	:	val_out <= 4'hf8f9;
         4'h3273 	:	val_out <= 4'hf8f9;
         4'h3278 	:	val_out <= 4'hf901;
         4'h3279 	:	val_out <= 4'hf901;
         4'h327a 	:	val_out <= 4'hf901;
         4'h327b 	:	val_out <= 4'hf901;
         4'h3280 	:	val_out <= 4'hf909;
         4'h3281 	:	val_out <= 4'hf909;
         4'h3282 	:	val_out <= 4'hf909;
         4'h3283 	:	val_out <= 4'hf909;
         4'h3288 	:	val_out <= 4'hf911;
         4'h3289 	:	val_out <= 4'hf911;
         4'h328a 	:	val_out <= 4'hf911;
         4'h328b 	:	val_out <= 4'hf911;
         4'h3290 	:	val_out <= 4'hf919;
         4'h3291 	:	val_out <= 4'hf919;
         4'h3292 	:	val_out <= 4'hf919;
         4'h3293 	:	val_out <= 4'hf919;
         4'h3298 	:	val_out <= 4'hf922;
         4'h3299 	:	val_out <= 4'hf922;
         4'h329a 	:	val_out <= 4'hf922;
         4'h329b 	:	val_out <= 4'hf922;
         4'h32a0 	:	val_out <= 4'hf92a;
         4'h32a1 	:	val_out <= 4'hf92a;
         4'h32a2 	:	val_out <= 4'hf92a;
         4'h32a3 	:	val_out <= 4'hf92a;
         4'h32a8 	:	val_out <= 4'hf932;
         4'h32a9 	:	val_out <= 4'hf932;
         4'h32aa 	:	val_out <= 4'hf932;
         4'h32ab 	:	val_out <= 4'hf932;
         4'h32b0 	:	val_out <= 4'hf93a;
         4'h32b1 	:	val_out <= 4'hf93a;
         4'h32b2 	:	val_out <= 4'hf93a;
         4'h32b3 	:	val_out <= 4'hf93a;
         4'h32b8 	:	val_out <= 4'hf942;
         4'h32b9 	:	val_out <= 4'hf942;
         4'h32ba 	:	val_out <= 4'hf942;
         4'h32bb 	:	val_out <= 4'hf942;
         4'h32c0 	:	val_out <= 4'hf94a;
         4'h32c1 	:	val_out <= 4'hf94a;
         4'h32c2 	:	val_out <= 4'hf94a;
         4'h32c3 	:	val_out <= 4'hf94a;
         4'h32c8 	:	val_out <= 4'hf952;
         4'h32c9 	:	val_out <= 4'hf952;
         4'h32ca 	:	val_out <= 4'hf952;
         4'h32cb 	:	val_out <= 4'hf952;
         4'h32d0 	:	val_out <= 4'hf95a;
         4'h32d1 	:	val_out <= 4'hf95a;
         4'h32d2 	:	val_out <= 4'hf95a;
         4'h32d3 	:	val_out <= 4'hf95a;
         4'h32d8 	:	val_out <= 4'hf962;
         4'h32d9 	:	val_out <= 4'hf962;
         4'h32da 	:	val_out <= 4'hf962;
         4'h32db 	:	val_out <= 4'hf962;
         4'h32e0 	:	val_out <= 4'hf96a;
         4'h32e1 	:	val_out <= 4'hf96a;
         4'h32e2 	:	val_out <= 4'hf96a;
         4'h32e3 	:	val_out <= 4'hf96a;
         4'h32e8 	:	val_out <= 4'hf972;
         4'h32e9 	:	val_out <= 4'hf972;
         4'h32ea 	:	val_out <= 4'hf972;
         4'h32eb 	:	val_out <= 4'hf972;
         4'h32f0 	:	val_out <= 4'hf97a;
         4'h32f1 	:	val_out <= 4'hf97a;
         4'h32f2 	:	val_out <= 4'hf97a;
         4'h32f3 	:	val_out <= 4'hf97a;
         4'h32f8 	:	val_out <= 4'hf982;
         4'h32f9 	:	val_out <= 4'hf982;
         4'h32fa 	:	val_out <= 4'hf982;
         4'h32fb 	:	val_out <= 4'hf982;
         4'h3300 	:	val_out <= 4'hf98a;
         4'h3301 	:	val_out <= 4'hf98a;
         4'h3302 	:	val_out <= 4'hf98a;
         4'h3303 	:	val_out <= 4'hf98a;
         4'h3308 	:	val_out <= 4'hf992;
         4'h3309 	:	val_out <= 4'hf992;
         4'h330a 	:	val_out <= 4'hf992;
         4'h330b 	:	val_out <= 4'hf992;
         4'h3310 	:	val_out <= 4'hf999;
         4'h3311 	:	val_out <= 4'hf999;
         4'h3312 	:	val_out <= 4'hf999;
         4'h3313 	:	val_out <= 4'hf999;
         4'h3318 	:	val_out <= 4'hf9a1;
         4'h3319 	:	val_out <= 4'hf9a1;
         4'h331a 	:	val_out <= 4'hf9a1;
         4'h331b 	:	val_out <= 4'hf9a1;
         4'h3320 	:	val_out <= 4'hf9a9;
         4'h3321 	:	val_out <= 4'hf9a9;
         4'h3322 	:	val_out <= 4'hf9a9;
         4'h3323 	:	val_out <= 4'hf9a9;
         4'h3328 	:	val_out <= 4'hf9b1;
         4'h3329 	:	val_out <= 4'hf9b1;
         4'h332a 	:	val_out <= 4'hf9b1;
         4'h332b 	:	val_out <= 4'hf9b1;
         4'h3330 	:	val_out <= 4'hf9b9;
         4'h3331 	:	val_out <= 4'hf9b9;
         4'h3332 	:	val_out <= 4'hf9b9;
         4'h3333 	:	val_out <= 4'hf9b9;
         4'h3338 	:	val_out <= 4'hf9c0;
         4'h3339 	:	val_out <= 4'hf9c0;
         4'h333a 	:	val_out <= 4'hf9c0;
         4'h333b 	:	val_out <= 4'hf9c0;
         4'h3340 	:	val_out <= 4'hf9c8;
         4'h3341 	:	val_out <= 4'hf9c8;
         4'h3342 	:	val_out <= 4'hf9c8;
         4'h3343 	:	val_out <= 4'hf9c8;
         4'h3348 	:	val_out <= 4'hf9d0;
         4'h3349 	:	val_out <= 4'hf9d0;
         4'h334a 	:	val_out <= 4'hf9d0;
         4'h334b 	:	val_out <= 4'hf9d0;
         4'h3350 	:	val_out <= 4'hf9d8;
         4'h3351 	:	val_out <= 4'hf9d8;
         4'h3352 	:	val_out <= 4'hf9d8;
         4'h3353 	:	val_out <= 4'hf9d8;
         4'h3358 	:	val_out <= 4'hf9df;
         4'h3359 	:	val_out <= 4'hf9df;
         4'h335a 	:	val_out <= 4'hf9df;
         4'h335b 	:	val_out <= 4'hf9df;
         4'h3360 	:	val_out <= 4'hf9e7;
         4'h3361 	:	val_out <= 4'hf9e7;
         4'h3362 	:	val_out <= 4'hf9e7;
         4'h3363 	:	val_out <= 4'hf9e7;
         4'h3368 	:	val_out <= 4'hf9ef;
         4'h3369 	:	val_out <= 4'hf9ef;
         4'h336a 	:	val_out <= 4'hf9ef;
         4'h336b 	:	val_out <= 4'hf9ef;
         4'h3370 	:	val_out <= 4'hf9f6;
         4'h3371 	:	val_out <= 4'hf9f6;
         4'h3372 	:	val_out <= 4'hf9f6;
         4'h3373 	:	val_out <= 4'hf9f6;
         4'h3378 	:	val_out <= 4'hf9fe;
         4'h3379 	:	val_out <= 4'hf9fe;
         4'h337a 	:	val_out <= 4'hf9fe;
         4'h337b 	:	val_out <= 4'hf9fe;
         4'h3380 	:	val_out <= 4'hfa05;
         4'h3381 	:	val_out <= 4'hfa05;
         4'h3382 	:	val_out <= 4'hfa05;
         4'h3383 	:	val_out <= 4'hfa05;
         4'h3388 	:	val_out <= 4'hfa0d;
         4'h3389 	:	val_out <= 4'hfa0d;
         4'h338a 	:	val_out <= 4'hfa0d;
         4'h338b 	:	val_out <= 4'hfa0d;
         4'h3390 	:	val_out <= 4'hfa15;
         4'h3391 	:	val_out <= 4'hfa15;
         4'h3392 	:	val_out <= 4'hfa15;
         4'h3393 	:	val_out <= 4'hfa15;
         4'h3398 	:	val_out <= 4'hfa1c;
         4'h3399 	:	val_out <= 4'hfa1c;
         4'h339a 	:	val_out <= 4'hfa1c;
         4'h339b 	:	val_out <= 4'hfa1c;
         4'h33a0 	:	val_out <= 4'hfa24;
         4'h33a1 	:	val_out <= 4'hfa24;
         4'h33a2 	:	val_out <= 4'hfa24;
         4'h33a3 	:	val_out <= 4'hfa24;
         4'h33a8 	:	val_out <= 4'hfa2b;
         4'h33a9 	:	val_out <= 4'hfa2b;
         4'h33aa 	:	val_out <= 4'hfa2b;
         4'h33ab 	:	val_out <= 4'hfa2b;
         4'h33b0 	:	val_out <= 4'hfa33;
         4'h33b1 	:	val_out <= 4'hfa33;
         4'h33b2 	:	val_out <= 4'hfa33;
         4'h33b3 	:	val_out <= 4'hfa33;
         4'h33b8 	:	val_out <= 4'hfa3a;
         4'h33b9 	:	val_out <= 4'hfa3a;
         4'h33ba 	:	val_out <= 4'hfa3a;
         4'h33bb 	:	val_out <= 4'hfa3a;
         4'h33c0 	:	val_out <= 4'hfa42;
         4'h33c1 	:	val_out <= 4'hfa42;
         4'h33c2 	:	val_out <= 4'hfa42;
         4'h33c3 	:	val_out <= 4'hfa42;
         4'h33c8 	:	val_out <= 4'hfa49;
         4'h33c9 	:	val_out <= 4'hfa49;
         4'h33ca 	:	val_out <= 4'hfa49;
         4'h33cb 	:	val_out <= 4'hfa49;
         4'h33d0 	:	val_out <= 4'hfa50;
         4'h33d1 	:	val_out <= 4'hfa50;
         4'h33d2 	:	val_out <= 4'hfa50;
         4'h33d3 	:	val_out <= 4'hfa50;
         4'h33d8 	:	val_out <= 4'hfa58;
         4'h33d9 	:	val_out <= 4'hfa58;
         4'h33da 	:	val_out <= 4'hfa58;
         4'h33db 	:	val_out <= 4'hfa58;
         4'h33e0 	:	val_out <= 4'hfa5f;
         4'h33e1 	:	val_out <= 4'hfa5f;
         4'h33e2 	:	val_out <= 4'hfa5f;
         4'h33e3 	:	val_out <= 4'hfa5f;
         4'h33e8 	:	val_out <= 4'hfa67;
         4'h33e9 	:	val_out <= 4'hfa67;
         4'h33ea 	:	val_out <= 4'hfa67;
         4'h33eb 	:	val_out <= 4'hfa67;
         4'h33f0 	:	val_out <= 4'hfa6e;
         4'h33f1 	:	val_out <= 4'hfa6e;
         4'h33f2 	:	val_out <= 4'hfa6e;
         4'h33f3 	:	val_out <= 4'hfa6e;
         4'h33f8 	:	val_out <= 4'hfa75;
         4'h33f9 	:	val_out <= 4'hfa75;
         4'h33fa 	:	val_out <= 4'hfa75;
         4'h33fb 	:	val_out <= 4'hfa75;
         4'h3400 	:	val_out <= 4'hfa7d;
         4'h3401 	:	val_out <= 4'hfa7d;
         4'h3402 	:	val_out <= 4'hfa7d;
         4'h3403 	:	val_out <= 4'hfa7d;
         4'h3408 	:	val_out <= 4'hfa84;
         4'h3409 	:	val_out <= 4'hfa84;
         4'h340a 	:	val_out <= 4'hfa84;
         4'h340b 	:	val_out <= 4'hfa84;
         4'h3410 	:	val_out <= 4'hfa8b;
         4'h3411 	:	val_out <= 4'hfa8b;
         4'h3412 	:	val_out <= 4'hfa8b;
         4'h3413 	:	val_out <= 4'hfa8b;
         4'h3418 	:	val_out <= 4'hfa92;
         4'h3419 	:	val_out <= 4'hfa92;
         4'h341a 	:	val_out <= 4'hfa92;
         4'h341b 	:	val_out <= 4'hfa92;
         4'h3420 	:	val_out <= 4'hfa9a;
         4'h3421 	:	val_out <= 4'hfa9a;
         4'h3422 	:	val_out <= 4'hfa9a;
         4'h3423 	:	val_out <= 4'hfa9a;
         4'h3428 	:	val_out <= 4'hfaa1;
         4'h3429 	:	val_out <= 4'hfaa1;
         4'h342a 	:	val_out <= 4'hfaa1;
         4'h342b 	:	val_out <= 4'hfaa1;
         4'h3430 	:	val_out <= 4'hfaa8;
         4'h3431 	:	val_out <= 4'hfaa8;
         4'h3432 	:	val_out <= 4'hfaa8;
         4'h3433 	:	val_out <= 4'hfaa8;
         4'h3438 	:	val_out <= 4'hfaaf;
         4'h3439 	:	val_out <= 4'hfaaf;
         4'h343a 	:	val_out <= 4'hfaaf;
         4'h343b 	:	val_out <= 4'hfaaf;
         4'h3440 	:	val_out <= 4'hfab6;
         4'h3441 	:	val_out <= 4'hfab6;
         4'h3442 	:	val_out <= 4'hfab6;
         4'h3443 	:	val_out <= 4'hfab6;
         4'h3448 	:	val_out <= 4'hfabd;
         4'h3449 	:	val_out <= 4'hfabd;
         4'h344a 	:	val_out <= 4'hfabd;
         4'h344b 	:	val_out <= 4'hfabd;
         4'h3450 	:	val_out <= 4'hfac5;
         4'h3451 	:	val_out <= 4'hfac5;
         4'h3452 	:	val_out <= 4'hfac5;
         4'h3453 	:	val_out <= 4'hfac5;
         4'h3458 	:	val_out <= 4'hfacc;
         4'h3459 	:	val_out <= 4'hfacc;
         4'h345a 	:	val_out <= 4'hfacc;
         4'h345b 	:	val_out <= 4'hfacc;
         4'h3460 	:	val_out <= 4'hfad3;
         4'h3461 	:	val_out <= 4'hfad3;
         4'h3462 	:	val_out <= 4'hfad3;
         4'h3463 	:	val_out <= 4'hfad3;
         4'h3468 	:	val_out <= 4'hfada;
         4'h3469 	:	val_out <= 4'hfada;
         4'h346a 	:	val_out <= 4'hfada;
         4'h346b 	:	val_out <= 4'hfada;
         4'h3470 	:	val_out <= 4'hfae1;
         4'h3471 	:	val_out <= 4'hfae1;
         4'h3472 	:	val_out <= 4'hfae1;
         4'h3473 	:	val_out <= 4'hfae1;
         4'h3478 	:	val_out <= 4'hfae8;
         4'h3479 	:	val_out <= 4'hfae8;
         4'h347a 	:	val_out <= 4'hfae8;
         4'h347b 	:	val_out <= 4'hfae8;
         4'h3480 	:	val_out <= 4'hfaef;
         4'h3481 	:	val_out <= 4'hfaef;
         4'h3482 	:	val_out <= 4'hfaef;
         4'h3483 	:	val_out <= 4'hfaef;
         4'h3488 	:	val_out <= 4'hfaf6;
         4'h3489 	:	val_out <= 4'hfaf6;
         4'h348a 	:	val_out <= 4'hfaf6;
         4'h348b 	:	val_out <= 4'hfaf6;
         4'h3490 	:	val_out <= 4'hfafd;
         4'h3491 	:	val_out <= 4'hfafd;
         4'h3492 	:	val_out <= 4'hfafd;
         4'h3493 	:	val_out <= 4'hfafd;
         4'h3498 	:	val_out <= 4'hfb04;
         4'h3499 	:	val_out <= 4'hfb04;
         4'h349a 	:	val_out <= 4'hfb04;
         4'h349b 	:	val_out <= 4'hfb04;
         4'h34a0 	:	val_out <= 4'hfb0b;
         4'h34a1 	:	val_out <= 4'hfb0b;
         4'h34a2 	:	val_out <= 4'hfb0b;
         4'h34a3 	:	val_out <= 4'hfb0b;
         4'h34a8 	:	val_out <= 4'hfb12;
         4'h34a9 	:	val_out <= 4'hfb12;
         4'h34aa 	:	val_out <= 4'hfb12;
         4'h34ab 	:	val_out <= 4'hfb12;
         4'h34b0 	:	val_out <= 4'hfb19;
         4'h34b1 	:	val_out <= 4'hfb19;
         4'h34b2 	:	val_out <= 4'hfb19;
         4'h34b3 	:	val_out <= 4'hfb19;
         4'h34b8 	:	val_out <= 4'hfb1f;
         4'h34b9 	:	val_out <= 4'hfb1f;
         4'h34ba 	:	val_out <= 4'hfb1f;
         4'h34bb 	:	val_out <= 4'hfb1f;
         4'h34c0 	:	val_out <= 4'hfb26;
         4'h34c1 	:	val_out <= 4'hfb26;
         4'h34c2 	:	val_out <= 4'hfb26;
         4'h34c3 	:	val_out <= 4'hfb26;
         4'h34c8 	:	val_out <= 4'hfb2d;
         4'h34c9 	:	val_out <= 4'hfb2d;
         4'h34ca 	:	val_out <= 4'hfb2d;
         4'h34cb 	:	val_out <= 4'hfb2d;
         4'h34d0 	:	val_out <= 4'hfb34;
         4'h34d1 	:	val_out <= 4'hfb34;
         4'h34d2 	:	val_out <= 4'hfb34;
         4'h34d3 	:	val_out <= 4'hfb34;
         4'h34d8 	:	val_out <= 4'hfb3b;
         4'h34d9 	:	val_out <= 4'hfb3b;
         4'h34da 	:	val_out <= 4'hfb3b;
         4'h34db 	:	val_out <= 4'hfb3b;
         4'h34e0 	:	val_out <= 4'hfb42;
         4'h34e1 	:	val_out <= 4'hfb42;
         4'h34e2 	:	val_out <= 4'hfb42;
         4'h34e3 	:	val_out <= 4'hfb42;
         4'h34e8 	:	val_out <= 4'hfb48;
         4'h34e9 	:	val_out <= 4'hfb48;
         4'h34ea 	:	val_out <= 4'hfb48;
         4'h34eb 	:	val_out <= 4'hfb48;
         4'h34f0 	:	val_out <= 4'hfb4f;
         4'h34f1 	:	val_out <= 4'hfb4f;
         4'h34f2 	:	val_out <= 4'hfb4f;
         4'h34f3 	:	val_out <= 4'hfb4f;
         4'h34f8 	:	val_out <= 4'hfb56;
         4'h34f9 	:	val_out <= 4'hfb56;
         4'h34fa 	:	val_out <= 4'hfb56;
         4'h34fb 	:	val_out <= 4'hfb56;
         4'h3500 	:	val_out <= 4'hfb5d;
         4'h3501 	:	val_out <= 4'hfb5d;
         4'h3502 	:	val_out <= 4'hfb5d;
         4'h3503 	:	val_out <= 4'hfb5d;
         4'h3508 	:	val_out <= 4'hfb63;
         4'h3509 	:	val_out <= 4'hfb63;
         4'h350a 	:	val_out <= 4'hfb63;
         4'h350b 	:	val_out <= 4'hfb63;
         4'h3510 	:	val_out <= 4'hfb6a;
         4'h3511 	:	val_out <= 4'hfb6a;
         4'h3512 	:	val_out <= 4'hfb6a;
         4'h3513 	:	val_out <= 4'hfb6a;
         4'h3518 	:	val_out <= 4'hfb71;
         4'h3519 	:	val_out <= 4'hfb71;
         4'h351a 	:	val_out <= 4'hfb71;
         4'h351b 	:	val_out <= 4'hfb71;
         4'h3520 	:	val_out <= 4'hfb77;
         4'h3521 	:	val_out <= 4'hfb77;
         4'h3522 	:	val_out <= 4'hfb77;
         4'h3523 	:	val_out <= 4'hfb77;
         4'h3528 	:	val_out <= 4'hfb7e;
         4'h3529 	:	val_out <= 4'hfb7e;
         4'h352a 	:	val_out <= 4'hfb7e;
         4'h352b 	:	val_out <= 4'hfb7e;
         4'h3530 	:	val_out <= 4'hfb84;
         4'h3531 	:	val_out <= 4'hfb84;
         4'h3532 	:	val_out <= 4'hfb84;
         4'h3533 	:	val_out <= 4'hfb84;
         4'h3538 	:	val_out <= 4'hfb8b;
         4'h3539 	:	val_out <= 4'hfb8b;
         4'h353a 	:	val_out <= 4'hfb8b;
         4'h353b 	:	val_out <= 4'hfb8b;
         4'h3540 	:	val_out <= 4'hfb92;
         4'h3541 	:	val_out <= 4'hfb92;
         4'h3542 	:	val_out <= 4'hfb92;
         4'h3543 	:	val_out <= 4'hfb92;
         4'h3548 	:	val_out <= 4'hfb98;
         4'h3549 	:	val_out <= 4'hfb98;
         4'h354a 	:	val_out <= 4'hfb98;
         4'h354b 	:	val_out <= 4'hfb98;
         4'h3550 	:	val_out <= 4'hfb9f;
         4'h3551 	:	val_out <= 4'hfb9f;
         4'h3552 	:	val_out <= 4'hfb9f;
         4'h3553 	:	val_out <= 4'hfb9f;
         4'h3558 	:	val_out <= 4'hfba5;
         4'h3559 	:	val_out <= 4'hfba5;
         4'h355a 	:	val_out <= 4'hfba5;
         4'h355b 	:	val_out <= 4'hfba5;
         4'h3560 	:	val_out <= 4'hfbac;
         4'h3561 	:	val_out <= 4'hfbac;
         4'h3562 	:	val_out <= 4'hfbac;
         4'h3563 	:	val_out <= 4'hfbac;
         4'h3568 	:	val_out <= 4'hfbb2;
         4'h3569 	:	val_out <= 4'hfbb2;
         4'h356a 	:	val_out <= 4'hfbb2;
         4'h356b 	:	val_out <= 4'hfbb2;
         4'h3570 	:	val_out <= 4'hfbb9;
         4'h3571 	:	val_out <= 4'hfbb9;
         4'h3572 	:	val_out <= 4'hfbb9;
         4'h3573 	:	val_out <= 4'hfbb9;
         4'h3578 	:	val_out <= 4'hfbbf;
         4'h3579 	:	val_out <= 4'hfbbf;
         4'h357a 	:	val_out <= 4'hfbbf;
         4'h357b 	:	val_out <= 4'hfbbf;
         4'h3580 	:	val_out <= 4'hfbc5;
         4'h3581 	:	val_out <= 4'hfbc5;
         4'h3582 	:	val_out <= 4'hfbc5;
         4'h3583 	:	val_out <= 4'hfbc5;
         4'h3588 	:	val_out <= 4'hfbcc;
         4'h3589 	:	val_out <= 4'hfbcc;
         4'h358a 	:	val_out <= 4'hfbcc;
         4'h358b 	:	val_out <= 4'hfbcc;
         4'h3590 	:	val_out <= 4'hfbd2;
         4'h3591 	:	val_out <= 4'hfbd2;
         4'h3592 	:	val_out <= 4'hfbd2;
         4'h3593 	:	val_out <= 4'hfbd2;
         4'h3598 	:	val_out <= 4'hfbd9;
         4'h3599 	:	val_out <= 4'hfbd9;
         4'h359a 	:	val_out <= 4'hfbd9;
         4'h359b 	:	val_out <= 4'hfbd9;
         4'h35a0 	:	val_out <= 4'hfbdf;
         4'h35a1 	:	val_out <= 4'hfbdf;
         4'h35a2 	:	val_out <= 4'hfbdf;
         4'h35a3 	:	val_out <= 4'hfbdf;
         4'h35a8 	:	val_out <= 4'hfbe5;
         4'h35a9 	:	val_out <= 4'hfbe5;
         4'h35aa 	:	val_out <= 4'hfbe5;
         4'h35ab 	:	val_out <= 4'hfbe5;
         4'h35b0 	:	val_out <= 4'hfbeb;
         4'h35b1 	:	val_out <= 4'hfbeb;
         4'h35b2 	:	val_out <= 4'hfbeb;
         4'h35b3 	:	val_out <= 4'hfbeb;
         4'h35b8 	:	val_out <= 4'hfbf2;
         4'h35b9 	:	val_out <= 4'hfbf2;
         4'h35ba 	:	val_out <= 4'hfbf2;
         4'h35bb 	:	val_out <= 4'hfbf2;
         4'h35c0 	:	val_out <= 4'hfbf8;
         4'h35c1 	:	val_out <= 4'hfbf8;
         4'h35c2 	:	val_out <= 4'hfbf8;
         4'h35c3 	:	val_out <= 4'hfbf8;
         4'h35c8 	:	val_out <= 4'hfbfe;
         4'h35c9 	:	val_out <= 4'hfbfe;
         4'h35ca 	:	val_out <= 4'hfbfe;
         4'h35cb 	:	val_out <= 4'hfbfe;
         4'h35d0 	:	val_out <= 4'hfc05;
         4'h35d1 	:	val_out <= 4'hfc05;
         4'h35d2 	:	val_out <= 4'hfc05;
         4'h35d3 	:	val_out <= 4'hfc05;
         4'h35d8 	:	val_out <= 4'hfc0b;
         4'h35d9 	:	val_out <= 4'hfc0b;
         4'h35da 	:	val_out <= 4'hfc0b;
         4'h35db 	:	val_out <= 4'hfc0b;
         4'h35e0 	:	val_out <= 4'hfc11;
         4'h35e1 	:	val_out <= 4'hfc11;
         4'h35e2 	:	val_out <= 4'hfc11;
         4'h35e3 	:	val_out <= 4'hfc11;
         4'h35e8 	:	val_out <= 4'hfc17;
         4'h35e9 	:	val_out <= 4'hfc17;
         4'h35ea 	:	val_out <= 4'hfc17;
         4'h35eb 	:	val_out <= 4'hfc17;
         4'h35f0 	:	val_out <= 4'hfc1d;
         4'h35f1 	:	val_out <= 4'hfc1d;
         4'h35f2 	:	val_out <= 4'hfc1d;
         4'h35f3 	:	val_out <= 4'hfc1d;
         4'h35f8 	:	val_out <= 4'hfc23;
         4'h35f9 	:	val_out <= 4'hfc23;
         4'h35fa 	:	val_out <= 4'hfc23;
         4'h35fb 	:	val_out <= 4'hfc23;
         4'h3600 	:	val_out <= 4'hfc29;
         4'h3601 	:	val_out <= 4'hfc29;
         4'h3602 	:	val_out <= 4'hfc29;
         4'h3603 	:	val_out <= 4'hfc29;
         4'h3608 	:	val_out <= 4'hfc30;
         4'h3609 	:	val_out <= 4'hfc30;
         4'h360a 	:	val_out <= 4'hfc30;
         4'h360b 	:	val_out <= 4'hfc30;
         4'h3610 	:	val_out <= 4'hfc36;
         4'h3611 	:	val_out <= 4'hfc36;
         4'h3612 	:	val_out <= 4'hfc36;
         4'h3613 	:	val_out <= 4'hfc36;
         4'h3618 	:	val_out <= 4'hfc3c;
         4'h3619 	:	val_out <= 4'hfc3c;
         4'h361a 	:	val_out <= 4'hfc3c;
         4'h361b 	:	val_out <= 4'hfc3c;
         4'h3620 	:	val_out <= 4'hfc42;
         4'h3621 	:	val_out <= 4'hfc42;
         4'h3622 	:	val_out <= 4'hfc42;
         4'h3623 	:	val_out <= 4'hfc42;
         4'h3628 	:	val_out <= 4'hfc48;
         4'h3629 	:	val_out <= 4'hfc48;
         4'h362a 	:	val_out <= 4'hfc48;
         4'h362b 	:	val_out <= 4'hfc48;
         4'h3630 	:	val_out <= 4'hfc4e;
         4'h3631 	:	val_out <= 4'hfc4e;
         4'h3632 	:	val_out <= 4'hfc4e;
         4'h3633 	:	val_out <= 4'hfc4e;
         4'h3638 	:	val_out <= 4'hfc54;
         4'h3639 	:	val_out <= 4'hfc54;
         4'h363a 	:	val_out <= 4'hfc54;
         4'h363b 	:	val_out <= 4'hfc54;
         4'h3640 	:	val_out <= 4'hfc5a;
         4'h3641 	:	val_out <= 4'hfc5a;
         4'h3642 	:	val_out <= 4'hfc5a;
         4'h3643 	:	val_out <= 4'hfc5a;
         4'h3648 	:	val_out <= 4'hfc60;
         4'h3649 	:	val_out <= 4'hfc60;
         4'h364a 	:	val_out <= 4'hfc60;
         4'h364b 	:	val_out <= 4'hfc60;
         4'h3650 	:	val_out <= 4'hfc66;
         4'h3651 	:	val_out <= 4'hfc66;
         4'h3652 	:	val_out <= 4'hfc66;
         4'h3653 	:	val_out <= 4'hfc66;
         4'h3658 	:	val_out <= 4'hfc6c;
         4'h3659 	:	val_out <= 4'hfc6c;
         4'h365a 	:	val_out <= 4'hfc6c;
         4'h365b 	:	val_out <= 4'hfc6c;
         4'h3660 	:	val_out <= 4'hfc71;
         4'h3661 	:	val_out <= 4'hfc71;
         4'h3662 	:	val_out <= 4'hfc71;
         4'h3663 	:	val_out <= 4'hfc71;
         4'h3668 	:	val_out <= 4'hfc77;
         4'h3669 	:	val_out <= 4'hfc77;
         4'h366a 	:	val_out <= 4'hfc77;
         4'h366b 	:	val_out <= 4'hfc77;
         4'h3670 	:	val_out <= 4'hfc7d;
         4'h3671 	:	val_out <= 4'hfc7d;
         4'h3672 	:	val_out <= 4'hfc7d;
         4'h3673 	:	val_out <= 4'hfc7d;
         4'h3678 	:	val_out <= 4'hfc83;
         4'h3679 	:	val_out <= 4'hfc83;
         4'h367a 	:	val_out <= 4'hfc83;
         4'h367b 	:	val_out <= 4'hfc83;
         4'h3680 	:	val_out <= 4'hfc89;
         4'h3681 	:	val_out <= 4'hfc89;
         4'h3682 	:	val_out <= 4'hfc89;
         4'h3683 	:	val_out <= 4'hfc89;
         4'h3688 	:	val_out <= 4'hfc8f;
         4'h3689 	:	val_out <= 4'hfc8f;
         4'h368a 	:	val_out <= 4'hfc8f;
         4'h368b 	:	val_out <= 4'hfc8f;
         4'h3690 	:	val_out <= 4'hfc94;
         4'h3691 	:	val_out <= 4'hfc94;
         4'h3692 	:	val_out <= 4'hfc94;
         4'h3693 	:	val_out <= 4'hfc94;
         4'h3698 	:	val_out <= 4'hfc9a;
         4'h3699 	:	val_out <= 4'hfc9a;
         4'h369a 	:	val_out <= 4'hfc9a;
         4'h369b 	:	val_out <= 4'hfc9a;
         4'h36a0 	:	val_out <= 4'hfca0;
         4'h36a1 	:	val_out <= 4'hfca0;
         4'h36a2 	:	val_out <= 4'hfca0;
         4'h36a3 	:	val_out <= 4'hfca0;
         4'h36a8 	:	val_out <= 4'hfca6;
         4'h36a9 	:	val_out <= 4'hfca6;
         4'h36aa 	:	val_out <= 4'hfca6;
         4'h36ab 	:	val_out <= 4'hfca6;
         4'h36b0 	:	val_out <= 4'hfcab;
         4'h36b1 	:	val_out <= 4'hfcab;
         4'h36b2 	:	val_out <= 4'hfcab;
         4'h36b3 	:	val_out <= 4'hfcab;
         4'h36b8 	:	val_out <= 4'hfcb1;
         4'h36b9 	:	val_out <= 4'hfcb1;
         4'h36ba 	:	val_out <= 4'hfcb1;
         4'h36bb 	:	val_out <= 4'hfcb1;
         4'h36c0 	:	val_out <= 4'hfcb7;
         4'h36c1 	:	val_out <= 4'hfcb7;
         4'h36c2 	:	val_out <= 4'hfcb7;
         4'h36c3 	:	val_out <= 4'hfcb7;
         4'h36c8 	:	val_out <= 4'hfcbc;
         4'h36c9 	:	val_out <= 4'hfcbc;
         4'h36ca 	:	val_out <= 4'hfcbc;
         4'h36cb 	:	val_out <= 4'hfcbc;
         4'h36d0 	:	val_out <= 4'hfcc2;
         4'h36d1 	:	val_out <= 4'hfcc2;
         4'h36d2 	:	val_out <= 4'hfcc2;
         4'h36d3 	:	val_out <= 4'hfcc2;
         4'h36d8 	:	val_out <= 4'hfcc8;
         4'h36d9 	:	val_out <= 4'hfcc8;
         4'h36da 	:	val_out <= 4'hfcc8;
         4'h36db 	:	val_out <= 4'hfcc8;
         4'h36e0 	:	val_out <= 4'hfccd;
         4'h36e1 	:	val_out <= 4'hfccd;
         4'h36e2 	:	val_out <= 4'hfccd;
         4'h36e3 	:	val_out <= 4'hfccd;
         4'h36e8 	:	val_out <= 4'hfcd3;
         4'h36e9 	:	val_out <= 4'hfcd3;
         4'h36ea 	:	val_out <= 4'hfcd3;
         4'h36eb 	:	val_out <= 4'hfcd3;
         4'h36f0 	:	val_out <= 4'hfcd8;
         4'h36f1 	:	val_out <= 4'hfcd8;
         4'h36f2 	:	val_out <= 4'hfcd8;
         4'h36f3 	:	val_out <= 4'hfcd8;
         4'h36f8 	:	val_out <= 4'hfcde;
         4'h36f9 	:	val_out <= 4'hfcde;
         4'h36fa 	:	val_out <= 4'hfcde;
         4'h36fb 	:	val_out <= 4'hfcde;
         4'h3700 	:	val_out <= 4'hfce3;
         4'h3701 	:	val_out <= 4'hfce3;
         4'h3702 	:	val_out <= 4'hfce3;
         4'h3703 	:	val_out <= 4'hfce3;
         4'h3708 	:	val_out <= 4'hfce9;
         4'h3709 	:	val_out <= 4'hfce9;
         4'h370a 	:	val_out <= 4'hfce9;
         4'h370b 	:	val_out <= 4'hfce9;
         4'h3710 	:	val_out <= 4'hfcee;
         4'h3711 	:	val_out <= 4'hfcee;
         4'h3712 	:	val_out <= 4'hfcee;
         4'h3713 	:	val_out <= 4'hfcee;
         4'h3718 	:	val_out <= 4'hfcf4;
         4'h3719 	:	val_out <= 4'hfcf4;
         4'h371a 	:	val_out <= 4'hfcf4;
         4'h371b 	:	val_out <= 4'hfcf4;
         4'h3720 	:	val_out <= 4'hfcf9;
         4'h3721 	:	val_out <= 4'hfcf9;
         4'h3722 	:	val_out <= 4'hfcf9;
         4'h3723 	:	val_out <= 4'hfcf9;
         4'h3728 	:	val_out <= 4'hfcff;
         4'h3729 	:	val_out <= 4'hfcff;
         4'h372a 	:	val_out <= 4'hfcff;
         4'h372b 	:	val_out <= 4'hfcff;
         4'h3730 	:	val_out <= 4'hfd04;
         4'h3731 	:	val_out <= 4'hfd04;
         4'h3732 	:	val_out <= 4'hfd04;
         4'h3733 	:	val_out <= 4'hfd04;
         4'h3738 	:	val_out <= 4'hfd09;
         4'h3739 	:	val_out <= 4'hfd09;
         4'h373a 	:	val_out <= 4'hfd09;
         4'h373b 	:	val_out <= 4'hfd09;
         4'h3740 	:	val_out <= 4'hfd0f;
         4'h3741 	:	val_out <= 4'hfd0f;
         4'h3742 	:	val_out <= 4'hfd0f;
         4'h3743 	:	val_out <= 4'hfd0f;
         4'h3748 	:	val_out <= 4'hfd14;
         4'h3749 	:	val_out <= 4'hfd14;
         4'h374a 	:	val_out <= 4'hfd14;
         4'h374b 	:	val_out <= 4'hfd14;
         4'h3750 	:	val_out <= 4'hfd19;
         4'h3751 	:	val_out <= 4'hfd19;
         4'h3752 	:	val_out <= 4'hfd19;
         4'h3753 	:	val_out <= 4'hfd19;
         4'h3758 	:	val_out <= 4'hfd1f;
         4'h3759 	:	val_out <= 4'hfd1f;
         4'h375a 	:	val_out <= 4'hfd1f;
         4'h375b 	:	val_out <= 4'hfd1f;
         4'h3760 	:	val_out <= 4'hfd24;
         4'h3761 	:	val_out <= 4'hfd24;
         4'h3762 	:	val_out <= 4'hfd24;
         4'h3763 	:	val_out <= 4'hfd24;
         4'h3768 	:	val_out <= 4'hfd29;
         4'h3769 	:	val_out <= 4'hfd29;
         4'h376a 	:	val_out <= 4'hfd29;
         4'h376b 	:	val_out <= 4'hfd29;
         4'h3770 	:	val_out <= 4'hfd2f;
         4'h3771 	:	val_out <= 4'hfd2f;
         4'h3772 	:	val_out <= 4'hfd2f;
         4'h3773 	:	val_out <= 4'hfd2f;
         4'h3778 	:	val_out <= 4'hfd34;
         4'h3779 	:	val_out <= 4'hfd34;
         4'h377a 	:	val_out <= 4'hfd34;
         4'h377b 	:	val_out <= 4'hfd34;
         4'h3780 	:	val_out <= 4'hfd39;
         4'h3781 	:	val_out <= 4'hfd39;
         4'h3782 	:	val_out <= 4'hfd39;
         4'h3783 	:	val_out <= 4'hfd39;
         4'h3788 	:	val_out <= 4'hfd3e;
         4'h3789 	:	val_out <= 4'hfd3e;
         4'h378a 	:	val_out <= 4'hfd3e;
         4'h378b 	:	val_out <= 4'hfd3e;
         4'h3790 	:	val_out <= 4'hfd43;
         4'h3791 	:	val_out <= 4'hfd43;
         4'h3792 	:	val_out <= 4'hfd43;
         4'h3793 	:	val_out <= 4'hfd43;
         4'h3798 	:	val_out <= 4'hfd49;
         4'h3799 	:	val_out <= 4'hfd49;
         4'h379a 	:	val_out <= 4'hfd49;
         4'h379b 	:	val_out <= 4'hfd49;
         4'h37a0 	:	val_out <= 4'hfd4e;
         4'h37a1 	:	val_out <= 4'hfd4e;
         4'h37a2 	:	val_out <= 4'hfd4e;
         4'h37a3 	:	val_out <= 4'hfd4e;
         4'h37a8 	:	val_out <= 4'hfd53;
         4'h37a9 	:	val_out <= 4'hfd53;
         4'h37aa 	:	val_out <= 4'hfd53;
         4'h37ab 	:	val_out <= 4'hfd53;
         4'h37b0 	:	val_out <= 4'hfd58;
         4'h37b1 	:	val_out <= 4'hfd58;
         4'h37b2 	:	val_out <= 4'hfd58;
         4'h37b3 	:	val_out <= 4'hfd58;
         4'h37b8 	:	val_out <= 4'hfd5d;
         4'h37b9 	:	val_out <= 4'hfd5d;
         4'h37ba 	:	val_out <= 4'hfd5d;
         4'h37bb 	:	val_out <= 4'hfd5d;
         4'h37c0 	:	val_out <= 4'hfd62;
         4'h37c1 	:	val_out <= 4'hfd62;
         4'h37c2 	:	val_out <= 4'hfd62;
         4'h37c3 	:	val_out <= 4'hfd62;
         4'h37c8 	:	val_out <= 4'hfd67;
         4'h37c9 	:	val_out <= 4'hfd67;
         4'h37ca 	:	val_out <= 4'hfd67;
         4'h37cb 	:	val_out <= 4'hfd67;
         4'h37d0 	:	val_out <= 4'hfd6c;
         4'h37d1 	:	val_out <= 4'hfd6c;
         4'h37d2 	:	val_out <= 4'hfd6c;
         4'h37d3 	:	val_out <= 4'hfd6c;
         4'h37d8 	:	val_out <= 4'hfd71;
         4'h37d9 	:	val_out <= 4'hfd71;
         4'h37da 	:	val_out <= 4'hfd71;
         4'h37db 	:	val_out <= 4'hfd71;
         4'h37e0 	:	val_out <= 4'hfd76;
         4'h37e1 	:	val_out <= 4'hfd76;
         4'h37e2 	:	val_out <= 4'hfd76;
         4'h37e3 	:	val_out <= 4'hfd76;
         4'h37e8 	:	val_out <= 4'hfd7b;
         4'h37e9 	:	val_out <= 4'hfd7b;
         4'h37ea 	:	val_out <= 4'hfd7b;
         4'h37eb 	:	val_out <= 4'hfd7b;
         4'h37f0 	:	val_out <= 4'hfd80;
         4'h37f1 	:	val_out <= 4'hfd80;
         4'h37f2 	:	val_out <= 4'hfd80;
         4'h37f3 	:	val_out <= 4'hfd80;
         4'h37f8 	:	val_out <= 4'hfd85;
         4'h37f9 	:	val_out <= 4'hfd85;
         4'h37fa 	:	val_out <= 4'hfd85;
         4'h37fb 	:	val_out <= 4'hfd85;
         4'h3800 	:	val_out <= 4'hfd8a;
         4'h3801 	:	val_out <= 4'hfd8a;
         4'h3802 	:	val_out <= 4'hfd8a;
         4'h3803 	:	val_out <= 4'hfd8a;
         4'h3808 	:	val_out <= 4'hfd8f;
         4'h3809 	:	val_out <= 4'hfd8f;
         4'h380a 	:	val_out <= 4'hfd8f;
         4'h380b 	:	val_out <= 4'hfd8f;
         4'h3810 	:	val_out <= 4'hfd94;
         4'h3811 	:	val_out <= 4'hfd94;
         4'h3812 	:	val_out <= 4'hfd94;
         4'h3813 	:	val_out <= 4'hfd94;
         4'h3818 	:	val_out <= 4'hfd98;
         4'h3819 	:	val_out <= 4'hfd98;
         4'h381a 	:	val_out <= 4'hfd98;
         4'h381b 	:	val_out <= 4'hfd98;
         4'h3820 	:	val_out <= 4'hfd9d;
         4'h3821 	:	val_out <= 4'hfd9d;
         4'h3822 	:	val_out <= 4'hfd9d;
         4'h3823 	:	val_out <= 4'hfd9d;
         4'h3828 	:	val_out <= 4'hfda2;
         4'h3829 	:	val_out <= 4'hfda2;
         4'h382a 	:	val_out <= 4'hfda2;
         4'h382b 	:	val_out <= 4'hfda2;
         4'h3830 	:	val_out <= 4'hfda7;
         4'h3831 	:	val_out <= 4'hfda7;
         4'h3832 	:	val_out <= 4'hfda7;
         4'h3833 	:	val_out <= 4'hfda7;
         4'h3838 	:	val_out <= 4'hfdac;
         4'h3839 	:	val_out <= 4'hfdac;
         4'h383a 	:	val_out <= 4'hfdac;
         4'h383b 	:	val_out <= 4'hfdac;
         4'h3840 	:	val_out <= 4'hfdb0;
         4'h3841 	:	val_out <= 4'hfdb0;
         4'h3842 	:	val_out <= 4'hfdb0;
         4'h3843 	:	val_out <= 4'hfdb0;
         4'h3848 	:	val_out <= 4'hfdb5;
         4'h3849 	:	val_out <= 4'hfdb5;
         4'h384a 	:	val_out <= 4'hfdb5;
         4'h384b 	:	val_out <= 4'hfdb5;
         4'h3850 	:	val_out <= 4'hfdba;
         4'h3851 	:	val_out <= 4'hfdba;
         4'h3852 	:	val_out <= 4'hfdba;
         4'h3853 	:	val_out <= 4'hfdba;
         4'h3858 	:	val_out <= 4'hfdbf;
         4'h3859 	:	val_out <= 4'hfdbf;
         4'h385a 	:	val_out <= 4'hfdbf;
         4'h385b 	:	val_out <= 4'hfdbf;
         4'h3860 	:	val_out <= 4'hfdc3;
         4'h3861 	:	val_out <= 4'hfdc3;
         4'h3862 	:	val_out <= 4'hfdc3;
         4'h3863 	:	val_out <= 4'hfdc3;
         4'h3868 	:	val_out <= 4'hfdc8;
         4'h3869 	:	val_out <= 4'hfdc8;
         4'h386a 	:	val_out <= 4'hfdc8;
         4'h386b 	:	val_out <= 4'hfdc8;
         4'h3870 	:	val_out <= 4'hfdcd;
         4'h3871 	:	val_out <= 4'hfdcd;
         4'h3872 	:	val_out <= 4'hfdcd;
         4'h3873 	:	val_out <= 4'hfdcd;
         4'h3878 	:	val_out <= 4'hfdd1;
         4'h3879 	:	val_out <= 4'hfdd1;
         4'h387a 	:	val_out <= 4'hfdd1;
         4'h387b 	:	val_out <= 4'hfdd1;
         4'h3880 	:	val_out <= 4'hfdd6;
         4'h3881 	:	val_out <= 4'hfdd6;
         4'h3882 	:	val_out <= 4'hfdd6;
         4'h3883 	:	val_out <= 4'hfdd6;
         4'h3888 	:	val_out <= 4'hfdda;
         4'h3889 	:	val_out <= 4'hfdda;
         4'h388a 	:	val_out <= 4'hfdda;
         4'h388b 	:	val_out <= 4'hfdda;
         4'h3890 	:	val_out <= 4'hfddf;
         4'h3891 	:	val_out <= 4'hfddf;
         4'h3892 	:	val_out <= 4'hfddf;
         4'h3893 	:	val_out <= 4'hfddf;
         4'h3898 	:	val_out <= 4'hfde4;
         4'h3899 	:	val_out <= 4'hfde4;
         4'h389a 	:	val_out <= 4'hfde4;
         4'h389b 	:	val_out <= 4'hfde4;
         4'h38a0 	:	val_out <= 4'hfde8;
         4'h38a1 	:	val_out <= 4'hfde8;
         4'h38a2 	:	val_out <= 4'hfde8;
         4'h38a3 	:	val_out <= 4'hfde8;
         4'h38a8 	:	val_out <= 4'hfded;
         4'h38a9 	:	val_out <= 4'hfded;
         4'h38aa 	:	val_out <= 4'hfded;
         4'h38ab 	:	val_out <= 4'hfded;
         4'h38b0 	:	val_out <= 4'hfdf1;
         4'h38b1 	:	val_out <= 4'hfdf1;
         4'h38b2 	:	val_out <= 4'hfdf1;
         4'h38b3 	:	val_out <= 4'hfdf1;
         4'h38b8 	:	val_out <= 4'hfdf6;
         4'h38b9 	:	val_out <= 4'hfdf6;
         4'h38ba 	:	val_out <= 4'hfdf6;
         4'h38bb 	:	val_out <= 4'hfdf6;
         4'h38c0 	:	val_out <= 4'hfdfa;
         4'h38c1 	:	val_out <= 4'hfdfa;
         4'h38c2 	:	val_out <= 4'hfdfa;
         4'h38c3 	:	val_out <= 4'hfdfa;
         4'h38c8 	:	val_out <= 4'hfdff;
         4'h38c9 	:	val_out <= 4'hfdff;
         4'h38ca 	:	val_out <= 4'hfdff;
         4'h38cb 	:	val_out <= 4'hfdff;
         4'h38d0 	:	val_out <= 4'hfe03;
         4'h38d1 	:	val_out <= 4'hfe03;
         4'h38d2 	:	val_out <= 4'hfe03;
         4'h38d3 	:	val_out <= 4'hfe03;
         4'h38d8 	:	val_out <= 4'hfe07;
         4'h38d9 	:	val_out <= 4'hfe07;
         4'h38da 	:	val_out <= 4'hfe07;
         4'h38db 	:	val_out <= 4'hfe07;
         4'h38e0 	:	val_out <= 4'hfe0c;
         4'h38e1 	:	val_out <= 4'hfe0c;
         4'h38e2 	:	val_out <= 4'hfe0c;
         4'h38e3 	:	val_out <= 4'hfe0c;
         4'h38e8 	:	val_out <= 4'hfe10;
         4'h38e9 	:	val_out <= 4'hfe10;
         4'h38ea 	:	val_out <= 4'hfe10;
         4'h38eb 	:	val_out <= 4'hfe10;
         4'h38f0 	:	val_out <= 4'hfe14;
         4'h38f1 	:	val_out <= 4'hfe14;
         4'h38f2 	:	val_out <= 4'hfe14;
         4'h38f3 	:	val_out <= 4'hfe14;
         4'h38f8 	:	val_out <= 4'hfe19;
         4'h38f9 	:	val_out <= 4'hfe19;
         4'h38fa 	:	val_out <= 4'hfe19;
         4'h38fb 	:	val_out <= 4'hfe19;
         4'h3900 	:	val_out <= 4'hfe1d;
         4'h3901 	:	val_out <= 4'hfe1d;
         4'h3902 	:	val_out <= 4'hfe1d;
         4'h3903 	:	val_out <= 4'hfe1d;
         4'h3908 	:	val_out <= 4'hfe21;
         4'h3909 	:	val_out <= 4'hfe21;
         4'h390a 	:	val_out <= 4'hfe21;
         4'h390b 	:	val_out <= 4'hfe21;
         4'h3910 	:	val_out <= 4'hfe26;
         4'h3911 	:	val_out <= 4'hfe26;
         4'h3912 	:	val_out <= 4'hfe26;
         4'h3913 	:	val_out <= 4'hfe26;
         4'h3918 	:	val_out <= 4'hfe2a;
         4'h3919 	:	val_out <= 4'hfe2a;
         4'h391a 	:	val_out <= 4'hfe2a;
         4'h391b 	:	val_out <= 4'hfe2a;
         4'h3920 	:	val_out <= 4'hfe2e;
         4'h3921 	:	val_out <= 4'hfe2e;
         4'h3922 	:	val_out <= 4'hfe2e;
         4'h3923 	:	val_out <= 4'hfe2e;
         4'h3928 	:	val_out <= 4'hfe32;
         4'h3929 	:	val_out <= 4'hfe32;
         4'h392a 	:	val_out <= 4'hfe32;
         4'h392b 	:	val_out <= 4'hfe32;
         4'h3930 	:	val_out <= 4'hfe37;
         4'h3931 	:	val_out <= 4'hfe37;
         4'h3932 	:	val_out <= 4'hfe37;
         4'h3933 	:	val_out <= 4'hfe37;
         4'h3938 	:	val_out <= 4'hfe3b;
         4'h3939 	:	val_out <= 4'hfe3b;
         4'h393a 	:	val_out <= 4'hfe3b;
         4'h393b 	:	val_out <= 4'hfe3b;
         4'h3940 	:	val_out <= 4'hfe3f;
         4'h3941 	:	val_out <= 4'hfe3f;
         4'h3942 	:	val_out <= 4'hfe3f;
         4'h3943 	:	val_out <= 4'hfe3f;
         4'h3948 	:	val_out <= 4'hfe43;
         4'h3949 	:	val_out <= 4'hfe43;
         4'h394a 	:	val_out <= 4'hfe43;
         4'h394b 	:	val_out <= 4'hfe43;
         4'h3950 	:	val_out <= 4'hfe47;
         4'h3951 	:	val_out <= 4'hfe47;
         4'h3952 	:	val_out <= 4'hfe47;
         4'h3953 	:	val_out <= 4'hfe47;
         4'h3958 	:	val_out <= 4'hfe4b;
         4'h3959 	:	val_out <= 4'hfe4b;
         4'h395a 	:	val_out <= 4'hfe4b;
         4'h395b 	:	val_out <= 4'hfe4b;
         4'h3960 	:	val_out <= 4'hfe4f;
         4'h3961 	:	val_out <= 4'hfe4f;
         4'h3962 	:	val_out <= 4'hfe4f;
         4'h3963 	:	val_out <= 4'hfe4f;
         4'h3968 	:	val_out <= 4'hfe53;
         4'h3969 	:	val_out <= 4'hfe53;
         4'h396a 	:	val_out <= 4'hfe53;
         4'h396b 	:	val_out <= 4'hfe53;
         4'h3970 	:	val_out <= 4'hfe57;
         4'h3971 	:	val_out <= 4'hfe57;
         4'h3972 	:	val_out <= 4'hfe57;
         4'h3973 	:	val_out <= 4'hfe57;
         4'h3978 	:	val_out <= 4'hfe5b;
         4'h3979 	:	val_out <= 4'hfe5b;
         4'h397a 	:	val_out <= 4'hfe5b;
         4'h397b 	:	val_out <= 4'hfe5b;
         4'h3980 	:	val_out <= 4'hfe5f;
         4'h3981 	:	val_out <= 4'hfe5f;
         4'h3982 	:	val_out <= 4'hfe5f;
         4'h3983 	:	val_out <= 4'hfe5f;
         4'h3988 	:	val_out <= 4'hfe63;
         4'h3989 	:	val_out <= 4'hfe63;
         4'h398a 	:	val_out <= 4'hfe63;
         4'h398b 	:	val_out <= 4'hfe63;
         4'h3990 	:	val_out <= 4'hfe67;
         4'h3991 	:	val_out <= 4'hfe67;
         4'h3992 	:	val_out <= 4'hfe67;
         4'h3993 	:	val_out <= 4'hfe67;
         4'h3998 	:	val_out <= 4'hfe6b;
         4'h3999 	:	val_out <= 4'hfe6b;
         4'h399a 	:	val_out <= 4'hfe6b;
         4'h399b 	:	val_out <= 4'hfe6b;
         4'h39a0 	:	val_out <= 4'hfe6f;
         4'h39a1 	:	val_out <= 4'hfe6f;
         4'h39a2 	:	val_out <= 4'hfe6f;
         4'h39a3 	:	val_out <= 4'hfe6f;
         4'h39a8 	:	val_out <= 4'hfe73;
         4'h39a9 	:	val_out <= 4'hfe73;
         4'h39aa 	:	val_out <= 4'hfe73;
         4'h39ab 	:	val_out <= 4'hfe73;
         4'h39b0 	:	val_out <= 4'hfe77;
         4'h39b1 	:	val_out <= 4'hfe77;
         4'h39b2 	:	val_out <= 4'hfe77;
         4'h39b3 	:	val_out <= 4'hfe77;
         4'h39b8 	:	val_out <= 4'hfe7b;
         4'h39b9 	:	val_out <= 4'hfe7b;
         4'h39ba 	:	val_out <= 4'hfe7b;
         4'h39bb 	:	val_out <= 4'hfe7b;
         4'h39c0 	:	val_out <= 4'hfe7f;
         4'h39c1 	:	val_out <= 4'hfe7f;
         4'h39c2 	:	val_out <= 4'hfe7f;
         4'h39c3 	:	val_out <= 4'hfe7f;
         4'h39c8 	:	val_out <= 4'hfe83;
         4'h39c9 	:	val_out <= 4'hfe83;
         4'h39ca 	:	val_out <= 4'hfe83;
         4'h39cb 	:	val_out <= 4'hfe83;
         4'h39d0 	:	val_out <= 4'hfe86;
         4'h39d1 	:	val_out <= 4'hfe86;
         4'h39d2 	:	val_out <= 4'hfe86;
         4'h39d3 	:	val_out <= 4'hfe86;
         4'h39d8 	:	val_out <= 4'hfe8a;
         4'h39d9 	:	val_out <= 4'hfe8a;
         4'h39da 	:	val_out <= 4'hfe8a;
         4'h39db 	:	val_out <= 4'hfe8a;
         4'h39e0 	:	val_out <= 4'hfe8e;
         4'h39e1 	:	val_out <= 4'hfe8e;
         4'h39e2 	:	val_out <= 4'hfe8e;
         4'h39e3 	:	val_out <= 4'hfe8e;
         4'h39e8 	:	val_out <= 4'hfe92;
         4'h39e9 	:	val_out <= 4'hfe92;
         4'h39ea 	:	val_out <= 4'hfe92;
         4'h39eb 	:	val_out <= 4'hfe92;
         4'h39f0 	:	val_out <= 4'hfe95;
         4'h39f1 	:	val_out <= 4'hfe95;
         4'h39f2 	:	val_out <= 4'hfe95;
         4'h39f3 	:	val_out <= 4'hfe95;
         4'h39f8 	:	val_out <= 4'hfe99;
         4'h39f9 	:	val_out <= 4'hfe99;
         4'h39fa 	:	val_out <= 4'hfe99;
         4'h39fb 	:	val_out <= 4'hfe99;
         4'h3a00 	:	val_out <= 4'hfe9d;
         4'h3a01 	:	val_out <= 4'hfe9d;
         4'h3a02 	:	val_out <= 4'hfe9d;
         4'h3a03 	:	val_out <= 4'hfe9d;
         4'h3a08 	:	val_out <= 4'hfea1;
         4'h3a09 	:	val_out <= 4'hfea1;
         4'h3a0a 	:	val_out <= 4'hfea1;
         4'h3a0b 	:	val_out <= 4'hfea1;
         4'h3a10 	:	val_out <= 4'hfea4;
         4'h3a11 	:	val_out <= 4'hfea4;
         4'h3a12 	:	val_out <= 4'hfea4;
         4'h3a13 	:	val_out <= 4'hfea4;
         4'h3a18 	:	val_out <= 4'hfea8;
         4'h3a19 	:	val_out <= 4'hfea8;
         4'h3a1a 	:	val_out <= 4'hfea8;
         4'h3a1b 	:	val_out <= 4'hfea8;
         4'h3a20 	:	val_out <= 4'hfeab;
         4'h3a21 	:	val_out <= 4'hfeab;
         4'h3a22 	:	val_out <= 4'hfeab;
         4'h3a23 	:	val_out <= 4'hfeab;
         4'h3a28 	:	val_out <= 4'hfeaf;
         4'h3a29 	:	val_out <= 4'hfeaf;
         4'h3a2a 	:	val_out <= 4'hfeaf;
         4'h3a2b 	:	val_out <= 4'hfeaf;
         4'h3a30 	:	val_out <= 4'hfeb3;
         4'h3a31 	:	val_out <= 4'hfeb3;
         4'h3a32 	:	val_out <= 4'hfeb3;
         4'h3a33 	:	val_out <= 4'hfeb3;
         4'h3a38 	:	val_out <= 4'hfeb6;
         4'h3a39 	:	val_out <= 4'hfeb6;
         4'h3a3a 	:	val_out <= 4'hfeb6;
         4'h3a3b 	:	val_out <= 4'hfeb6;
         4'h3a40 	:	val_out <= 4'hfeba;
         4'h3a41 	:	val_out <= 4'hfeba;
         4'h3a42 	:	val_out <= 4'hfeba;
         4'h3a43 	:	val_out <= 4'hfeba;
         4'h3a48 	:	val_out <= 4'hfebd;
         4'h3a49 	:	val_out <= 4'hfebd;
         4'h3a4a 	:	val_out <= 4'hfebd;
         4'h3a4b 	:	val_out <= 4'hfebd;
         4'h3a50 	:	val_out <= 4'hfec1;
         4'h3a51 	:	val_out <= 4'hfec1;
         4'h3a52 	:	val_out <= 4'hfec1;
         4'h3a53 	:	val_out <= 4'hfec1;
         4'h3a58 	:	val_out <= 4'hfec4;
         4'h3a59 	:	val_out <= 4'hfec4;
         4'h3a5a 	:	val_out <= 4'hfec4;
         4'h3a5b 	:	val_out <= 4'hfec4;
         4'h3a60 	:	val_out <= 4'hfec8;
         4'h3a61 	:	val_out <= 4'hfec8;
         4'h3a62 	:	val_out <= 4'hfec8;
         4'h3a63 	:	val_out <= 4'hfec8;
         4'h3a68 	:	val_out <= 4'hfecb;
         4'h3a69 	:	val_out <= 4'hfecb;
         4'h3a6a 	:	val_out <= 4'hfecb;
         4'h3a6b 	:	val_out <= 4'hfecb;
         4'h3a70 	:	val_out <= 4'hfecf;
         4'h3a71 	:	val_out <= 4'hfecf;
         4'h3a72 	:	val_out <= 4'hfecf;
         4'h3a73 	:	val_out <= 4'hfecf;
         4'h3a78 	:	val_out <= 4'hfed2;
         4'h3a79 	:	val_out <= 4'hfed2;
         4'h3a7a 	:	val_out <= 4'hfed2;
         4'h3a7b 	:	val_out <= 4'hfed2;
         4'h3a80 	:	val_out <= 4'hfed5;
         4'h3a81 	:	val_out <= 4'hfed5;
         4'h3a82 	:	val_out <= 4'hfed5;
         4'h3a83 	:	val_out <= 4'hfed5;
         4'h3a88 	:	val_out <= 4'hfed9;
         4'h3a89 	:	val_out <= 4'hfed9;
         4'h3a8a 	:	val_out <= 4'hfed9;
         4'h3a8b 	:	val_out <= 4'hfed9;
         4'h3a90 	:	val_out <= 4'hfedc;
         4'h3a91 	:	val_out <= 4'hfedc;
         4'h3a92 	:	val_out <= 4'hfedc;
         4'h3a93 	:	val_out <= 4'hfedc;
         4'h3a98 	:	val_out <= 4'hfedf;
         4'h3a99 	:	val_out <= 4'hfedf;
         4'h3a9a 	:	val_out <= 4'hfedf;
         4'h3a9b 	:	val_out <= 4'hfedf;
         4'h3aa0 	:	val_out <= 4'hfee3;
         4'h3aa1 	:	val_out <= 4'hfee3;
         4'h3aa2 	:	val_out <= 4'hfee3;
         4'h3aa3 	:	val_out <= 4'hfee3;
         4'h3aa8 	:	val_out <= 4'hfee6;
         4'h3aa9 	:	val_out <= 4'hfee6;
         4'h3aaa 	:	val_out <= 4'hfee6;
         4'h3aab 	:	val_out <= 4'hfee6;
         4'h3ab0 	:	val_out <= 4'hfee9;
         4'h3ab1 	:	val_out <= 4'hfee9;
         4'h3ab2 	:	val_out <= 4'hfee9;
         4'h3ab3 	:	val_out <= 4'hfee9;
         4'h3ab8 	:	val_out <= 4'hfeed;
         4'h3ab9 	:	val_out <= 4'hfeed;
         4'h3aba 	:	val_out <= 4'hfeed;
         4'h3abb 	:	val_out <= 4'hfeed;
         4'h3ac0 	:	val_out <= 4'hfef0;
         4'h3ac1 	:	val_out <= 4'hfef0;
         4'h3ac2 	:	val_out <= 4'hfef0;
         4'h3ac3 	:	val_out <= 4'hfef0;
         4'h3ac8 	:	val_out <= 4'hfef3;
         4'h3ac9 	:	val_out <= 4'hfef3;
         4'h3aca 	:	val_out <= 4'hfef3;
         4'h3acb 	:	val_out <= 4'hfef3;
         4'h3ad0 	:	val_out <= 4'hfef6;
         4'h3ad1 	:	val_out <= 4'hfef6;
         4'h3ad2 	:	val_out <= 4'hfef6;
         4'h3ad3 	:	val_out <= 4'hfef6;
         4'h3ad8 	:	val_out <= 4'hfef9;
         4'h3ad9 	:	val_out <= 4'hfef9;
         4'h3ada 	:	val_out <= 4'hfef9;
         4'h3adb 	:	val_out <= 4'hfef9;
         4'h3ae0 	:	val_out <= 4'hfefd;
         4'h3ae1 	:	val_out <= 4'hfefd;
         4'h3ae2 	:	val_out <= 4'hfefd;
         4'h3ae3 	:	val_out <= 4'hfefd;
         4'h3ae8 	:	val_out <= 4'hff00;
         4'h3ae9 	:	val_out <= 4'hff00;
         4'h3aea 	:	val_out <= 4'hff00;
         4'h3aeb 	:	val_out <= 4'hff00;
         4'h3af0 	:	val_out <= 4'hff03;
         4'h3af1 	:	val_out <= 4'hff03;
         4'h3af2 	:	val_out <= 4'hff03;
         4'h3af3 	:	val_out <= 4'hff03;
         4'h3af8 	:	val_out <= 4'hff06;
         4'h3af9 	:	val_out <= 4'hff06;
         4'h3afa 	:	val_out <= 4'hff06;
         4'h3afb 	:	val_out <= 4'hff06;
         4'h3b00 	:	val_out <= 4'hff09;
         4'h3b01 	:	val_out <= 4'hff09;
         4'h3b02 	:	val_out <= 4'hff09;
         4'h3b03 	:	val_out <= 4'hff09;
         4'h3b08 	:	val_out <= 4'hff0c;
         4'h3b09 	:	val_out <= 4'hff0c;
         4'h3b0a 	:	val_out <= 4'hff0c;
         4'h3b0b 	:	val_out <= 4'hff0c;
         4'h3b10 	:	val_out <= 4'hff0f;
         4'h3b11 	:	val_out <= 4'hff0f;
         4'h3b12 	:	val_out <= 4'hff0f;
         4'h3b13 	:	val_out <= 4'hff0f;
         4'h3b18 	:	val_out <= 4'hff12;
         4'h3b19 	:	val_out <= 4'hff12;
         4'h3b1a 	:	val_out <= 4'hff12;
         4'h3b1b 	:	val_out <= 4'hff12;
         4'h3b20 	:	val_out <= 4'hff15;
         4'h3b21 	:	val_out <= 4'hff15;
         4'h3b22 	:	val_out <= 4'hff15;
         4'h3b23 	:	val_out <= 4'hff15;
         4'h3b28 	:	val_out <= 4'hff18;
         4'h3b29 	:	val_out <= 4'hff18;
         4'h3b2a 	:	val_out <= 4'hff18;
         4'h3b2b 	:	val_out <= 4'hff18;
         4'h3b30 	:	val_out <= 4'hff1b;
         4'h3b31 	:	val_out <= 4'hff1b;
         4'h3b32 	:	val_out <= 4'hff1b;
         4'h3b33 	:	val_out <= 4'hff1b;
         4'h3b38 	:	val_out <= 4'hff1e;
         4'h3b39 	:	val_out <= 4'hff1e;
         4'h3b3a 	:	val_out <= 4'hff1e;
         4'h3b3b 	:	val_out <= 4'hff1e;
         4'h3b40 	:	val_out <= 4'hff21;
         4'h3b41 	:	val_out <= 4'hff21;
         4'h3b42 	:	val_out <= 4'hff21;
         4'h3b43 	:	val_out <= 4'hff21;
         4'h3b48 	:	val_out <= 4'hff24;
         4'h3b49 	:	val_out <= 4'hff24;
         4'h3b4a 	:	val_out <= 4'hff24;
         4'h3b4b 	:	val_out <= 4'hff24;
         4'h3b50 	:	val_out <= 4'hff27;
         4'h3b51 	:	val_out <= 4'hff27;
         4'h3b52 	:	val_out <= 4'hff27;
         4'h3b53 	:	val_out <= 4'hff27;
         4'h3b58 	:	val_out <= 4'hff2a;
         4'h3b59 	:	val_out <= 4'hff2a;
         4'h3b5a 	:	val_out <= 4'hff2a;
         4'h3b5b 	:	val_out <= 4'hff2a;
         4'h3b60 	:	val_out <= 4'hff2d;
         4'h3b61 	:	val_out <= 4'hff2d;
         4'h3b62 	:	val_out <= 4'hff2d;
         4'h3b63 	:	val_out <= 4'hff2d;
         4'h3b68 	:	val_out <= 4'hff2f;
         4'h3b69 	:	val_out <= 4'hff2f;
         4'h3b6a 	:	val_out <= 4'hff2f;
         4'h3b6b 	:	val_out <= 4'hff2f;
         4'h3b70 	:	val_out <= 4'hff32;
         4'h3b71 	:	val_out <= 4'hff32;
         4'h3b72 	:	val_out <= 4'hff32;
         4'h3b73 	:	val_out <= 4'hff32;
         4'h3b78 	:	val_out <= 4'hff35;
         4'h3b79 	:	val_out <= 4'hff35;
         4'h3b7a 	:	val_out <= 4'hff35;
         4'h3b7b 	:	val_out <= 4'hff35;
         4'h3b80 	:	val_out <= 4'hff38;
         4'h3b81 	:	val_out <= 4'hff38;
         4'h3b82 	:	val_out <= 4'hff38;
         4'h3b83 	:	val_out <= 4'hff38;
         4'h3b88 	:	val_out <= 4'hff3b;
         4'h3b89 	:	val_out <= 4'hff3b;
         4'h3b8a 	:	val_out <= 4'hff3b;
         4'h3b8b 	:	val_out <= 4'hff3b;
         4'h3b90 	:	val_out <= 4'hff3d;
         4'h3b91 	:	val_out <= 4'hff3d;
         4'h3b92 	:	val_out <= 4'hff3d;
         4'h3b93 	:	val_out <= 4'hff3d;
         4'h3b98 	:	val_out <= 4'hff40;
         4'h3b99 	:	val_out <= 4'hff40;
         4'h3b9a 	:	val_out <= 4'hff40;
         4'h3b9b 	:	val_out <= 4'hff40;
         4'h3ba0 	:	val_out <= 4'hff43;
         4'h3ba1 	:	val_out <= 4'hff43;
         4'h3ba2 	:	val_out <= 4'hff43;
         4'h3ba3 	:	val_out <= 4'hff43;
         4'h3ba8 	:	val_out <= 4'hff45;
         4'h3ba9 	:	val_out <= 4'hff45;
         4'h3baa 	:	val_out <= 4'hff45;
         4'h3bab 	:	val_out <= 4'hff45;
         4'h3bb0 	:	val_out <= 4'hff48;
         4'h3bb1 	:	val_out <= 4'hff48;
         4'h3bb2 	:	val_out <= 4'hff48;
         4'h3bb3 	:	val_out <= 4'hff48;
         4'h3bb8 	:	val_out <= 4'hff4b;
         4'h3bb9 	:	val_out <= 4'hff4b;
         4'h3bba 	:	val_out <= 4'hff4b;
         4'h3bbb 	:	val_out <= 4'hff4b;
         4'h3bc0 	:	val_out <= 4'hff4d;
         4'h3bc1 	:	val_out <= 4'hff4d;
         4'h3bc2 	:	val_out <= 4'hff4d;
         4'h3bc3 	:	val_out <= 4'hff4d;
         4'h3bc8 	:	val_out <= 4'hff50;
         4'h3bc9 	:	val_out <= 4'hff50;
         4'h3bca 	:	val_out <= 4'hff50;
         4'h3bcb 	:	val_out <= 4'hff50;
         4'h3bd0 	:	val_out <= 4'hff53;
         4'h3bd1 	:	val_out <= 4'hff53;
         4'h3bd2 	:	val_out <= 4'hff53;
         4'h3bd3 	:	val_out <= 4'hff53;
         4'h3bd8 	:	val_out <= 4'hff55;
         4'h3bd9 	:	val_out <= 4'hff55;
         4'h3bda 	:	val_out <= 4'hff55;
         4'h3bdb 	:	val_out <= 4'hff55;
         4'h3be0 	:	val_out <= 4'hff58;
         4'h3be1 	:	val_out <= 4'hff58;
         4'h3be2 	:	val_out <= 4'hff58;
         4'h3be3 	:	val_out <= 4'hff58;
         4'h3be8 	:	val_out <= 4'hff5a;
         4'h3be9 	:	val_out <= 4'hff5a;
         4'h3bea 	:	val_out <= 4'hff5a;
         4'h3beb 	:	val_out <= 4'hff5a;
         4'h3bf0 	:	val_out <= 4'hff5d;
         4'h3bf1 	:	val_out <= 4'hff5d;
         4'h3bf2 	:	val_out <= 4'hff5d;
         4'h3bf3 	:	val_out <= 4'hff5d;
         4'h3bf8 	:	val_out <= 4'hff5f;
         4'h3bf9 	:	val_out <= 4'hff5f;
         4'h3bfa 	:	val_out <= 4'hff5f;
         4'h3bfb 	:	val_out <= 4'hff5f;
         4'h3c00 	:	val_out <= 4'hff62;
         4'h3c01 	:	val_out <= 4'hff62;
         4'h3c02 	:	val_out <= 4'hff62;
         4'h3c03 	:	val_out <= 4'hff62;
         4'h3c08 	:	val_out <= 4'hff64;
         4'h3c09 	:	val_out <= 4'hff64;
         4'h3c0a 	:	val_out <= 4'hff64;
         4'h3c0b 	:	val_out <= 4'hff64;
         4'h3c10 	:	val_out <= 4'hff67;
         4'h3c11 	:	val_out <= 4'hff67;
         4'h3c12 	:	val_out <= 4'hff67;
         4'h3c13 	:	val_out <= 4'hff67;
         4'h3c18 	:	val_out <= 4'hff69;
         4'h3c19 	:	val_out <= 4'hff69;
         4'h3c1a 	:	val_out <= 4'hff69;
         4'h3c1b 	:	val_out <= 4'hff69;
         4'h3c20 	:	val_out <= 4'hff6b;
         4'h3c21 	:	val_out <= 4'hff6b;
         4'h3c22 	:	val_out <= 4'hff6b;
         4'h3c23 	:	val_out <= 4'hff6b;
         4'h3c28 	:	val_out <= 4'hff6e;
         4'h3c29 	:	val_out <= 4'hff6e;
         4'h3c2a 	:	val_out <= 4'hff6e;
         4'h3c2b 	:	val_out <= 4'hff6e;
         4'h3c30 	:	val_out <= 4'hff70;
         4'h3c31 	:	val_out <= 4'hff70;
         4'h3c32 	:	val_out <= 4'hff70;
         4'h3c33 	:	val_out <= 4'hff70;
         4'h3c38 	:	val_out <= 4'hff72;
         4'h3c39 	:	val_out <= 4'hff72;
         4'h3c3a 	:	val_out <= 4'hff72;
         4'h3c3b 	:	val_out <= 4'hff72;
         4'h3c40 	:	val_out <= 4'hff75;
         4'h3c41 	:	val_out <= 4'hff75;
         4'h3c42 	:	val_out <= 4'hff75;
         4'h3c43 	:	val_out <= 4'hff75;
         4'h3c48 	:	val_out <= 4'hff77;
         4'h3c49 	:	val_out <= 4'hff77;
         4'h3c4a 	:	val_out <= 4'hff77;
         4'h3c4b 	:	val_out <= 4'hff77;
         4'h3c50 	:	val_out <= 4'hff79;
         4'h3c51 	:	val_out <= 4'hff79;
         4'h3c52 	:	val_out <= 4'hff79;
         4'h3c53 	:	val_out <= 4'hff79;
         4'h3c58 	:	val_out <= 4'hff7c;
         4'h3c59 	:	val_out <= 4'hff7c;
         4'h3c5a 	:	val_out <= 4'hff7c;
         4'h3c5b 	:	val_out <= 4'hff7c;
         4'h3c60 	:	val_out <= 4'hff7e;
         4'h3c61 	:	val_out <= 4'hff7e;
         4'h3c62 	:	val_out <= 4'hff7e;
         4'h3c63 	:	val_out <= 4'hff7e;
         4'h3c68 	:	val_out <= 4'hff80;
         4'h3c69 	:	val_out <= 4'hff80;
         4'h3c6a 	:	val_out <= 4'hff80;
         4'h3c6b 	:	val_out <= 4'hff80;
         4'h3c70 	:	val_out <= 4'hff82;
         4'h3c71 	:	val_out <= 4'hff82;
         4'h3c72 	:	val_out <= 4'hff82;
         4'h3c73 	:	val_out <= 4'hff82;
         4'h3c78 	:	val_out <= 4'hff85;
         4'h3c79 	:	val_out <= 4'hff85;
         4'h3c7a 	:	val_out <= 4'hff85;
         4'h3c7b 	:	val_out <= 4'hff85;
         4'h3c80 	:	val_out <= 4'hff87;
         4'h3c81 	:	val_out <= 4'hff87;
         4'h3c82 	:	val_out <= 4'hff87;
         4'h3c83 	:	val_out <= 4'hff87;
         4'h3c88 	:	val_out <= 4'hff89;
         4'h3c89 	:	val_out <= 4'hff89;
         4'h3c8a 	:	val_out <= 4'hff89;
         4'h3c8b 	:	val_out <= 4'hff89;
         4'h3c90 	:	val_out <= 4'hff8b;
         4'h3c91 	:	val_out <= 4'hff8b;
         4'h3c92 	:	val_out <= 4'hff8b;
         4'h3c93 	:	val_out <= 4'hff8b;
         4'h3c98 	:	val_out <= 4'hff8d;
         4'h3c99 	:	val_out <= 4'hff8d;
         4'h3c9a 	:	val_out <= 4'hff8d;
         4'h3c9b 	:	val_out <= 4'hff8d;
         4'h3ca0 	:	val_out <= 4'hff8f;
         4'h3ca1 	:	val_out <= 4'hff8f;
         4'h3ca2 	:	val_out <= 4'hff8f;
         4'h3ca3 	:	val_out <= 4'hff8f;
         4'h3ca8 	:	val_out <= 4'hff91;
         4'h3ca9 	:	val_out <= 4'hff91;
         4'h3caa 	:	val_out <= 4'hff91;
         4'h3cab 	:	val_out <= 4'hff91;
         4'h3cb0 	:	val_out <= 4'hff93;
         4'h3cb1 	:	val_out <= 4'hff93;
         4'h3cb2 	:	val_out <= 4'hff93;
         4'h3cb3 	:	val_out <= 4'hff93;
         4'h3cb8 	:	val_out <= 4'hff95;
         4'h3cb9 	:	val_out <= 4'hff95;
         4'h3cba 	:	val_out <= 4'hff95;
         4'h3cbb 	:	val_out <= 4'hff95;
         4'h3cc0 	:	val_out <= 4'hff97;
         4'h3cc1 	:	val_out <= 4'hff97;
         4'h3cc2 	:	val_out <= 4'hff97;
         4'h3cc3 	:	val_out <= 4'hff97;
         4'h3cc8 	:	val_out <= 4'hff99;
         4'h3cc9 	:	val_out <= 4'hff99;
         4'h3cca 	:	val_out <= 4'hff99;
         4'h3ccb 	:	val_out <= 4'hff99;
         4'h3cd0 	:	val_out <= 4'hff9b;
         4'h3cd1 	:	val_out <= 4'hff9b;
         4'h3cd2 	:	val_out <= 4'hff9b;
         4'h3cd3 	:	val_out <= 4'hff9b;
         4'h3cd8 	:	val_out <= 4'hff9d;
         4'h3cd9 	:	val_out <= 4'hff9d;
         4'h3cda 	:	val_out <= 4'hff9d;
         4'h3cdb 	:	val_out <= 4'hff9d;
         4'h3ce0 	:	val_out <= 4'hff9f;
         4'h3ce1 	:	val_out <= 4'hff9f;
         4'h3ce2 	:	val_out <= 4'hff9f;
         4'h3ce3 	:	val_out <= 4'hff9f;
         4'h3ce8 	:	val_out <= 4'hffa1;
         4'h3ce9 	:	val_out <= 4'hffa1;
         4'h3cea 	:	val_out <= 4'hffa1;
         4'h3ceb 	:	val_out <= 4'hffa1;
         4'h3cf0 	:	val_out <= 4'hffa3;
         4'h3cf1 	:	val_out <= 4'hffa3;
         4'h3cf2 	:	val_out <= 4'hffa3;
         4'h3cf3 	:	val_out <= 4'hffa3;
         4'h3cf8 	:	val_out <= 4'hffa5;
         4'h3cf9 	:	val_out <= 4'hffa5;
         4'h3cfa 	:	val_out <= 4'hffa5;
         4'h3cfb 	:	val_out <= 4'hffa5;
         4'h3d00 	:	val_out <= 4'hffa7;
         4'h3d01 	:	val_out <= 4'hffa7;
         4'h3d02 	:	val_out <= 4'hffa7;
         4'h3d03 	:	val_out <= 4'hffa7;
         4'h3d08 	:	val_out <= 4'hffa9;
         4'h3d09 	:	val_out <= 4'hffa9;
         4'h3d0a 	:	val_out <= 4'hffa9;
         4'h3d0b 	:	val_out <= 4'hffa9;
         4'h3d10 	:	val_out <= 4'hffaa;
         4'h3d11 	:	val_out <= 4'hffaa;
         4'h3d12 	:	val_out <= 4'hffaa;
         4'h3d13 	:	val_out <= 4'hffaa;
         4'h3d18 	:	val_out <= 4'hffac;
         4'h3d19 	:	val_out <= 4'hffac;
         4'h3d1a 	:	val_out <= 4'hffac;
         4'h3d1b 	:	val_out <= 4'hffac;
         4'h3d20 	:	val_out <= 4'hffae;
         4'h3d21 	:	val_out <= 4'hffae;
         4'h3d22 	:	val_out <= 4'hffae;
         4'h3d23 	:	val_out <= 4'hffae;
         4'h3d28 	:	val_out <= 4'hffb0;
         4'h3d29 	:	val_out <= 4'hffb0;
         4'h3d2a 	:	val_out <= 4'hffb0;
         4'h3d2b 	:	val_out <= 4'hffb0;
         4'h3d30 	:	val_out <= 4'hffb1;
         4'h3d31 	:	val_out <= 4'hffb1;
         4'h3d32 	:	val_out <= 4'hffb1;
         4'h3d33 	:	val_out <= 4'hffb1;
         4'h3d38 	:	val_out <= 4'hffb3;
         4'h3d39 	:	val_out <= 4'hffb3;
         4'h3d3a 	:	val_out <= 4'hffb3;
         4'h3d3b 	:	val_out <= 4'hffb3;
         4'h3d40 	:	val_out <= 4'hffb5;
         4'h3d41 	:	val_out <= 4'hffb5;
         4'h3d42 	:	val_out <= 4'hffb5;
         4'h3d43 	:	val_out <= 4'hffb5;
         4'h3d48 	:	val_out <= 4'hffb7;
         4'h3d49 	:	val_out <= 4'hffb7;
         4'h3d4a 	:	val_out <= 4'hffb7;
         4'h3d4b 	:	val_out <= 4'hffb7;
         4'h3d50 	:	val_out <= 4'hffb8;
         4'h3d51 	:	val_out <= 4'hffb8;
         4'h3d52 	:	val_out <= 4'hffb8;
         4'h3d53 	:	val_out <= 4'hffb8;
         4'h3d58 	:	val_out <= 4'hffba;
         4'h3d59 	:	val_out <= 4'hffba;
         4'h3d5a 	:	val_out <= 4'hffba;
         4'h3d5b 	:	val_out <= 4'hffba;
         4'h3d60 	:	val_out <= 4'hffbc;
         4'h3d61 	:	val_out <= 4'hffbc;
         4'h3d62 	:	val_out <= 4'hffbc;
         4'h3d63 	:	val_out <= 4'hffbc;
         4'h3d68 	:	val_out <= 4'hffbd;
         4'h3d69 	:	val_out <= 4'hffbd;
         4'h3d6a 	:	val_out <= 4'hffbd;
         4'h3d6b 	:	val_out <= 4'hffbd;
         4'h3d70 	:	val_out <= 4'hffbf;
         4'h3d71 	:	val_out <= 4'hffbf;
         4'h3d72 	:	val_out <= 4'hffbf;
         4'h3d73 	:	val_out <= 4'hffbf;
         4'h3d78 	:	val_out <= 4'hffc0;
         4'h3d79 	:	val_out <= 4'hffc0;
         4'h3d7a 	:	val_out <= 4'hffc0;
         4'h3d7b 	:	val_out <= 4'hffc0;
         4'h3d80 	:	val_out <= 4'hffc2;
         4'h3d81 	:	val_out <= 4'hffc2;
         4'h3d82 	:	val_out <= 4'hffc2;
         4'h3d83 	:	val_out <= 4'hffc2;
         4'h3d88 	:	val_out <= 4'hffc3;
         4'h3d89 	:	val_out <= 4'hffc3;
         4'h3d8a 	:	val_out <= 4'hffc3;
         4'h3d8b 	:	val_out <= 4'hffc3;
         4'h3d90 	:	val_out <= 4'hffc5;
         4'h3d91 	:	val_out <= 4'hffc5;
         4'h3d92 	:	val_out <= 4'hffc5;
         4'h3d93 	:	val_out <= 4'hffc5;
         4'h3d98 	:	val_out <= 4'hffc6;
         4'h3d99 	:	val_out <= 4'hffc6;
         4'h3d9a 	:	val_out <= 4'hffc6;
         4'h3d9b 	:	val_out <= 4'hffc6;
         4'h3da0 	:	val_out <= 4'hffc8;
         4'h3da1 	:	val_out <= 4'hffc8;
         4'h3da2 	:	val_out <= 4'hffc8;
         4'h3da3 	:	val_out <= 4'hffc8;
         4'h3da8 	:	val_out <= 4'hffc9;
         4'h3da9 	:	val_out <= 4'hffc9;
         4'h3daa 	:	val_out <= 4'hffc9;
         4'h3dab 	:	val_out <= 4'hffc9;
         4'h3db0 	:	val_out <= 4'hffcb;
         4'h3db1 	:	val_out <= 4'hffcb;
         4'h3db2 	:	val_out <= 4'hffcb;
         4'h3db3 	:	val_out <= 4'hffcb;
         4'h3db8 	:	val_out <= 4'hffcc;
         4'h3db9 	:	val_out <= 4'hffcc;
         4'h3dba 	:	val_out <= 4'hffcc;
         4'h3dbb 	:	val_out <= 4'hffcc;
         4'h3dc0 	:	val_out <= 4'hffce;
         4'h3dc1 	:	val_out <= 4'hffce;
         4'h3dc2 	:	val_out <= 4'hffce;
         4'h3dc3 	:	val_out <= 4'hffce;
         4'h3dc8 	:	val_out <= 4'hffcf;
         4'h3dc9 	:	val_out <= 4'hffcf;
         4'h3dca 	:	val_out <= 4'hffcf;
         4'h3dcb 	:	val_out <= 4'hffcf;
         4'h3dd0 	:	val_out <= 4'hffd0;
         4'h3dd1 	:	val_out <= 4'hffd0;
         4'h3dd2 	:	val_out <= 4'hffd0;
         4'h3dd3 	:	val_out <= 4'hffd0;
         4'h3dd8 	:	val_out <= 4'hffd2;
         4'h3dd9 	:	val_out <= 4'hffd2;
         4'h3dda 	:	val_out <= 4'hffd2;
         4'h3ddb 	:	val_out <= 4'hffd2;
         4'h3de0 	:	val_out <= 4'hffd3;
         4'h3de1 	:	val_out <= 4'hffd3;
         4'h3de2 	:	val_out <= 4'hffd3;
         4'h3de3 	:	val_out <= 4'hffd3;
         4'h3de8 	:	val_out <= 4'hffd4;
         4'h3de9 	:	val_out <= 4'hffd4;
         4'h3dea 	:	val_out <= 4'hffd4;
         4'h3deb 	:	val_out <= 4'hffd4;
         4'h3df0 	:	val_out <= 4'hffd6;
         4'h3df1 	:	val_out <= 4'hffd6;
         4'h3df2 	:	val_out <= 4'hffd6;
         4'h3df3 	:	val_out <= 4'hffd6;
         4'h3df8 	:	val_out <= 4'hffd7;
         4'h3df9 	:	val_out <= 4'hffd7;
         4'h3dfa 	:	val_out <= 4'hffd7;
         4'h3dfb 	:	val_out <= 4'hffd7;
         4'h3e00 	:	val_out <= 4'hffd8;
         4'h3e01 	:	val_out <= 4'hffd8;
         4'h3e02 	:	val_out <= 4'hffd8;
         4'h3e03 	:	val_out <= 4'hffd8;
         4'h3e08 	:	val_out <= 4'hffd9;
         4'h3e09 	:	val_out <= 4'hffd9;
         4'h3e0a 	:	val_out <= 4'hffd9;
         4'h3e0b 	:	val_out <= 4'hffd9;
         4'h3e10 	:	val_out <= 4'hffda;
         4'h3e11 	:	val_out <= 4'hffda;
         4'h3e12 	:	val_out <= 4'hffda;
         4'h3e13 	:	val_out <= 4'hffda;
         4'h3e18 	:	val_out <= 4'hffdc;
         4'h3e19 	:	val_out <= 4'hffdc;
         4'h3e1a 	:	val_out <= 4'hffdc;
         4'h3e1b 	:	val_out <= 4'hffdc;
         4'h3e20 	:	val_out <= 4'hffdd;
         4'h3e21 	:	val_out <= 4'hffdd;
         4'h3e22 	:	val_out <= 4'hffdd;
         4'h3e23 	:	val_out <= 4'hffdd;
         4'h3e28 	:	val_out <= 4'hffde;
         4'h3e29 	:	val_out <= 4'hffde;
         4'h3e2a 	:	val_out <= 4'hffde;
         4'h3e2b 	:	val_out <= 4'hffde;
         4'h3e30 	:	val_out <= 4'hffdf;
         4'h3e31 	:	val_out <= 4'hffdf;
         4'h3e32 	:	val_out <= 4'hffdf;
         4'h3e33 	:	val_out <= 4'hffdf;
         4'h3e38 	:	val_out <= 4'hffe0;
         4'h3e39 	:	val_out <= 4'hffe0;
         4'h3e3a 	:	val_out <= 4'hffe0;
         4'h3e3b 	:	val_out <= 4'hffe0;
         4'h3e40 	:	val_out <= 4'hffe1;
         4'h3e41 	:	val_out <= 4'hffe1;
         4'h3e42 	:	val_out <= 4'hffe1;
         4'h3e43 	:	val_out <= 4'hffe1;
         4'h3e48 	:	val_out <= 4'hffe2;
         4'h3e49 	:	val_out <= 4'hffe2;
         4'h3e4a 	:	val_out <= 4'hffe2;
         4'h3e4b 	:	val_out <= 4'hffe2;
         4'h3e50 	:	val_out <= 4'hffe3;
         4'h3e51 	:	val_out <= 4'hffe3;
         4'h3e52 	:	val_out <= 4'hffe3;
         4'h3e53 	:	val_out <= 4'hffe3;
         4'h3e58 	:	val_out <= 4'hffe4;
         4'h3e59 	:	val_out <= 4'hffe4;
         4'h3e5a 	:	val_out <= 4'hffe4;
         4'h3e5b 	:	val_out <= 4'hffe4;
         4'h3e60 	:	val_out <= 4'hffe5;
         4'h3e61 	:	val_out <= 4'hffe5;
         4'h3e62 	:	val_out <= 4'hffe5;
         4'h3e63 	:	val_out <= 4'hffe5;
         4'h3e68 	:	val_out <= 4'hffe6;
         4'h3e69 	:	val_out <= 4'hffe6;
         4'h3e6a 	:	val_out <= 4'hffe6;
         4'h3e6b 	:	val_out <= 4'hffe6;
         4'h3e70 	:	val_out <= 4'hffe7;
         4'h3e71 	:	val_out <= 4'hffe7;
         4'h3e72 	:	val_out <= 4'hffe7;
         4'h3e73 	:	val_out <= 4'hffe7;
         4'h3e78 	:	val_out <= 4'hffe8;
         4'h3e79 	:	val_out <= 4'hffe8;
         4'h3e7a 	:	val_out <= 4'hffe8;
         4'h3e7b 	:	val_out <= 4'hffe8;
         4'h3e80 	:	val_out <= 4'hffe9;
         4'h3e81 	:	val_out <= 4'hffe9;
         4'h3e82 	:	val_out <= 4'hffe9;
         4'h3e83 	:	val_out <= 4'hffe9;
         4'h3e88 	:	val_out <= 4'hffea;
         4'h3e89 	:	val_out <= 4'hffea;
         4'h3e8a 	:	val_out <= 4'hffea;
         4'h3e8b 	:	val_out <= 4'hffea;
         4'h3e90 	:	val_out <= 4'hffeb;
         4'h3e91 	:	val_out <= 4'hffeb;
         4'h3e92 	:	val_out <= 4'hffeb;
         4'h3e93 	:	val_out <= 4'hffeb;
         4'h3e98 	:	val_out <= 4'hffec;
         4'h3e99 	:	val_out <= 4'hffec;
         4'h3e9a 	:	val_out <= 4'hffec;
         4'h3e9b 	:	val_out <= 4'hffec;
         4'h3ea0 	:	val_out <= 4'hffed;
         4'h3ea1 	:	val_out <= 4'hffed;
         4'h3ea2 	:	val_out <= 4'hffed;
         4'h3ea3 	:	val_out <= 4'hffed;
         4'h3ea8 	:	val_out <= 4'hffee;
         4'h3ea9 	:	val_out <= 4'hffee;
         4'h3eaa 	:	val_out <= 4'hffee;
         4'h3eab 	:	val_out <= 4'hffee;
         4'h3eb0 	:	val_out <= 4'hffee;
         4'h3eb1 	:	val_out <= 4'hffee;
         4'h3eb2 	:	val_out <= 4'hffee;
         4'h3eb3 	:	val_out <= 4'hffee;
         4'h3eb8 	:	val_out <= 4'hffef;
         4'h3eb9 	:	val_out <= 4'hffef;
         4'h3eba 	:	val_out <= 4'hffef;
         4'h3ebb 	:	val_out <= 4'hffef;
         4'h3ec0 	:	val_out <= 4'hfff0;
         4'h3ec1 	:	val_out <= 4'hfff0;
         4'h3ec2 	:	val_out <= 4'hfff0;
         4'h3ec3 	:	val_out <= 4'hfff0;
         4'h3ec8 	:	val_out <= 4'hfff1;
         4'h3ec9 	:	val_out <= 4'hfff1;
         4'h3eca 	:	val_out <= 4'hfff1;
         4'h3ecb 	:	val_out <= 4'hfff1;
         4'h3ed0 	:	val_out <= 4'hfff2;
         4'h3ed1 	:	val_out <= 4'hfff2;
         4'h3ed2 	:	val_out <= 4'hfff2;
         4'h3ed3 	:	val_out <= 4'hfff2;
         4'h3ed8 	:	val_out <= 4'hfff2;
         4'h3ed9 	:	val_out <= 4'hfff2;
         4'h3eda 	:	val_out <= 4'hfff2;
         4'h3edb 	:	val_out <= 4'hfff2;
         4'h3ee0 	:	val_out <= 4'hfff3;
         4'h3ee1 	:	val_out <= 4'hfff3;
         4'h3ee2 	:	val_out <= 4'hfff3;
         4'h3ee3 	:	val_out <= 4'hfff3;
         4'h3ee8 	:	val_out <= 4'hfff4;
         4'h3ee9 	:	val_out <= 4'hfff4;
         4'h3eea 	:	val_out <= 4'hfff4;
         4'h3eeb 	:	val_out <= 4'hfff4;
         4'h3ef0 	:	val_out <= 4'hfff4;
         4'h3ef1 	:	val_out <= 4'hfff4;
         4'h3ef2 	:	val_out <= 4'hfff4;
         4'h3ef3 	:	val_out <= 4'hfff4;
         4'h3ef8 	:	val_out <= 4'hfff5;
         4'h3ef9 	:	val_out <= 4'hfff5;
         4'h3efa 	:	val_out <= 4'hfff5;
         4'h3efb 	:	val_out <= 4'hfff5;
         4'h3f00 	:	val_out <= 4'hfff6;
         4'h3f01 	:	val_out <= 4'hfff6;
         4'h3f02 	:	val_out <= 4'hfff6;
         4'h3f03 	:	val_out <= 4'hfff6;
         4'h3f08 	:	val_out <= 4'hfff6;
         4'h3f09 	:	val_out <= 4'hfff6;
         4'h3f0a 	:	val_out <= 4'hfff6;
         4'h3f0b 	:	val_out <= 4'hfff6;
         4'h3f10 	:	val_out <= 4'hfff7;
         4'h3f11 	:	val_out <= 4'hfff7;
         4'h3f12 	:	val_out <= 4'hfff7;
         4'h3f13 	:	val_out <= 4'hfff7;
         4'h3f18 	:	val_out <= 4'hfff7;
         4'h3f19 	:	val_out <= 4'hfff7;
         4'h3f1a 	:	val_out <= 4'hfff7;
         4'h3f1b 	:	val_out <= 4'hfff7;
         4'h3f20 	:	val_out <= 4'hfff8;
         4'h3f21 	:	val_out <= 4'hfff8;
         4'h3f22 	:	val_out <= 4'hfff8;
         4'h3f23 	:	val_out <= 4'hfff8;
         4'h3f28 	:	val_out <= 4'hfff8;
         4'h3f29 	:	val_out <= 4'hfff8;
         4'h3f2a 	:	val_out <= 4'hfff8;
         4'h3f2b 	:	val_out <= 4'hfff8;
         4'h3f30 	:	val_out <= 4'hfff9;
         4'h3f31 	:	val_out <= 4'hfff9;
         4'h3f32 	:	val_out <= 4'hfff9;
         4'h3f33 	:	val_out <= 4'hfff9;
         4'h3f38 	:	val_out <= 4'hfff9;
         4'h3f39 	:	val_out <= 4'hfff9;
         4'h3f3a 	:	val_out <= 4'hfff9;
         4'h3f3b 	:	val_out <= 4'hfff9;
         4'h3f40 	:	val_out <= 4'hfffa;
         4'h3f41 	:	val_out <= 4'hfffa;
         4'h3f42 	:	val_out <= 4'hfffa;
         4'h3f43 	:	val_out <= 4'hfffa;
         4'h3f48 	:	val_out <= 4'hfffa;
         4'h3f49 	:	val_out <= 4'hfffa;
         4'h3f4a 	:	val_out <= 4'hfffa;
         4'h3f4b 	:	val_out <= 4'hfffa;
         4'h3f50 	:	val_out <= 4'hfffb;
         4'h3f51 	:	val_out <= 4'hfffb;
         4'h3f52 	:	val_out <= 4'hfffb;
         4'h3f53 	:	val_out <= 4'hfffb;
         4'h3f58 	:	val_out <= 4'hfffb;
         4'h3f59 	:	val_out <= 4'hfffb;
         4'h3f5a 	:	val_out <= 4'hfffb;
         4'h3f5b 	:	val_out <= 4'hfffb;
         4'h3f60 	:	val_out <= 4'hfffc;
         4'h3f61 	:	val_out <= 4'hfffc;
         4'h3f62 	:	val_out <= 4'hfffc;
         4'h3f63 	:	val_out <= 4'hfffc;
         4'h3f68 	:	val_out <= 4'hfffc;
         4'h3f69 	:	val_out <= 4'hfffc;
         4'h3f6a 	:	val_out <= 4'hfffc;
         4'h3f6b 	:	val_out <= 4'hfffc;
         4'h3f70 	:	val_out <= 4'hfffc;
         4'h3f71 	:	val_out <= 4'hfffc;
         4'h3f72 	:	val_out <= 4'hfffc;
         4'h3f73 	:	val_out <= 4'hfffc;
         4'h3f78 	:	val_out <= 4'hfffd;
         4'h3f79 	:	val_out <= 4'hfffd;
         4'h3f7a 	:	val_out <= 4'hfffd;
         4'h3f7b 	:	val_out <= 4'hfffd;
         4'h3f80 	:	val_out <= 4'hfffd;
         4'h3f81 	:	val_out <= 4'hfffd;
         4'h3f82 	:	val_out <= 4'hfffd;
         4'h3f83 	:	val_out <= 4'hfffd;
         4'h3f88 	:	val_out <= 4'hfffd;
         4'h3f89 	:	val_out <= 4'hfffd;
         4'h3f8a 	:	val_out <= 4'hfffd;
         4'h3f8b 	:	val_out <= 4'hfffd;
         4'h3f90 	:	val_out <= 4'hfffe;
         4'h3f91 	:	val_out <= 4'hfffe;
         4'h3f92 	:	val_out <= 4'hfffe;
         4'h3f93 	:	val_out <= 4'hfffe;
         4'h3f98 	:	val_out <= 4'hfffe;
         4'h3f99 	:	val_out <= 4'hfffe;
         4'h3f9a 	:	val_out <= 4'hfffe;
         4'h3f9b 	:	val_out <= 4'hfffe;
         4'h3fa0 	:	val_out <= 4'hfffe;
         4'h3fa1 	:	val_out <= 4'hfffe;
         4'h3fa2 	:	val_out <= 4'hfffe;
         4'h3fa3 	:	val_out <= 4'hfffe;
         4'h3fa8 	:	val_out <= 4'hfffe;
         4'h3fa9 	:	val_out <= 4'hfffe;
         4'h3faa 	:	val_out <= 4'hfffe;
         4'h3fab 	:	val_out <= 4'hfffe;
         4'h3fb0 	:	val_out <= 4'hffff;
         4'h3fb1 	:	val_out <= 4'hffff;
         4'h3fb2 	:	val_out <= 4'hffff;
         4'h3fb3 	:	val_out <= 4'hffff;
         4'h3fb8 	:	val_out <= 4'hffff;
         4'h3fb9 	:	val_out <= 4'hffff;
         4'h3fba 	:	val_out <= 4'hffff;
         4'h3fbb 	:	val_out <= 4'hffff;
         4'h3fc0 	:	val_out <= 4'hffff;
         4'h3fc1 	:	val_out <= 4'hffff;
         4'h3fc2 	:	val_out <= 4'hffff;
         4'h3fc3 	:	val_out <= 4'hffff;
         4'h3fc8 	:	val_out <= 4'hffff;
         4'h3fc9 	:	val_out <= 4'hffff;
         4'h3fca 	:	val_out <= 4'hffff;
         4'h3fcb 	:	val_out <= 4'hffff;
         4'h3fd0 	:	val_out <= 4'hffff;
         4'h3fd1 	:	val_out <= 4'hffff;
         4'h3fd2 	:	val_out <= 4'hffff;
         4'h3fd3 	:	val_out <= 4'hffff;
         4'h3fd8 	:	val_out <= 4'hffff;
         4'h3fd9 	:	val_out <= 4'hffff;
         4'h3fda 	:	val_out <= 4'hffff;
         4'h3fdb 	:	val_out <= 4'hffff;
         4'h3fe0 	:	val_out <= 4'hffff;
         4'h3fe1 	:	val_out <= 4'hffff;
         4'h3fe2 	:	val_out <= 4'hffff;
         4'h3fe3 	:	val_out <= 4'hffff;
         4'h3fe8 	:	val_out <= 4'hffff;
         4'h3fe9 	:	val_out <= 4'hffff;
         4'h3fea 	:	val_out <= 4'hffff;
         4'h3feb 	:	val_out <= 4'hffff;
         4'h3ff0 	:	val_out <= 4'hffff;
         4'h3ff1 	:	val_out <= 4'hffff;
         4'h3ff2 	:	val_out <= 4'hffff;
         4'h3ff3 	:	val_out <= 4'hffff;
         4'h3ff8 	:	val_out <= 4'hffff;
         4'h3ff9 	:	val_out <= 4'hffff;
         4'h3ffa 	:	val_out <= 4'hffff;
         4'h3ffb 	:	val_out <= 4'hffff;
         4'h4000 	:	val_out <= 4'h10000;
         4'h4001 	:	val_out <= 4'h10000;
         4'h4002 	:	val_out <= 4'h10000;
         4'h4003 	:	val_out <= 4'h10000;
         4'h4008 	:	val_out <= 4'hffff;
         4'h4009 	:	val_out <= 4'hffff;
         4'h400a 	:	val_out <= 4'hffff;
         4'h400b 	:	val_out <= 4'hffff;
         4'h4010 	:	val_out <= 4'hffff;
         4'h4011 	:	val_out <= 4'hffff;
         4'h4012 	:	val_out <= 4'hffff;
         4'h4013 	:	val_out <= 4'hffff;
         4'h4018 	:	val_out <= 4'hffff;
         4'h4019 	:	val_out <= 4'hffff;
         4'h401a 	:	val_out <= 4'hffff;
         4'h401b 	:	val_out <= 4'hffff;
         4'h4020 	:	val_out <= 4'hffff;
         4'h4021 	:	val_out <= 4'hffff;
         4'h4022 	:	val_out <= 4'hffff;
         4'h4023 	:	val_out <= 4'hffff;
         4'h4028 	:	val_out <= 4'hffff;
         4'h4029 	:	val_out <= 4'hffff;
         4'h402a 	:	val_out <= 4'hffff;
         4'h402b 	:	val_out <= 4'hffff;
         4'h4030 	:	val_out <= 4'hffff;
         4'h4031 	:	val_out <= 4'hffff;
         4'h4032 	:	val_out <= 4'hffff;
         4'h4033 	:	val_out <= 4'hffff;
         4'h4038 	:	val_out <= 4'hffff;
         4'h4039 	:	val_out <= 4'hffff;
         4'h403a 	:	val_out <= 4'hffff;
         4'h403b 	:	val_out <= 4'hffff;
         4'h4040 	:	val_out <= 4'hffff;
         4'h4041 	:	val_out <= 4'hffff;
         4'h4042 	:	val_out <= 4'hffff;
         4'h4043 	:	val_out <= 4'hffff;
         4'h4048 	:	val_out <= 4'hffff;
         4'h4049 	:	val_out <= 4'hffff;
         4'h404a 	:	val_out <= 4'hffff;
         4'h404b 	:	val_out <= 4'hffff;
         4'h4050 	:	val_out <= 4'hffff;
         4'h4051 	:	val_out <= 4'hffff;
         4'h4052 	:	val_out <= 4'hffff;
         4'h4053 	:	val_out <= 4'hffff;
         4'h4058 	:	val_out <= 4'hfffe;
         4'h4059 	:	val_out <= 4'hfffe;
         4'h405a 	:	val_out <= 4'hfffe;
         4'h405b 	:	val_out <= 4'hfffe;
         4'h4060 	:	val_out <= 4'hfffe;
         4'h4061 	:	val_out <= 4'hfffe;
         4'h4062 	:	val_out <= 4'hfffe;
         4'h4063 	:	val_out <= 4'hfffe;
         4'h4068 	:	val_out <= 4'hfffe;
         4'h4069 	:	val_out <= 4'hfffe;
         4'h406a 	:	val_out <= 4'hfffe;
         4'h406b 	:	val_out <= 4'hfffe;
         4'h4070 	:	val_out <= 4'hfffe;
         4'h4071 	:	val_out <= 4'hfffe;
         4'h4072 	:	val_out <= 4'hfffe;
         4'h4073 	:	val_out <= 4'hfffe;
         4'h4078 	:	val_out <= 4'hfffd;
         4'h4079 	:	val_out <= 4'hfffd;
         4'h407a 	:	val_out <= 4'hfffd;
         4'h407b 	:	val_out <= 4'hfffd;
         4'h4080 	:	val_out <= 4'hfffd;
         4'h4081 	:	val_out <= 4'hfffd;
         4'h4082 	:	val_out <= 4'hfffd;
         4'h4083 	:	val_out <= 4'hfffd;
         4'h4088 	:	val_out <= 4'hfffd;
         4'h4089 	:	val_out <= 4'hfffd;
         4'h408a 	:	val_out <= 4'hfffd;
         4'h408b 	:	val_out <= 4'hfffd;
         4'h4090 	:	val_out <= 4'hfffc;
         4'h4091 	:	val_out <= 4'hfffc;
         4'h4092 	:	val_out <= 4'hfffc;
         4'h4093 	:	val_out <= 4'hfffc;
         4'h4098 	:	val_out <= 4'hfffc;
         4'h4099 	:	val_out <= 4'hfffc;
         4'h409a 	:	val_out <= 4'hfffc;
         4'h409b 	:	val_out <= 4'hfffc;
         4'h40a0 	:	val_out <= 4'hfffc;
         4'h40a1 	:	val_out <= 4'hfffc;
         4'h40a2 	:	val_out <= 4'hfffc;
         4'h40a3 	:	val_out <= 4'hfffc;
         4'h40a8 	:	val_out <= 4'hfffb;
         4'h40a9 	:	val_out <= 4'hfffb;
         4'h40aa 	:	val_out <= 4'hfffb;
         4'h40ab 	:	val_out <= 4'hfffb;
         4'h40b0 	:	val_out <= 4'hfffb;
         4'h40b1 	:	val_out <= 4'hfffb;
         4'h40b2 	:	val_out <= 4'hfffb;
         4'h40b3 	:	val_out <= 4'hfffb;
         4'h40b8 	:	val_out <= 4'hfffa;
         4'h40b9 	:	val_out <= 4'hfffa;
         4'h40ba 	:	val_out <= 4'hfffa;
         4'h40bb 	:	val_out <= 4'hfffa;
         4'h40c0 	:	val_out <= 4'hfffa;
         4'h40c1 	:	val_out <= 4'hfffa;
         4'h40c2 	:	val_out <= 4'hfffa;
         4'h40c3 	:	val_out <= 4'hfffa;
         4'h40c8 	:	val_out <= 4'hfff9;
         4'h40c9 	:	val_out <= 4'hfff9;
         4'h40ca 	:	val_out <= 4'hfff9;
         4'h40cb 	:	val_out <= 4'hfff9;
         4'h40d0 	:	val_out <= 4'hfff9;
         4'h40d1 	:	val_out <= 4'hfff9;
         4'h40d2 	:	val_out <= 4'hfff9;
         4'h40d3 	:	val_out <= 4'hfff9;
         4'h40d8 	:	val_out <= 4'hfff8;
         4'h40d9 	:	val_out <= 4'hfff8;
         4'h40da 	:	val_out <= 4'hfff8;
         4'h40db 	:	val_out <= 4'hfff8;
         4'h40e0 	:	val_out <= 4'hfff8;
         4'h40e1 	:	val_out <= 4'hfff8;
         4'h40e2 	:	val_out <= 4'hfff8;
         4'h40e3 	:	val_out <= 4'hfff8;
         4'h40e8 	:	val_out <= 4'hfff7;
         4'h40e9 	:	val_out <= 4'hfff7;
         4'h40ea 	:	val_out <= 4'hfff7;
         4'h40eb 	:	val_out <= 4'hfff7;
         4'h40f0 	:	val_out <= 4'hfff7;
         4'h40f1 	:	val_out <= 4'hfff7;
         4'h40f2 	:	val_out <= 4'hfff7;
         4'h40f3 	:	val_out <= 4'hfff7;
         4'h40f8 	:	val_out <= 4'hfff6;
         4'h40f9 	:	val_out <= 4'hfff6;
         4'h40fa 	:	val_out <= 4'hfff6;
         4'h40fb 	:	val_out <= 4'hfff6;
         4'h4100 	:	val_out <= 4'hfff6;
         4'h4101 	:	val_out <= 4'hfff6;
         4'h4102 	:	val_out <= 4'hfff6;
         4'h4103 	:	val_out <= 4'hfff6;
         4'h4108 	:	val_out <= 4'hfff5;
         4'h4109 	:	val_out <= 4'hfff5;
         4'h410a 	:	val_out <= 4'hfff5;
         4'h410b 	:	val_out <= 4'hfff5;
         4'h4110 	:	val_out <= 4'hfff4;
         4'h4111 	:	val_out <= 4'hfff4;
         4'h4112 	:	val_out <= 4'hfff4;
         4'h4113 	:	val_out <= 4'hfff4;
         4'h4118 	:	val_out <= 4'hfff4;
         4'h4119 	:	val_out <= 4'hfff4;
         4'h411a 	:	val_out <= 4'hfff4;
         4'h411b 	:	val_out <= 4'hfff4;
         4'h4120 	:	val_out <= 4'hfff3;
         4'h4121 	:	val_out <= 4'hfff3;
         4'h4122 	:	val_out <= 4'hfff3;
         4'h4123 	:	val_out <= 4'hfff3;
         4'h4128 	:	val_out <= 4'hfff2;
         4'h4129 	:	val_out <= 4'hfff2;
         4'h412a 	:	val_out <= 4'hfff2;
         4'h412b 	:	val_out <= 4'hfff2;
         4'h4130 	:	val_out <= 4'hfff2;
         4'h4131 	:	val_out <= 4'hfff2;
         4'h4132 	:	val_out <= 4'hfff2;
         4'h4133 	:	val_out <= 4'hfff2;
         4'h4138 	:	val_out <= 4'hfff1;
         4'h4139 	:	val_out <= 4'hfff1;
         4'h413a 	:	val_out <= 4'hfff1;
         4'h413b 	:	val_out <= 4'hfff1;
         4'h4140 	:	val_out <= 4'hfff0;
         4'h4141 	:	val_out <= 4'hfff0;
         4'h4142 	:	val_out <= 4'hfff0;
         4'h4143 	:	val_out <= 4'hfff0;
         4'h4148 	:	val_out <= 4'hffef;
         4'h4149 	:	val_out <= 4'hffef;
         4'h414a 	:	val_out <= 4'hffef;
         4'h414b 	:	val_out <= 4'hffef;
         4'h4150 	:	val_out <= 4'hffee;
         4'h4151 	:	val_out <= 4'hffee;
         4'h4152 	:	val_out <= 4'hffee;
         4'h4153 	:	val_out <= 4'hffee;
         4'h4158 	:	val_out <= 4'hffee;
         4'h4159 	:	val_out <= 4'hffee;
         4'h415a 	:	val_out <= 4'hffee;
         4'h415b 	:	val_out <= 4'hffee;
         4'h4160 	:	val_out <= 4'hffed;
         4'h4161 	:	val_out <= 4'hffed;
         4'h4162 	:	val_out <= 4'hffed;
         4'h4163 	:	val_out <= 4'hffed;
         4'h4168 	:	val_out <= 4'hffec;
         4'h4169 	:	val_out <= 4'hffec;
         4'h416a 	:	val_out <= 4'hffec;
         4'h416b 	:	val_out <= 4'hffec;
         4'h4170 	:	val_out <= 4'hffeb;
         4'h4171 	:	val_out <= 4'hffeb;
         4'h4172 	:	val_out <= 4'hffeb;
         4'h4173 	:	val_out <= 4'hffeb;
         4'h4178 	:	val_out <= 4'hffea;
         4'h4179 	:	val_out <= 4'hffea;
         4'h417a 	:	val_out <= 4'hffea;
         4'h417b 	:	val_out <= 4'hffea;
         4'h4180 	:	val_out <= 4'hffe9;
         4'h4181 	:	val_out <= 4'hffe9;
         4'h4182 	:	val_out <= 4'hffe9;
         4'h4183 	:	val_out <= 4'hffe9;
         4'h4188 	:	val_out <= 4'hffe8;
         4'h4189 	:	val_out <= 4'hffe8;
         4'h418a 	:	val_out <= 4'hffe8;
         4'h418b 	:	val_out <= 4'hffe8;
         4'h4190 	:	val_out <= 4'hffe7;
         4'h4191 	:	val_out <= 4'hffe7;
         4'h4192 	:	val_out <= 4'hffe7;
         4'h4193 	:	val_out <= 4'hffe7;
         4'h4198 	:	val_out <= 4'hffe6;
         4'h4199 	:	val_out <= 4'hffe6;
         4'h419a 	:	val_out <= 4'hffe6;
         4'h419b 	:	val_out <= 4'hffe6;
         4'h41a0 	:	val_out <= 4'hffe5;
         4'h41a1 	:	val_out <= 4'hffe5;
         4'h41a2 	:	val_out <= 4'hffe5;
         4'h41a3 	:	val_out <= 4'hffe5;
         4'h41a8 	:	val_out <= 4'hffe4;
         4'h41a9 	:	val_out <= 4'hffe4;
         4'h41aa 	:	val_out <= 4'hffe4;
         4'h41ab 	:	val_out <= 4'hffe4;
         4'h41b0 	:	val_out <= 4'hffe3;
         4'h41b1 	:	val_out <= 4'hffe3;
         4'h41b2 	:	val_out <= 4'hffe3;
         4'h41b3 	:	val_out <= 4'hffe3;
         4'h41b8 	:	val_out <= 4'hffe2;
         4'h41b9 	:	val_out <= 4'hffe2;
         4'h41ba 	:	val_out <= 4'hffe2;
         4'h41bb 	:	val_out <= 4'hffe2;
         4'h41c0 	:	val_out <= 4'hffe1;
         4'h41c1 	:	val_out <= 4'hffe1;
         4'h41c2 	:	val_out <= 4'hffe1;
         4'h41c3 	:	val_out <= 4'hffe1;
         4'h41c8 	:	val_out <= 4'hffe0;
         4'h41c9 	:	val_out <= 4'hffe0;
         4'h41ca 	:	val_out <= 4'hffe0;
         4'h41cb 	:	val_out <= 4'hffe0;
         4'h41d0 	:	val_out <= 4'hffdf;
         4'h41d1 	:	val_out <= 4'hffdf;
         4'h41d2 	:	val_out <= 4'hffdf;
         4'h41d3 	:	val_out <= 4'hffdf;
         4'h41d8 	:	val_out <= 4'hffde;
         4'h41d9 	:	val_out <= 4'hffde;
         4'h41da 	:	val_out <= 4'hffde;
         4'h41db 	:	val_out <= 4'hffde;
         4'h41e0 	:	val_out <= 4'hffdd;
         4'h41e1 	:	val_out <= 4'hffdd;
         4'h41e2 	:	val_out <= 4'hffdd;
         4'h41e3 	:	val_out <= 4'hffdd;
         4'h41e8 	:	val_out <= 4'hffdc;
         4'h41e9 	:	val_out <= 4'hffdc;
         4'h41ea 	:	val_out <= 4'hffdc;
         4'h41eb 	:	val_out <= 4'hffdc;
         4'h41f0 	:	val_out <= 4'hffda;
         4'h41f1 	:	val_out <= 4'hffda;
         4'h41f2 	:	val_out <= 4'hffda;
         4'h41f3 	:	val_out <= 4'hffda;
         4'h41f8 	:	val_out <= 4'hffd9;
         4'h41f9 	:	val_out <= 4'hffd9;
         4'h41fa 	:	val_out <= 4'hffd9;
         4'h41fb 	:	val_out <= 4'hffd9;
         4'h4200 	:	val_out <= 4'hffd8;
         4'h4201 	:	val_out <= 4'hffd8;
         4'h4202 	:	val_out <= 4'hffd8;
         4'h4203 	:	val_out <= 4'hffd8;
         4'h4208 	:	val_out <= 4'hffd7;
         4'h4209 	:	val_out <= 4'hffd7;
         4'h420a 	:	val_out <= 4'hffd7;
         4'h420b 	:	val_out <= 4'hffd7;
         4'h4210 	:	val_out <= 4'hffd6;
         4'h4211 	:	val_out <= 4'hffd6;
         4'h4212 	:	val_out <= 4'hffd6;
         4'h4213 	:	val_out <= 4'hffd6;
         4'h4218 	:	val_out <= 4'hffd4;
         4'h4219 	:	val_out <= 4'hffd4;
         4'h421a 	:	val_out <= 4'hffd4;
         4'h421b 	:	val_out <= 4'hffd4;
         4'h4220 	:	val_out <= 4'hffd3;
         4'h4221 	:	val_out <= 4'hffd3;
         4'h4222 	:	val_out <= 4'hffd3;
         4'h4223 	:	val_out <= 4'hffd3;
         4'h4228 	:	val_out <= 4'hffd2;
         4'h4229 	:	val_out <= 4'hffd2;
         4'h422a 	:	val_out <= 4'hffd2;
         4'h422b 	:	val_out <= 4'hffd2;
         4'h4230 	:	val_out <= 4'hffd0;
         4'h4231 	:	val_out <= 4'hffd0;
         4'h4232 	:	val_out <= 4'hffd0;
         4'h4233 	:	val_out <= 4'hffd0;
         4'h4238 	:	val_out <= 4'hffcf;
         4'h4239 	:	val_out <= 4'hffcf;
         4'h423a 	:	val_out <= 4'hffcf;
         4'h423b 	:	val_out <= 4'hffcf;
         4'h4240 	:	val_out <= 4'hffce;
         4'h4241 	:	val_out <= 4'hffce;
         4'h4242 	:	val_out <= 4'hffce;
         4'h4243 	:	val_out <= 4'hffce;
         4'h4248 	:	val_out <= 4'hffcc;
         4'h4249 	:	val_out <= 4'hffcc;
         4'h424a 	:	val_out <= 4'hffcc;
         4'h424b 	:	val_out <= 4'hffcc;
         4'h4250 	:	val_out <= 4'hffcb;
         4'h4251 	:	val_out <= 4'hffcb;
         4'h4252 	:	val_out <= 4'hffcb;
         4'h4253 	:	val_out <= 4'hffcb;
         4'h4258 	:	val_out <= 4'hffc9;
         4'h4259 	:	val_out <= 4'hffc9;
         4'h425a 	:	val_out <= 4'hffc9;
         4'h425b 	:	val_out <= 4'hffc9;
         4'h4260 	:	val_out <= 4'hffc8;
         4'h4261 	:	val_out <= 4'hffc8;
         4'h4262 	:	val_out <= 4'hffc8;
         4'h4263 	:	val_out <= 4'hffc8;
         4'h4268 	:	val_out <= 4'hffc6;
         4'h4269 	:	val_out <= 4'hffc6;
         4'h426a 	:	val_out <= 4'hffc6;
         4'h426b 	:	val_out <= 4'hffc6;
         4'h4270 	:	val_out <= 4'hffc5;
         4'h4271 	:	val_out <= 4'hffc5;
         4'h4272 	:	val_out <= 4'hffc5;
         4'h4273 	:	val_out <= 4'hffc5;
         4'h4278 	:	val_out <= 4'hffc3;
         4'h4279 	:	val_out <= 4'hffc3;
         4'h427a 	:	val_out <= 4'hffc3;
         4'h427b 	:	val_out <= 4'hffc3;
         4'h4280 	:	val_out <= 4'hffc2;
         4'h4281 	:	val_out <= 4'hffc2;
         4'h4282 	:	val_out <= 4'hffc2;
         4'h4283 	:	val_out <= 4'hffc2;
         4'h4288 	:	val_out <= 4'hffc0;
         4'h4289 	:	val_out <= 4'hffc0;
         4'h428a 	:	val_out <= 4'hffc0;
         4'h428b 	:	val_out <= 4'hffc0;
         4'h4290 	:	val_out <= 4'hffbf;
         4'h4291 	:	val_out <= 4'hffbf;
         4'h4292 	:	val_out <= 4'hffbf;
         4'h4293 	:	val_out <= 4'hffbf;
         4'h4298 	:	val_out <= 4'hffbd;
         4'h4299 	:	val_out <= 4'hffbd;
         4'h429a 	:	val_out <= 4'hffbd;
         4'h429b 	:	val_out <= 4'hffbd;
         4'h42a0 	:	val_out <= 4'hffbc;
         4'h42a1 	:	val_out <= 4'hffbc;
         4'h42a2 	:	val_out <= 4'hffbc;
         4'h42a3 	:	val_out <= 4'hffbc;
         4'h42a8 	:	val_out <= 4'hffba;
         4'h42a9 	:	val_out <= 4'hffba;
         4'h42aa 	:	val_out <= 4'hffba;
         4'h42ab 	:	val_out <= 4'hffba;
         4'h42b0 	:	val_out <= 4'hffb8;
         4'h42b1 	:	val_out <= 4'hffb8;
         4'h42b2 	:	val_out <= 4'hffb8;
         4'h42b3 	:	val_out <= 4'hffb8;
         4'h42b8 	:	val_out <= 4'hffb7;
         4'h42b9 	:	val_out <= 4'hffb7;
         4'h42ba 	:	val_out <= 4'hffb7;
         4'h42bb 	:	val_out <= 4'hffb7;
         4'h42c0 	:	val_out <= 4'hffb5;
         4'h42c1 	:	val_out <= 4'hffb5;
         4'h42c2 	:	val_out <= 4'hffb5;
         4'h42c3 	:	val_out <= 4'hffb5;
         4'h42c8 	:	val_out <= 4'hffb3;
         4'h42c9 	:	val_out <= 4'hffb3;
         4'h42ca 	:	val_out <= 4'hffb3;
         4'h42cb 	:	val_out <= 4'hffb3;
         4'h42d0 	:	val_out <= 4'hffb1;
         4'h42d1 	:	val_out <= 4'hffb1;
         4'h42d2 	:	val_out <= 4'hffb1;
         4'h42d3 	:	val_out <= 4'hffb1;
         4'h42d8 	:	val_out <= 4'hffb0;
         4'h42d9 	:	val_out <= 4'hffb0;
         4'h42da 	:	val_out <= 4'hffb0;
         4'h42db 	:	val_out <= 4'hffb0;
         4'h42e0 	:	val_out <= 4'hffae;
         4'h42e1 	:	val_out <= 4'hffae;
         4'h42e2 	:	val_out <= 4'hffae;
         4'h42e3 	:	val_out <= 4'hffae;
         4'h42e8 	:	val_out <= 4'hffac;
         4'h42e9 	:	val_out <= 4'hffac;
         4'h42ea 	:	val_out <= 4'hffac;
         4'h42eb 	:	val_out <= 4'hffac;
         4'h42f0 	:	val_out <= 4'hffaa;
         4'h42f1 	:	val_out <= 4'hffaa;
         4'h42f2 	:	val_out <= 4'hffaa;
         4'h42f3 	:	val_out <= 4'hffaa;
         4'h42f8 	:	val_out <= 4'hffa9;
         4'h42f9 	:	val_out <= 4'hffa9;
         4'h42fa 	:	val_out <= 4'hffa9;
         4'h42fb 	:	val_out <= 4'hffa9;
         4'h4300 	:	val_out <= 4'hffa7;
         4'h4301 	:	val_out <= 4'hffa7;
         4'h4302 	:	val_out <= 4'hffa7;
         4'h4303 	:	val_out <= 4'hffa7;
         4'h4308 	:	val_out <= 4'hffa5;
         4'h4309 	:	val_out <= 4'hffa5;
         4'h430a 	:	val_out <= 4'hffa5;
         4'h430b 	:	val_out <= 4'hffa5;
         4'h4310 	:	val_out <= 4'hffa3;
         4'h4311 	:	val_out <= 4'hffa3;
         4'h4312 	:	val_out <= 4'hffa3;
         4'h4313 	:	val_out <= 4'hffa3;
         4'h4318 	:	val_out <= 4'hffa1;
         4'h4319 	:	val_out <= 4'hffa1;
         4'h431a 	:	val_out <= 4'hffa1;
         4'h431b 	:	val_out <= 4'hffa1;
         4'h4320 	:	val_out <= 4'hff9f;
         4'h4321 	:	val_out <= 4'hff9f;
         4'h4322 	:	val_out <= 4'hff9f;
         4'h4323 	:	val_out <= 4'hff9f;
         4'h4328 	:	val_out <= 4'hff9d;
         4'h4329 	:	val_out <= 4'hff9d;
         4'h432a 	:	val_out <= 4'hff9d;
         4'h432b 	:	val_out <= 4'hff9d;
         4'h4330 	:	val_out <= 4'hff9b;
         4'h4331 	:	val_out <= 4'hff9b;
         4'h4332 	:	val_out <= 4'hff9b;
         4'h4333 	:	val_out <= 4'hff9b;
         4'h4338 	:	val_out <= 4'hff99;
         4'h4339 	:	val_out <= 4'hff99;
         4'h433a 	:	val_out <= 4'hff99;
         4'h433b 	:	val_out <= 4'hff99;
         4'h4340 	:	val_out <= 4'hff97;
         4'h4341 	:	val_out <= 4'hff97;
         4'h4342 	:	val_out <= 4'hff97;
         4'h4343 	:	val_out <= 4'hff97;
         4'h4348 	:	val_out <= 4'hff95;
         4'h4349 	:	val_out <= 4'hff95;
         4'h434a 	:	val_out <= 4'hff95;
         4'h434b 	:	val_out <= 4'hff95;
         4'h4350 	:	val_out <= 4'hff93;
         4'h4351 	:	val_out <= 4'hff93;
         4'h4352 	:	val_out <= 4'hff93;
         4'h4353 	:	val_out <= 4'hff93;
         4'h4358 	:	val_out <= 4'hff91;
         4'h4359 	:	val_out <= 4'hff91;
         4'h435a 	:	val_out <= 4'hff91;
         4'h435b 	:	val_out <= 4'hff91;
         4'h4360 	:	val_out <= 4'hff8f;
         4'h4361 	:	val_out <= 4'hff8f;
         4'h4362 	:	val_out <= 4'hff8f;
         4'h4363 	:	val_out <= 4'hff8f;
         4'h4368 	:	val_out <= 4'hff8d;
         4'h4369 	:	val_out <= 4'hff8d;
         4'h436a 	:	val_out <= 4'hff8d;
         4'h436b 	:	val_out <= 4'hff8d;
         4'h4370 	:	val_out <= 4'hff8b;
         4'h4371 	:	val_out <= 4'hff8b;
         4'h4372 	:	val_out <= 4'hff8b;
         4'h4373 	:	val_out <= 4'hff8b;
         4'h4378 	:	val_out <= 4'hff89;
         4'h4379 	:	val_out <= 4'hff89;
         4'h437a 	:	val_out <= 4'hff89;
         4'h437b 	:	val_out <= 4'hff89;
         4'h4380 	:	val_out <= 4'hff87;
         4'h4381 	:	val_out <= 4'hff87;
         4'h4382 	:	val_out <= 4'hff87;
         4'h4383 	:	val_out <= 4'hff87;
         4'h4388 	:	val_out <= 4'hff85;
         4'h4389 	:	val_out <= 4'hff85;
         4'h438a 	:	val_out <= 4'hff85;
         4'h438b 	:	val_out <= 4'hff85;
         4'h4390 	:	val_out <= 4'hff82;
         4'h4391 	:	val_out <= 4'hff82;
         4'h4392 	:	val_out <= 4'hff82;
         4'h4393 	:	val_out <= 4'hff82;
         4'h4398 	:	val_out <= 4'hff80;
         4'h4399 	:	val_out <= 4'hff80;
         4'h439a 	:	val_out <= 4'hff80;
         4'h439b 	:	val_out <= 4'hff80;
         4'h43a0 	:	val_out <= 4'hff7e;
         4'h43a1 	:	val_out <= 4'hff7e;
         4'h43a2 	:	val_out <= 4'hff7e;
         4'h43a3 	:	val_out <= 4'hff7e;
         4'h43a8 	:	val_out <= 4'hff7c;
         4'h43a9 	:	val_out <= 4'hff7c;
         4'h43aa 	:	val_out <= 4'hff7c;
         4'h43ab 	:	val_out <= 4'hff7c;
         4'h43b0 	:	val_out <= 4'hff79;
         4'h43b1 	:	val_out <= 4'hff79;
         4'h43b2 	:	val_out <= 4'hff79;
         4'h43b3 	:	val_out <= 4'hff79;
         4'h43b8 	:	val_out <= 4'hff77;
         4'h43b9 	:	val_out <= 4'hff77;
         4'h43ba 	:	val_out <= 4'hff77;
         4'h43bb 	:	val_out <= 4'hff77;
         4'h43c0 	:	val_out <= 4'hff75;
         4'h43c1 	:	val_out <= 4'hff75;
         4'h43c2 	:	val_out <= 4'hff75;
         4'h43c3 	:	val_out <= 4'hff75;
         4'h43c8 	:	val_out <= 4'hff72;
         4'h43c9 	:	val_out <= 4'hff72;
         4'h43ca 	:	val_out <= 4'hff72;
         4'h43cb 	:	val_out <= 4'hff72;
         4'h43d0 	:	val_out <= 4'hff70;
         4'h43d1 	:	val_out <= 4'hff70;
         4'h43d2 	:	val_out <= 4'hff70;
         4'h43d3 	:	val_out <= 4'hff70;
         4'h43d8 	:	val_out <= 4'hff6e;
         4'h43d9 	:	val_out <= 4'hff6e;
         4'h43da 	:	val_out <= 4'hff6e;
         4'h43db 	:	val_out <= 4'hff6e;
         4'h43e0 	:	val_out <= 4'hff6b;
         4'h43e1 	:	val_out <= 4'hff6b;
         4'h43e2 	:	val_out <= 4'hff6b;
         4'h43e3 	:	val_out <= 4'hff6b;
         4'h43e8 	:	val_out <= 4'hff69;
         4'h43e9 	:	val_out <= 4'hff69;
         4'h43ea 	:	val_out <= 4'hff69;
         4'h43eb 	:	val_out <= 4'hff69;
         4'h43f0 	:	val_out <= 4'hff67;
         4'h43f1 	:	val_out <= 4'hff67;
         4'h43f2 	:	val_out <= 4'hff67;
         4'h43f3 	:	val_out <= 4'hff67;
         4'h43f8 	:	val_out <= 4'hff64;
         4'h43f9 	:	val_out <= 4'hff64;
         4'h43fa 	:	val_out <= 4'hff64;
         4'h43fb 	:	val_out <= 4'hff64;
         4'h4400 	:	val_out <= 4'hff62;
         4'h4401 	:	val_out <= 4'hff62;
         4'h4402 	:	val_out <= 4'hff62;
         4'h4403 	:	val_out <= 4'hff62;
         4'h4408 	:	val_out <= 4'hff5f;
         4'h4409 	:	val_out <= 4'hff5f;
         4'h440a 	:	val_out <= 4'hff5f;
         4'h440b 	:	val_out <= 4'hff5f;
         4'h4410 	:	val_out <= 4'hff5d;
         4'h4411 	:	val_out <= 4'hff5d;
         4'h4412 	:	val_out <= 4'hff5d;
         4'h4413 	:	val_out <= 4'hff5d;
         4'h4418 	:	val_out <= 4'hff5a;
         4'h4419 	:	val_out <= 4'hff5a;
         4'h441a 	:	val_out <= 4'hff5a;
         4'h441b 	:	val_out <= 4'hff5a;
         4'h4420 	:	val_out <= 4'hff58;
         4'h4421 	:	val_out <= 4'hff58;
         4'h4422 	:	val_out <= 4'hff58;
         4'h4423 	:	val_out <= 4'hff58;
         4'h4428 	:	val_out <= 4'hff55;
         4'h4429 	:	val_out <= 4'hff55;
         4'h442a 	:	val_out <= 4'hff55;
         4'h442b 	:	val_out <= 4'hff55;
         4'h4430 	:	val_out <= 4'hff53;
         4'h4431 	:	val_out <= 4'hff53;
         4'h4432 	:	val_out <= 4'hff53;
         4'h4433 	:	val_out <= 4'hff53;
         4'h4438 	:	val_out <= 4'hff50;
         4'h4439 	:	val_out <= 4'hff50;
         4'h443a 	:	val_out <= 4'hff50;
         4'h443b 	:	val_out <= 4'hff50;
         4'h4440 	:	val_out <= 4'hff4d;
         4'h4441 	:	val_out <= 4'hff4d;
         4'h4442 	:	val_out <= 4'hff4d;
         4'h4443 	:	val_out <= 4'hff4d;
         4'h4448 	:	val_out <= 4'hff4b;
         4'h4449 	:	val_out <= 4'hff4b;
         4'h444a 	:	val_out <= 4'hff4b;
         4'h444b 	:	val_out <= 4'hff4b;
         4'h4450 	:	val_out <= 4'hff48;
         4'h4451 	:	val_out <= 4'hff48;
         4'h4452 	:	val_out <= 4'hff48;
         4'h4453 	:	val_out <= 4'hff48;
         4'h4458 	:	val_out <= 4'hff45;
         4'h4459 	:	val_out <= 4'hff45;
         4'h445a 	:	val_out <= 4'hff45;
         4'h445b 	:	val_out <= 4'hff45;
         4'h4460 	:	val_out <= 4'hff43;
         4'h4461 	:	val_out <= 4'hff43;
         4'h4462 	:	val_out <= 4'hff43;
         4'h4463 	:	val_out <= 4'hff43;
         4'h4468 	:	val_out <= 4'hff40;
         4'h4469 	:	val_out <= 4'hff40;
         4'h446a 	:	val_out <= 4'hff40;
         4'h446b 	:	val_out <= 4'hff40;
         4'h4470 	:	val_out <= 4'hff3d;
         4'h4471 	:	val_out <= 4'hff3d;
         4'h4472 	:	val_out <= 4'hff3d;
         4'h4473 	:	val_out <= 4'hff3d;
         4'h4478 	:	val_out <= 4'hff3b;
         4'h4479 	:	val_out <= 4'hff3b;
         4'h447a 	:	val_out <= 4'hff3b;
         4'h447b 	:	val_out <= 4'hff3b;
         4'h4480 	:	val_out <= 4'hff38;
         4'h4481 	:	val_out <= 4'hff38;
         4'h4482 	:	val_out <= 4'hff38;
         4'h4483 	:	val_out <= 4'hff38;
         4'h4488 	:	val_out <= 4'hff35;
         4'h4489 	:	val_out <= 4'hff35;
         4'h448a 	:	val_out <= 4'hff35;
         4'h448b 	:	val_out <= 4'hff35;
         4'h4490 	:	val_out <= 4'hff32;
         4'h4491 	:	val_out <= 4'hff32;
         4'h4492 	:	val_out <= 4'hff32;
         4'h4493 	:	val_out <= 4'hff32;
         4'h4498 	:	val_out <= 4'hff2f;
         4'h4499 	:	val_out <= 4'hff2f;
         4'h449a 	:	val_out <= 4'hff2f;
         4'h449b 	:	val_out <= 4'hff2f;
         4'h44a0 	:	val_out <= 4'hff2d;
         4'h44a1 	:	val_out <= 4'hff2d;
         4'h44a2 	:	val_out <= 4'hff2d;
         4'h44a3 	:	val_out <= 4'hff2d;
         4'h44a8 	:	val_out <= 4'hff2a;
         4'h44a9 	:	val_out <= 4'hff2a;
         4'h44aa 	:	val_out <= 4'hff2a;
         4'h44ab 	:	val_out <= 4'hff2a;
         4'h44b0 	:	val_out <= 4'hff27;
         4'h44b1 	:	val_out <= 4'hff27;
         4'h44b2 	:	val_out <= 4'hff27;
         4'h44b3 	:	val_out <= 4'hff27;
         4'h44b8 	:	val_out <= 4'hff24;
         4'h44b9 	:	val_out <= 4'hff24;
         4'h44ba 	:	val_out <= 4'hff24;
         4'h44bb 	:	val_out <= 4'hff24;
         4'h44c0 	:	val_out <= 4'hff21;
         4'h44c1 	:	val_out <= 4'hff21;
         4'h44c2 	:	val_out <= 4'hff21;
         4'h44c3 	:	val_out <= 4'hff21;
         4'h44c8 	:	val_out <= 4'hff1e;
         4'h44c9 	:	val_out <= 4'hff1e;
         4'h44ca 	:	val_out <= 4'hff1e;
         4'h44cb 	:	val_out <= 4'hff1e;
         4'h44d0 	:	val_out <= 4'hff1b;
         4'h44d1 	:	val_out <= 4'hff1b;
         4'h44d2 	:	val_out <= 4'hff1b;
         4'h44d3 	:	val_out <= 4'hff1b;
         4'h44d8 	:	val_out <= 4'hff18;
         4'h44d9 	:	val_out <= 4'hff18;
         4'h44da 	:	val_out <= 4'hff18;
         4'h44db 	:	val_out <= 4'hff18;
         4'h44e0 	:	val_out <= 4'hff15;
         4'h44e1 	:	val_out <= 4'hff15;
         4'h44e2 	:	val_out <= 4'hff15;
         4'h44e3 	:	val_out <= 4'hff15;
         4'h44e8 	:	val_out <= 4'hff12;
         4'h44e9 	:	val_out <= 4'hff12;
         4'h44ea 	:	val_out <= 4'hff12;
         4'h44eb 	:	val_out <= 4'hff12;
         4'h44f0 	:	val_out <= 4'hff0f;
         4'h44f1 	:	val_out <= 4'hff0f;
         4'h44f2 	:	val_out <= 4'hff0f;
         4'h44f3 	:	val_out <= 4'hff0f;
         4'h44f8 	:	val_out <= 4'hff0c;
         4'h44f9 	:	val_out <= 4'hff0c;
         4'h44fa 	:	val_out <= 4'hff0c;
         4'h44fb 	:	val_out <= 4'hff0c;
         4'h4500 	:	val_out <= 4'hff09;
         4'h4501 	:	val_out <= 4'hff09;
         4'h4502 	:	val_out <= 4'hff09;
         4'h4503 	:	val_out <= 4'hff09;
         4'h4508 	:	val_out <= 4'hff06;
         4'h4509 	:	val_out <= 4'hff06;
         4'h450a 	:	val_out <= 4'hff06;
         4'h450b 	:	val_out <= 4'hff06;
         4'h4510 	:	val_out <= 4'hff03;
         4'h4511 	:	val_out <= 4'hff03;
         4'h4512 	:	val_out <= 4'hff03;
         4'h4513 	:	val_out <= 4'hff03;
         4'h4518 	:	val_out <= 4'hff00;
         4'h4519 	:	val_out <= 4'hff00;
         4'h451a 	:	val_out <= 4'hff00;
         4'h451b 	:	val_out <= 4'hff00;
         4'h4520 	:	val_out <= 4'hfefd;
         4'h4521 	:	val_out <= 4'hfefd;
         4'h4522 	:	val_out <= 4'hfefd;
         4'h4523 	:	val_out <= 4'hfefd;
         4'h4528 	:	val_out <= 4'hfef9;
         4'h4529 	:	val_out <= 4'hfef9;
         4'h452a 	:	val_out <= 4'hfef9;
         4'h452b 	:	val_out <= 4'hfef9;
         4'h4530 	:	val_out <= 4'hfef6;
         4'h4531 	:	val_out <= 4'hfef6;
         4'h4532 	:	val_out <= 4'hfef6;
         4'h4533 	:	val_out <= 4'hfef6;
         4'h4538 	:	val_out <= 4'hfef3;
         4'h4539 	:	val_out <= 4'hfef3;
         4'h453a 	:	val_out <= 4'hfef3;
         4'h453b 	:	val_out <= 4'hfef3;
         4'h4540 	:	val_out <= 4'hfef0;
         4'h4541 	:	val_out <= 4'hfef0;
         4'h4542 	:	val_out <= 4'hfef0;
         4'h4543 	:	val_out <= 4'hfef0;
         4'h4548 	:	val_out <= 4'hfeed;
         4'h4549 	:	val_out <= 4'hfeed;
         4'h454a 	:	val_out <= 4'hfeed;
         4'h454b 	:	val_out <= 4'hfeed;
         4'h4550 	:	val_out <= 4'hfee9;
         4'h4551 	:	val_out <= 4'hfee9;
         4'h4552 	:	val_out <= 4'hfee9;
         4'h4553 	:	val_out <= 4'hfee9;
         4'h4558 	:	val_out <= 4'hfee6;
         4'h4559 	:	val_out <= 4'hfee6;
         4'h455a 	:	val_out <= 4'hfee6;
         4'h455b 	:	val_out <= 4'hfee6;
         4'h4560 	:	val_out <= 4'hfee3;
         4'h4561 	:	val_out <= 4'hfee3;
         4'h4562 	:	val_out <= 4'hfee3;
         4'h4563 	:	val_out <= 4'hfee3;
         4'h4568 	:	val_out <= 4'hfedf;
         4'h4569 	:	val_out <= 4'hfedf;
         4'h456a 	:	val_out <= 4'hfedf;
         4'h456b 	:	val_out <= 4'hfedf;
         4'h4570 	:	val_out <= 4'hfedc;
         4'h4571 	:	val_out <= 4'hfedc;
         4'h4572 	:	val_out <= 4'hfedc;
         4'h4573 	:	val_out <= 4'hfedc;
         4'h4578 	:	val_out <= 4'hfed9;
         4'h4579 	:	val_out <= 4'hfed9;
         4'h457a 	:	val_out <= 4'hfed9;
         4'h457b 	:	val_out <= 4'hfed9;
         4'h4580 	:	val_out <= 4'hfed5;
         4'h4581 	:	val_out <= 4'hfed5;
         4'h4582 	:	val_out <= 4'hfed5;
         4'h4583 	:	val_out <= 4'hfed5;
         4'h4588 	:	val_out <= 4'hfed2;
         4'h4589 	:	val_out <= 4'hfed2;
         4'h458a 	:	val_out <= 4'hfed2;
         4'h458b 	:	val_out <= 4'hfed2;
         4'h4590 	:	val_out <= 4'hfecf;
         4'h4591 	:	val_out <= 4'hfecf;
         4'h4592 	:	val_out <= 4'hfecf;
         4'h4593 	:	val_out <= 4'hfecf;
         4'h4598 	:	val_out <= 4'hfecb;
         4'h4599 	:	val_out <= 4'hfecb;
         4'h459a 	:	val_out <= 4'hfecb;
         4'h459b 	:	val_out <= 4'hfecb;
         4'h45a0 	:	val_out <= 4'hfec8;
         4'h45a1 	:	val_out <= 4'hfec8;
         4'h45a2 	:	val_out <= 4'hfec8;
         4'h45a3 	:	val_out <= 4'hfec8;
         4'h45a8 	:	val_out <= 4'hfec4;
         4'h45a9 	:	val_out <= 4'hfec4;
         4'h45aa 	:	val_out <= 4'hfec4;
         4'h45ab 	:	val_out <= 4'hfec4;
         4'h45b0 	:	val_out <= 4'hfec1;
         4'h45b1 	:	val_out <= 4'hfec1;
         4'h45b2 	:	val_out <= 4'hfec1;
         4'h45b3 	:	val_out <= 4'hfec1;
         4'h45b8 	:	val_out <= 4'hfebd;
         4'h45b9 	:	val_out <= 4'hfebd;
         4'h45ba 	:	val_out <= 4'hfebd;
         4'h45bb 	:	val_out <= 4'hfebd;
         4'h45c0 	:	val_out <= 4'hfeba;
         4'h45c1 	:	val_out <= 4'hfeba;
         4'h45c2 	:	val_out <= 4'hfeba;
         4'h45c3 	:	val_out <= 4'hfeba;
         4'h45c8 	:	val_out <= 4'hfeb6;
         4'h45c9 	:	val_out <= 4'hfeb6;
         4'h45ca 	:	val_out <= 4'hfeb6;
         4'h45cb 	:	val_out <= 4'hfeb6;
         4'h45d0 	:	val_out <= 4'hfeb3;
         4'h45d1 	:	val_out <= 4'hfeb3;
         4'h45d2 	:	val_out <= 4'hfeb3;
         4'h45d3 	:	val_out <= 4'hfeb3;
         4'h45d8 	:	val_out <= 4'hfeaf;
         4'h45d9 	:	val_out <= 4'hfeaf;
         4'h45da 	:	val_out <= 4'hfeaf;
         4'h45db 	:	val_out <= 4'hfeaf;
         4'h45e0 	:	val_out <= 4'hfeab;
         4'h45e1 	:	val_out <= 4'hfeab;
         4'h45e2 	:	val_out <= 4'hfeab;
         4'h45e3 	:	val_out <= 4'hfeab;
         4'h45e8 	:	val_out <= 4'hfea8;
         4'h45e9 	:	val_out <= 4'hfea8;
         4'h45ea 	:	val_out <= 4'hfea8;
         4'h45eb 	:	val_out <= 4'hfea8;
         4'h45f0 	:	val_out <= 4'hfea4;
         4'h45f1 	:	val_out <= 4'hfea4;
         4'h45f2 	:	val_out <= 4'hfea4;
         4'h45f3 	:	val_out <= 4'hfea4;
         4'h45f8 	:	val_out <= 4'hfea1;
         4'h45f9 	:	val_out <= 4'hfea1;
         4'h45fa 	:	val_out <= 4'hfea1;
         4'h45fb 	:	val_out <= 4'hfea1;
         4'h4600 	:	val_out <= 4'hfe9d;
         4'h4601 	:	val_out <= 4'hfe9d;
         4'h4602 	:	val_out <= 4'hfe9d;
         4'h4603 	:	val_out <= 4'hfe9d;
         4'h4608 	:	val_out <= 4'hfe99;
         4'h4609 	:	val_out <= 4'hfe99;
         4'h460a 	:	val_out <= 4'hfe99;
         4'h460b 	:	val_out <= 4'hfe99;
         4'h4610 	:	val_out <= 4'hfe95;
         4'h4611 	:	val_out <= 4'hfe95;
         4'h4612 	:	val_out <= 4'hfe95;
         4'h4613 	:	val_out <= 4'hfe95;
         4'h4618 	:	val_out <= 4'hfe92;
         4'h4619 	:	val_out <= 4'hfe92;
         4'h461a 	:	val_out <= 4'hfe92;
         4'h461b 	:	val_out <= 4'hfe92;
         4'h4620 	:	val_out <= 4'hfe8e;
         4'h4621 	:	val_out <= 4'hfe8e;
         4'h4622 	:	val_out <= 4'hfe8e;
         4'h4623 	:	val_out <= 4'hfe8e;
         4'h4628 	:	val_out <= 4'hfe8a;
         4'h4629 	:	val_out <= 4'hfe8a;
         4'h462a 	:	val_out <= 4'hfe8a;
         4'h462b 	:	val_out <= 4'hfe8a;
         4'h4630 	:	val_out <= 4'hfe86;
         4'h4631 	:	val_out <= 4'hfe86;
         4'h4632 	:	val_out <= 4'hfe86;
         4'h4633 	:	val_out <= 4'hfe86;
         4'h4638 	:	val_out <= 4'hfe83;
         4'h4639 	:	val_out <= 4'hfe83;
         4'h463a 	:	val_out <= 4'hfe83;
         4'h463b 	:	val_out <= 4'hfe83;
         4'h4640 	:	val_out <= 4'hfe7f;
         4'h4641 	:	val_out <= 4'hfe7f;
         4'h4642 	:	val_out <= 4'hfe7f;
         4'h4643 	:	val_out <= 4'hfe7f;
         4'h4648 	:	val_out <= 4'hfe7b;
         4'h4649 	:	val_out <= 4'hfe7b;
         4'h464a 	:	val_out <= 4'hfe7b;
         4'h464b 	:	val_out <= 4'hfe7b;
         4'h4650 	:	val_out <= 4'hfe77;
         4'h4651 	:	val_out <= 4'hfe77;
         4'h4652 	:	val_out <= 4'hfe77;
         4'h4653 	:	val_out <= 4'hfe77;
         4'h4658 	:	val_out <= 4'hfe73;
         4'h4659 	:	val_out <= 4'hfe73;
         4'h465a 	:	val_out <= 4'hfe73;
         4'h465b 	:	val_out <= 4'hfe73;
         4'h4660 	:	val_out <= 4'hfe6f;
         4'h4661 	:	val_out <= 4'hfe6f;
         4'h4662 	:	val_out <= 4'hfe6f;
         4'h4663 	:	val_out <= 4'hfe6f;
         4'h4668 	:	val_out <= 4'hfe6b;
         4'h4669 	:	val_out <= 4'hfe6b;
         4'h466a 	:	val_out <= 4'hfe6b;
         4'h466b 	:	val_out <= 4'hfe6b;
         4'h4670 	:	val_out <= 4'hfe67;
         4'h4671 	:	val_out <= 4'hfe67;
         4'h4672 	:	val_out <= 4'hfe67;
         4'h4673 	:	val_out <= 4'hfe67;
         4'h4678 	:	val_out <= 4'hfe63;
         4'h4679 	:	val_out <= 4'hfe63;
         4'h467a 	:	val_out <= 4'hfe63;
         4'h467b 	:	val_out <= 4'hfe63;
         4'h4680 	:	val_out <= 4'hfe5f;
         4'h4681 	:	val_out <= 4'hfe5f;
         4'h4682 	:	val_out <= 4'hfe5f;
         4'h4683 	:	val_out <= 4'hfe5f;
         4'h4688 	:	val_out <= 4'hfe5b;
         4'h4689 	:	val_out <= 4'hfe5b;
         4'h468a 	:	val_out <= 4'hfe5b;
         4'h468b 	:	val_out <= 4'hfe5b;
         4'h4690 	:	val_out <= 4'hfe57;
         4'h4691 	:	val_out <= 4'hfe57;
         4'h4692 	:	val_out <= 4'hfe57;
         4'h4693 	:	val_out <= 4'hfe57;
         4'h4698 	:	val_out <= 4'hfe53;
         4'h4699 	:	val_out <= 4'hfe53;
         4'h469a 	:	val_out <= 4'hfe53;
         4'h469b 	:	val_out <= 4'hfe53;
         4'h46a0 	:	val_out <= 4'hfe4f;
         4'h46a1 	:	val_out <= 4'hfe4f;
         4'h46a2 	:	val_out <= 4'hfe4f;
         4'h46a3 	:	val_out <= 4'hfe4f;
         4'h46a8 	:	val_out <= 4'hfe4b;
         4'h46a9 	:	val_out <= 4'hfe4b;
         4'h46aa 	:	val_out <= 4'hfe4b;
         4'h46ab 	:	val_out <= 4'hfe4b;
         4'h46b0 	:	val_out <= 4'hfe47;
         4'h46b1 	:	val_out <= 4'hfe47;
         4'h46b2 	:	val_out <= 4'hfe47;
         4'h46b3 	:	val_out <= 4'hfe47;
         4'h46b8 	:	val_out <= 4'hfe43;
         4'h46b9 	:	val_out <= 4'hfe43;
         4'h46ba 	:	val_out <= 4'hfe43;
         4'h46bb 	:	val_out <= 4'hfe43;
         4'h46c0 	:	val_out <= 4'hfe3f;
         4'h46c1 	:	val_out <= 4'hfe3f;
         4'h46c2 	:	val_out <= 4'hfe3f;
         4'h46c3 	:	val_out <= 4'hfe3f;
         4'h46c8 	:	val_out <= 4'hfe3b;
         4'h46c9 	:	val_out <= 4'hfe3b;
         4'h46ca 	:	val_out <= 4'hfe3b;
         4'h46cb 	:	val_out <= 4'hfe3b;
         4'h46d0 	:	val_out <= 4'hfe37;
         4'h46d1 	:	val_out <= 4'hfe37;
         4'h46d2 	:	val_out <= 4'hfe37;
         4'h46d3 	:	val_out <= 4'hfe37;
         4'h46d8 	:	val_out <= 4'hfe32;
         4'h46d9 	:	val_out <= 4'hfe32;
         4'h46da 	:	val_out <= 4'hfe32;
         4'h46db 	:	val_out <= 4'hfe32;
         4'h46e0 	:	val_out <= 4'hfe2e;
         4'h46e1 	:	val_out <= 4'hfe2e;
         4'h46e2 	:	val_out <= 4'hfe2e;
         4'h46e3 	:	val_out <= 4'hfe2e;
         4'h46e8 	:	val_out <= 4'hfe2a;
         4'h46e9 	:	val_out <= 4'hfe2a;
         4'h46ea 	:	val_out <= 4'hfe2a;
         4'h46eb 	:	val_out <= 4'hfe2a;
         4'h46f0 	:	val_out <= 4'hfe26;
         4'h46f1 	:	val_out <= 4'hfe26;
         4'h46f2 	:	val_out <= 4'hfe26;
         4'h46f3 	:	val_out <= 4'hfe26;
         4'h46f8 	:	val_out <= 4'hfe21;
         4'h46f9 	:	val_out <= 4'hfe21;
         4'h46fa 	:	val_out <= 4'hfe21;
         4'h46fb 	:	val_out <= 4'hfe21;
         4'h4700 	:	val_out <= 4'hfe1d;
         4'h4701 	:	val_out <= 4'hfe1d;
         4'h4702 	:	val_out <= 4'hfe1d;
         4'h4703 	:	val_out <= 4'hfe1d;
         4'h4708 	:	val_out <= 4'hfe19;
         4'h4709 	:	val_out <= 4'hfe19;
         4'h470a 	:	val_out <= 4'hfe19;
         4'h470b 	:	val_out <= 4'hfe19;
         4'h4710 	:	val_out <= 4'hfe14;
         4'h4711 	:	val_out <= 4'hfe14;
         4'h4712 	:	val_out <= 4'hfe14;
         4'h4713 	:	val_out <= 4'hfe14;
         4'h4718 	:	val_out <= 4'hfe10;
         4'h4719 	:	val_out <= 4'hfe10;
         4'h471a 	:	val_out <= 4'hfe10;
         4'h471b 	:	val_out <= 4'hfe10;
         4'h4720 	:	val_out <= 4'hfe0c;
         4'h4721 	:	val_out <= 4'hfe0c;
         4'h4722 	:	val_out <= 4'hfe0c;
         4'h4723 	:	val_out <= 4'hfe0c;
         4'h4728 	:	val_out <= 4'hfe07;
         4'h4729 	:	val_out <= 4'hfe07;
         4'h472a 	:	val_out <= 4'hfe07;
         4'h472b 	:	val_out <= 4'hfe07;
         4'h4730 	:	val_out <= 4'hfe03;
         4'h4731 	:	val_out <= 4'hfe03;
         4'h4732 	:	val_out <= 4'hfe03;
         4'h4733 	:	val_out <= 4'hfe03;
         4'h4738 	:	val_out <= 4'hfdff;
         4'h4739 	:	val_out <= 4'hfdff;
         4'h473a 	:	val_out <= 4'hfdff;
         4'h473b 	:	val_out <= 4'hfdff;
         4'h4740 	:	val_out <= 4'hfdfa;
         4'h4741 	:	val_out <= 4'hfdfa;
         4'h4742 	:	val_out <= 4'hfdfa;
         4'h4743 	:	val_out <= 4'hfdfa;
         4'h4748 	:	val_out <= 4'hfdf6;
         4'h4749 	:	val_out <= 4'hfdf6;
         4'h474a 	:	val_out <= 4'hfdf6;
         4'h474b 	:	val_out <= 4'hfdf6;
         4'h4750 	:	val_out <= 4'hfdf1;
         4'h4751 	:	val_out <= 4'hfdf1;
         4'h4752 	:	val_out <= 4'hfdf1;
         4'h4753 	:	val_out <= 4'hfdf1;
         4'h4758 	:	val_out <= 4'hfded;
         4'h4759 	:	val_out <= 4'hfded;
         4'h475a 	:	val_out <= 4'hfded;
         4'h475b 	:	val_out <= 4'hfded;
         4'h4760 	:	val_out <= 4'hfde8;
         4'h4761 	:	val_out <= 4'hfde8;
         4'h4762 	:	val_out <= 4'hfde8;
         4'h4763 	:	val_out <= 4'hfde8;
         4'h4768 	:	val_out <= 4'hfde4;
         4'h4769 	:	val_out <= 4'hfde4;
         4'h476a 	:	val_out <= 4'hfde4;
         4'h476b 	:	val_out <= 4'hfde4;
         4'h4770 	:	val_out <= 4'hfddf;
         4'h4771 	:	val_out <= 4'hfddf;
         4'h4772 	:	val_out <= 4'hfddf;
         4'h4773 	:	val_out <= 4'hfddf;
         4'h4778 	:	val_out <= 4'hfdda;
         4'h4779 	:	val_out <= 4'hfdda;
         4'h477a 	:	val_out <= 4'hfdda;
         4'h477b 	:	val_out <= 4'hfdda;
         4'h4780 	:	val_out <= 4'hfdd6;
         4'h4781 	:	val_out <= 4'hfdd6;
         4'h4782 	:	val_out <= 4'hfdd6;
         4'h4783 	:	val_out <= 4'hfdd6;
         4'h4788 	:	val_out <= 4'hfdd1;
         4'h4789 	:	val_out <= 4'hfdd1;
         4'h478a 	:	val_out <= 4'hfdd1;
         4'h478b 	:	val_out <= 4'hfdd1;
         4'h4790 	:	val_out <= 4'hfdcd;
         4'h4791 	:	val_out <= 4'hfdcd;
         4'h4792 	:	val_out <= 4'hfdcd;
         4'h4793 	:	val_out <= 4'hfdcd;
         4'h4798 	:	val_out <= 4'hfdc8;
         4'h4799 	:	val_out <= 4'hfdc8;
         4'h479a 	:	val_out <= 4'hfdc8;
         4'h479b 	:	val_out <= 4'hfdc8;
         4'h47a0 	:	val_out <= 4'hfdc3;
         4'h47a1 	:	val_out <= 4'hfdc3;
         4'h47a2 	:	val_out <= 4'hfdc3;
         4'h47a3 	:	val_out <= 4'hfdc3;
         4'h47a8 	:	val_out <= 4'hfdbf;
         4'h47a9 	:	val_out <= 4'hfdbf;
         4'h47aa 	:	val_out <= 4'hfdbf;
         4'h47ab 	:	val_out <= 4'hfdbf;
         4'h47b0 	:	val_out <= 4'hfdba;
         4'h47b1 	:	val_out <= 4'hfdba;
         4'h47b2 	:	val_out <= 4'hfdba;
         4'h47b3 	:	val_out <= 4'hfdba;
         4'h47b8 	:	val_out <= 4'hfdb5;
         4'h47b9 	:	val_out <= 4'hfdb5;
         4'h47ba 	:	val_out <= 4'hfdb5;
         4'h47bb 	:	val_out <= 4'hfdb5;
         4'h47c0 	:	val_out <= 4'hfdb0;
         4'h47c1 	:	val_out <= 4'hfdb0;
         4'h47c2 	:	val_out <= 4'hfdb0;
         4'h47c3 	:	val_out <= 4'hfdb0;
         4'h47c8 	:	val_out <= 4'hfdac;
         4'h47c9 	:	val_out <= 4'hfdac;
         4'h47ca 	:	val_out <= 4'hfdac;
         4'h47cb 	:	val_out <= 4'hfdac;
         4'h47d0 	:	val_out <= 4'hfda7;
         4'h47d1 	:	val_out <= 4'hfda7;
         4'h47d2 	:	val_out <= 4'hfda7;
         4'h47d3 	:	val_out <= 4'hfda7;
         4'h47d8 	:	val_out <= 4'hfda2;
         4'h47d9 	:	val_out <= 4'hfda2;
         4'h47da 	:	val_out <= 4'hfda2;
         4'h47db 	:	val_out <= 4'hfda2;
         4'h47e0 	:	val_out <= 4'hfd9d;
         4'h47e1 	:	val_out <= 4'hfd9d;
         4'h47e2 	:	val_out <= 4'hfd9d;
         4'h47e3 	:	val_out <= 4'hfd9d;
         4'h47e8 	:	val_out <= 4'hfd98;
         4'h47e9 	:	val_out <= 4'hfd98;
         4'h47ea 	:	val_out <= 4'hfd98;
         4'h47eb 	:	val_out <= 4'hfd98;
         4'h47f0 	:	val_out <= 4'hfd94;
         4'h47f1 	:	val_out <= 4'hfd94;
         4'h47f2 	:	val_out <= 4'hfd94;
         4'h47f3 	:	val_out <= 4'hfd94;
         4'h47f8 	:	val_out <= 4'hfd8f;
         4'h47f9 	:	val_out <= 4'hfd8f;
         4'h47fa 	:	val_out <= 4'hfd8f;
         4'h47fb 	:	val_out <= 4'hfd8f;
         4'h4800 	:	val_out <= 4'hfd8a;
         4'h4801 	:	val_out <= 4'hfd8a;
         4'h4802 	:	val_out <= 4'hfd8a;
         4'h4803 	:	val_out <= 4'hfd8a;
         4'h4808 	:	val_out <= 4'hfd85;
         4'h4809 	:	val_out <= 4'hfd85;
         4'h480a 	:	val_out <= 4'hfd85;
         4'h480b 	:	val_out <= 4'hfd85;
         4'h4810 	:	val_out <= 4'hfd80;
         4'h4811 	:	val_out <= 4'hfd80;
         4'h4812 	:	val_out <= 4'hfd80;
         4'h4813 	:	val_out <= 4'hfd80;
         4'h4818 	:	val_out <= 4'hfd7b;
         4'h4819 	:	val_out <= 4'hfd7b;
         4'h481a 	:	val_out <= 4'hfd7b;
         4'h481b 	:	val_out <= 4'hfd7b;
         4'h4820 	:	val_out <= 4'hfd76;
         4'h4821 	:	val_out <= 4'hfd76;
         4'h4822 	:	val_out <= 4'hfd76;
         4'h4823 	:	val_out <= 4'hfd76;
         4'h4828 	:	val_out <= 4'hfd71;
         4'h4829 	:	val_out <= 4'hfd71;
         4'h482a 	:	val_out <= 4'hfd71;
         4'h482b 	:	val_out <= 4'hfd71;
         4'h4830 	:	val_out <= 4'hfd6c;
         4'h4831 	:	val_out <= 4'hfd6c;
         4'h4832 	:	val_out <= 4'hfd6c;
         4'h4833 	:	val_out <= 4'hfd6c;
         4'h4838 	:	val_out <= 4'hfd67;
         4'h4839 	:	val_out <= 4'hfd67;
         4'h483a 	:	val_out <= 4'hfd67;
         4'h483b 	:	val_out <= 4'hfd67;
         4'h4840 	:	val_out <= 4'hfd62;
         4'h4841 	:	val_out <= 4'hfd62;
         4'h4842 	:	val_out <= 4'hfd62;
         4'h4843 	:	val_out <= 4'hfd62;
         4'h4848 	:	val_out <= 4'hfd5d;
         4'h4849 	:	val_out <= 4'hfd5d;
         4'h484a 	:	val_out <= 4'hfd5d;
         4'h484b 	:	val_out <= 4'hfd5d;
         4'h4850 	:	val_out <= 4'hfd58;
         4'h4851 	:	val_out <= 4'hfd58;
         4'h4852 	:	val_out <= 4'hfd58;
         4'h4853 	:	val_out <= 4'hfd58;
         4'h4858 	:	val_out <= 4'hfd53;
         4'h4859 	:	val_out <= 4'hfd53;
         4'h485a 	:	val_out <= 4'hfd53;
         4'h485b 	:	val_out <= 4'hfd53;
         4'h4860 	:	val_out <= 4'hfd4e;
         4'h4861 	:	val_out <= 4'hfd4e;
         4'h4862 	:	val_out <= 4'hfd4e;
         4'h4863 	:	val_out <= 4'hfd4e;
         4'h4868 	:	val_out <= 4'hfd49;
         4'h4869 	:	val_out <= 4'hfd49;
         4'h486a 	:	val_out <= 4'hfd49;
         4'h486b 	:	val_out <= 4'hfd49;
         4'h4870 	:	val_out <= 4'hfd43;
         4'h4871 	:	val_out <= 4'hfd43;
         4'h4872 	:	val_out <= 4'hfd43;
         4'h4873 	:	val_out <= 4'hfd43;
         4'h4878 	:	val_out <= 4'hfd3e;
         4'h4879 	:	val_out <= 4'hfd3e;
         4'h487a 	:	val_out <= 4'hfd3e;
         4'h487b 	:	val_out <= 4'hfd3e;
         4'h4880 	:	val_out <= 4'hfd39;
         4'h4881 	:	val_out <= 4'hfd39;
         4'h4882 	:	val_out <= 4'hfd39;
         4'h4883 	:	val_out <= 4'hfd39;
         4'h4888 	:	val_out <= 4'hfd34;
         4'h4889 	:	val_out <= 4'hfd34;
         4'h488a 	:	val_out <= 4'hfd34;
         4'h488b 	:	val_out <= 4'hfd34;
         4'h4890 	:	val_out <= 4'hfd2f;
         4'h4891 	:	val_out <= 4'hfd2f;
         4'h4892 	:	val_out <= 4'hfd2f;
         4'h4893 	:	val_out <= 4'hfd2f;
         4'h4898 	:	val_out <= 4'hfd29;
         4'h4899 	:	val_out <= 4'hfd29;
         4'h489a 	:	val_out <= 4'hfd29;
         4'h489b 	:	val_out <= 4'hfd29;
         4'h48a0 	:	val_out <= 4'hfd24;
         4'h48a1 	:	val_out <= 4'hfd24;
         4'h48a2 	:	val_out <= 4'hfd24;
         4'h48a3 	:	val_out <= 4'hfd24;
         4'h48a8 	:	val_out <= 4'hfd1f;
         4'h48a9 	:	val_out <= 4'hfd1f;
         4'h48aa 	:	val_out <= 4'hfd1f;
         4'h48ab 	:	val_out <= 4'hfd1f;
         4'h48b0 	:	val_out <= 4'hfd19;
         4'h48b1 	:	val_out <= 4'hfd19;
         4'h48b2 	:	val_out <= 4'hfd19;
         4'h48b3 	:	val_out <= 4'hfd19;
         4'h48b8 	:	val_out <= 4'hfd14;
         4'h48b9 	:	val_out <= 4'hfd14;
         4'h48ba 	:	val_out <= 4'hfd14;
         4'h48bb 	:	val_out <= 4'hfd14;
         4'h48c0 	:	val_out <= 4'hfd0f;
         4'h48c1 	:	val_out <= 4'hfd0f;
         4'h48c2 	:	val_out <= 4'hfd0f;
         4'h48c3 	:	val_out <= 4'hfd0f;
         4'h48c8 	:	val_out <= 4'hfd09;
         4'h48c9 	:	val_out <= 4'hfd09;
         4'h48ca 	:	val_out <= 4'hfd09;
         4'h48cb 	:	val_out <= 4'hfd09;
         4'h48d0 	:	val_out <= 4'hfd04;
         4'h48d1 	:	val_out <= 4'hfd04;
         4'h48d2 	:	val_out <= 4'hfd04;
         4'h48d3 	:	val_out <= 4'hfd04;
         4'h48d8 	:	val_out <= 4'hfcff;
         4'h48d9 	:	val_out <= 4'hfcff;
         4'h48da 	:	val_out <= 4'hfcff;
         4'h48db 	:	val_out <= 4'hfcff;
         4'h48e0 	:	val_out <= 4'hfcf9;
         4'h48e1 	:	val_out <= 4'hfcf9;
         4'h48e2 	:	val_out <= 4'hfcf9;
         4'h48e3 	:	val_out <= 4'hfcf9;
         4'h48e8 	:	val_out <= 4'hfcf4;
         4'h48e9 	:	val_out <= 4'hfcf4;
         4'h48ea 	:	val_out <= 4'hfcf4;
         4'h48eb 	:	val_out <= 4'hfcf4;
         4'h48f0 	:	val_out <= 4'hfcee;
         4'h48f1 	:	val_out <= 4'hfcee;
         4'h48f2 	:	val_out <= 4'hfcee;
         4'h48f3 	:	val_out <= 4'hfcee;
         4'h48f8 	:	val_out <= 4'hfce9;
         4'h48f9 	:	val_out <= 4'hfce9;
         4'h48fa 	:	val_out <= 4'hfce9;
         4'h48fb 	:	val_out <= 4'hfce9;
         4'h4900 	:	val_out <= 4'hfce3;
         4'h4901 	:	val_out <= 4'hfce3;
         4'h4902 	:	val_out <= 4'hfce3;
         4'h4903 	:	val_out <= 4'hfce3;
         4'h4908 	:	val_out <= 4'hfcde;
         4'h4909 	:	val_out <= 4'hfcde;
         4'h490a 	:	val_out <= 4'hfcde;
         4'h490b 	:	val_out <= 4'hfcde;
         4'h4910 	:	val_out <= 4'hfcd8;
         4'h4911 	:	val_out <= 4'hfcd8;
         4'h4912 	:	val_out <= 4'hfcd8;
         4'h4913 	:	val_out <= 4'hfcd8;
         4'h4918 	:	val_out <= 4'hfcd3;
         4'h4919 	:	val_out <= 4'hfcd3;
         4'h491a 	:	val_out <= 4'hfcd3;
         4'h491b 	:	val_out <= 4'hfcd3;
         4'h4920 	:	val_out <= 4'hfccd;
         4'h4921 	:	val_out <= 4'hfccd;
         4'h4922 	:	val_out <= 4'hfccd;
         4'h4923 	:	val_out <= 4'hfccd;
         4'h4928 	:	val_out <= 4'hfcc8;
         4'h4929 	:	val_out <= 4'hfcc8;
         4'h492a 	:	val_out <= 4'hfcc8;
         4'h492b 	:	val_out <= 4'hfcc8;
         4'h4930 	:	val_out <= 4'hfcc2;
         4'h4931 	:	val_out <= 4'hfcc2;
         4'h4932 	:	val_out <= 4'hfcc2;
         4'h4933 	:	val_out <= 4'hfcc2;
         4'h4938 	:	val_out <= 4'hfcbc;
         4'h4939 	:	val_out <= 4'hfcbc;
         4'h493a 	:	val_out <= 4'hfcbc;
         4'h493b 	:	val_out <= 4'hfcbc;
         4'h4940 	:	val_out <= 4'hfcb7;
         4'h4941 	:	val_out <= 4'hfcb7;
         4'h4942 	:	val_out <= 4'hfcb7;
         4'h4943 	:	val_out <= 4'hfcb7;
         4'h4948 	:	val_out <= 4'hfcb1;
         4'h4949 	:	val_out <= 4'hfcb1;
         4'h494a 	:	val_out <= 4'hfcb1;
         4'h494b 	:	val_out <= 4'hfcb1;
         4'h4950 	:	val_out <= 4'hfcab;
         4'h4951 	:	val_out <= 4'hfcab;
         4'h4952 	:	val_out <= 4'hfcab;
         4'h4953 	:	val_out <= 4'hfcab;
         4'h4958 	:	val_out <= 4'hfca6;
         4'h4959 	:	val_out <= 4'hfca6;
         4'h495a 	:	val_out <= 4'hfca6;
         4'h495b 	:	val_out <= 4'hfca6;
         4'h4960 	:	val_out <= 4'hfca0;
         4'h4961 	:	val_out <= 4'hfca0;
         4'h4962 	:	val_out <= 4'hfca0;
         4'h4963 	:	val_out <= 4'hfca0;
         4'h4968 	:	val_out <= 4'hfc9a;
         4'h4969 	:	val_out <= 4'hfc9a;
         4'h496a 	:	val_out <= 4'hfc9a;
         4'h496b 	:	val_out <= 4'hfc9a;
         4'h4970 	:	val_out <= 4'hfc94;
         4'h4971 	:	val_out <= 4'hfc94;
         4'h4972 	:	val_out <= 4'hfc94;
         4'h4973 	:	val_out <= 4'hfc94;
         4'h4978 	:	val_out <= 4'hfc8f;
         4'h4979 	:	val_out <= 4'hfc8f;
         4'h497a 	:	val_out <= 4'hfc8f;
         4'h497b 	:	val_out <= 4'hfc8f;
         4'h4980 	:	val_out <= 4'hfc89;
         4'h4981 	:	val_out <= 4'hfc89;
         4'h4982 	:	val_out <= 4'hfc89;
         4'h4983 	:	val_out <= 4'hfc89;
         4'h4988 	:	val_out <= 4'hfc83;
         4'h4989 	:	val_out <= 4'hfc83;
         4'h498a 	:	val_out <= 4'hfc83;
         4'h498b 	:	val_out <= 4'hfc83;
         4'h4990 	:	val_out <= 4'hfc7d;
         4'h4991 	:	val_out <= 4'hfc7d;
         4'h4992 	:	val_out <= 4'hfc7d;
         4'h4993 	:	val_out <= 4'hfc7d;
         4'h4998 	:	val_out <= 4'hfc77;
         4'h4999 	:	val_out <= 4'hfc77;
         4'h499a 	:	val_out <= 4'hfc77;
         4'h499b 	:	val_out <= 4'hfc77;
         4'h49a0 	:	val_out <= 4'hfc71;
         4'h49a1 	:	val_out <= 4'hfc71;
         4'h49a2 	:	val_out <= 4'hfc71;
         4'h49a3 	:	val_out <= 4'hfc71;
         4'h49a8 	:	val_out <= 4'hfc6c;
         4'h49a9 	:	val_out <= 4'hfc6c;
         4'h49aa 	:	val_out <= 4'hfc6c;
         4'h49ab 	:	val_out <= 4'hfc6c;
         4'h49b0 	:	val_out <= 4'hfc66;
         4'h49b1 	:	val_out <= 4'hfc66;
         4'h49b2 	:	val_out <= 4'hfc66;
         4'h49b3 	:	val_out <= 4'hfc66;
         4'h49b8 	:	val_out <= 4'hfc60;
         4'h49b9 	:	val_out <= 4'hfc60;
         4'h49ba 	:	val_out <= 4'hfc60;
         4'h49bb 	:	val_out <= 4'hfc60;
         4'h49c0 	:	val_out <= 4'hfc5a;
         4'h49c1 	:	val_out <= 4'hfc5a;
         4'h49c2 	:	val_out <= 4'hfc5a;
         4'h49c3 	:	val_out <= 4'hfc5a;
         4'h49c8 	:	val_out <= 4'hfc54;
         4'h49c9 	:	val_out <= 4'hfc54;
         4'h49ca 	:	val_out <= 4'hfc54;
         4'h49cb 	:	val_out <= 4'hfc54;
         4'h49d0 	:	val_out <= 4'hfc4e;
         4'h49d1 	:	val_out <= 4'hfc4e;
         4'h49d2 	:	val_out <= 4'hfc4e;
         4'h49d3 	:	val_out <= 4'hfc4e;
         4'h49d8 	:	val_out <= 4'hfc48;
         4'h49d9 	:	val_out <= 4'hfc48;
         4'h49da 	:	val_out <= 4'hfc48;
         4'h49db 	:	val_out <= 4'hfc48;
         4'h49e0 	:	val_out <= 4'hfc42;
         4'h49e1 	:	val_out <= 4'hfc42;
         4'h49e2 	:	val_out <= 4'hfc42;
         4'h49e3 	:	val_out <= 4'hfc42;
         4'h49e8 	:	val_out <= 4'hfc3c;
         4'h49e9 	:	val_out <= 4'hfc3c;
         4'h49ea 	:	val_out <= 4'hfc3c;
         4'h49eb 	:	val_out <= 4'hfc3c;
         4'h49f0 	:	val_out <= 4'hfc36;
         4'h49f1 	:	val_out <= 4'hfc36;
         4'h49f2 	:	val_out <= 4'hfc36;
         4'h49f3 	:	val_out <= 4'hfc36;
         4'h49f8 	:	val_out <= 4'hfc30;
         4'h49f9 	:	val_out <= 4'hfc30;
         4'h49fa 	:	val_out <= 4'hfc30;
         4'h49fb 	:	val_out <= 4'hfc30;
         4'h4a00 	:	val_out <= 4'hfc29;
         4'h4a01 	:	val_out <= 4'hfc29;
         4'h4a02 	:	val_out <= 4'hfc29;
         4'h4a03 	:	val_out <= 4'hfc29;
         4'h4a08 	:	val_out <= 4'hfc23;
         4'h4a09 	:	val_out <= 4'hfc23;
         4'h4a0a 	:	val_out <= 4'hfc23;
         4'h4a0b 	:	val_out <= 4'hfc23;
         4'h4a10 	:	val_out <= 4'hfc1d;
         4'h4a11 	:	val_out <= 4'hfc1d;
         4'h4a12 	:	val_out <= 4'hfc1d;
         4'h4a13 	:	val_out <= 4'hfc1d;
         4'h4a18 	:	val_out <= 4'hfc17;
         4'h4a19 	:	val_out <= 4'hfc17;
         4'h4a1a 	:	val_out <= 4'hfc17;
         4'h4a1b 	:	val_out <= 4'hfc17;
         4'h4a20 	:	val_out <= 4'hfc11;
         4'h4a21 	:	val_out <= 4'hfc11;
         4'h4a22 	:	val_out <= 4'hfc11;
         4'h4a23 	:	val_out <= 4'hfc11;
         4'h4a28 	:	val_out <= 4'hfc0b;
         4'h4a29 	:	val_out <= 4'hfc0b;
         4'h4a2a 	:	val_out <= 4'hfc0b;
         4'h4a2b 	:	val_out <= 4'hfc0b;
         4'h4a30 	:	val_out <= 4'hfc05;
         4'h4a31 	:	val_out <= 4'hfc05;
         4'h4a32 	:	val_out <= 4'hfc05;
         4'h4a33 	:	val_out <= 4'hfc05;
         4'h4a38 	:	val_out <= 4'hfbfe;
         4'h4a39 	:	val_out <= 4'hfbfe;
         4'h4a3a 	:	val_out <= 4'hfbfe;
         4'h4a3b 	:	val_out <= 4'hfbfe;
         4'h4a40 	:	val_out <= 4'hfbf8;
         4'h4a41 	:	val_out <= 4'hfbf8;
         4'h4a42 	:	val_out <= 4'hfbf8;
         4'h4a43 	:	val_out <= 4'hfbf8;
         4'h4a48 	:	val_out <= 4'hfbf2;
         4'h4a49 	:	val_out <= 4'hfbf2;
         4'h4a4a 	:	val_out <= 4'hfbf2;
         4'h4a4b 	:	val_out <= 4'hfbf2;
         4'h4a50 	:	val_out <= 4'hfbeb;
         4'h4a51 	:	val_out <= 4'hfbeb;
         4'h4a52 	:	val_out <= 4'hfbeb;
         4'h4a53 	:	val_out <= 4'hfbeb;
         4'h4a58 	:	val_out <= 4'hfbe5;
         4'h4a59 	:	val_out <= 4'hfbe5;
         4'h4a5a 	:	val_out <= 4'hfbe5;
         4'h4a5b 	:	val_out <= 4'hfbe5;
         4'h4a60 	:	val_out <= 4'hfbdf;
         4'h4a61 	:	val_out <= 4'hfbdf;
         4'h4a62 	:	val_out <= 4'hfbdf;
         4'h4a63 	:	val_out <= 4'hfbdf;
         4'h4a68 	:	val_out <= 4'hfbd9;
         4'h4a69 	:	val_out <= 4'hfbd9;
         4'h4a6a 	:	val_out <= 4'hfbd9;
         4'h4a6b 	:	val_out <= 4'hfbd9;
         4'h4a70 	:	val_out <= 4'hfbd2;
         4'h4a71 	:	val_out <= 4'hfbd2;
         4'h4a72 	:	val_out <= 4'hfbd2;
         4'h4a73 	:	val_out <= 4'hfbd2;
         4'h4a78 	:	val_out <= 4'hfbcc;
         4'h4a79 	:	val_out <= 4'hfbcc;
         4'h4a7a 	:	val_out <= 4'hfbcc;
         4'h4a7b 	:	val_out <= 4'hfbcc;
         4'h4a80 	:	val_out <= 4'hfbc5;
         4'h4a81 	:	val_out <= 4'hfbc5;
         4'h4a82 	:	val_out <= 4'hfbc5;
         4'h4a83 	:	val_out <= 4'hfbc5;
         4'h4a88 	:	val_out <= 4'hfbbf;
         4'h4a89 	:	val_out <= 4'hfbbf;
         4'h4a8a 	:	val_out <= 4'hfbbf;
         4'h4a8b 	:	val_out <= 4'hfbbf;
         4'h4a90 	:	val_out <= 4'hfbb9;
         4'h4a91 	:	val_out <= 4'hfbb9;
         4'h4a92 	:	val_out <= 4'hfbb9;
         4'h4a93 	:	val_out <= 4'hfbb9;
         4'h4a98 	:	val_out <= 4'hfbb2;
         4'h4a99 	:	val_out <= 4'hfbb2;
         4'h4a9a 	:	val_out <= 4'hfbb2;
         4'h4a9b 	:	val_out <= 4'hfbb2;
         4'h4aa0 	:	val_out <= 4'hfbac;
         4'h4aa1 	:	val_out <= 4'hfbac;
         4'h4aa2 	:	val_out <= 4'hfbac;
         4'h4aa3 	:	val_out <= 4'hfbac;
         4'h4aa8 	:	val_out <= 4'hfba5;
         4'h4aa9 	:	val_out <= 4'hfba5;
         4'h4aaa 	:	val_out <= 4'hfba5;
         4'h4aab 	:	val_out <= 4'hfba5;
         4'h4ab0 	:	val_out <= 4'hfb9f;
         4'h4ab1 	:	val_out <= 4'hfb9f;
         4'h4ab2 	:	val_out <= 4'hfb9f;
         4'h4ab3 	:	val_out <= 4'hfb9f;
         4'h4ab8 	:	val_out <= 4'hfb98;
         4'h4ab9 	:	val_out <= 4'hfb98;
         4'h4aba 	:	val_out <= 4'hfb98;
         4'h4abb 	:	val_out <= 4'hfb98;
         4'h4ac0 	:	val_out <= 4'hfb92;
         4'h4ac1 	:	val_out <= 4'hfb92;
         4'h4ac2 	:	val_out <= 4'hfb92;
         4'h4ac3 	:	val_out <= 4'hfb92;
         4'h4ac8 	:	val_out <= 4'hfb8b;
         4'h4ac9 	:	val_out <= 4'hfb8b;
         4'h4aca 	:	val_out <= 4'hfb8b;
         4'h4acb 	:	val_out <= 4'hfb8b;
         4'h4ad0 	:	val_out <= 4'hfb84;
         4'h4ad1 	:	val_out <= 4'hfb84;
         4'h4ad2 	:	val_out <= 4'hfb84;
         4'h4ad3 	:	val_out <= 4'hfb84;
         4'h4ad8 	:	val_out <= 4'hfb7e;
         4'h4ad9 	:	val_out <= 4'hfb7e;
         4'h4ada 	:	val_out <= 4'hfb7e;
         4'h4adb 	:	val_out <= 4'hfb7e;
         4'h4ae0 	:	val_out <= 4'hfb77;
         4'h4ae1 	:	val_out <= 4'hfb77;
         4'h4ae2 	:	val_out <= 4'hfb77;
         4'h4ae3 	:	val_out <= 4'hfb77;
         4'h4ae8 	:	val_out <= 4'hfb71;
         4'h4ae9 	:	val_out <= 4'hfb71;
         4'h4aea 	:	val_out <= 4'hfb71;
         4'h4aeb 	:	val_out <= 4'hfb71;
         4'h4af0 	:	val_out <= 4'hfb6a;
         4'h4af1 	:	val_out <= 4'hfb6a;
         4'h4af2 	:	val_out <= 4'hfb6a;
         4'h4af3 	:	val_out <= 4'hfb6a;
         4'h4af8 	:	val_out <= 4'hfb63;
         4'h4af9 	:	val_out <= 4'hfb63;
         4'h4afa 	:	val_out <= 4'hfb63;
         4'h4afb 	:	val_out <= 4'hfb63;
         4'h4b00 	:	val_out <= 4'hfb5d;
         4'h4b01 	:	val_out <= 4'hfb5d;
         4'h4b02 	:	val_out <= 4'hfb5d;
         4'h4b03 	:	val_out <= 4'hfb5d;
         4'h4b08 	:	val_out <= 4'hfb56;
         4'h4b09 	:	val_out <= 4'hfb56;
         4'h4b0a 	:	val_out <= 4'hfb56;
         4'h4b0b 	:	val_out <= 4'hfb56;
         4'h4b10 	:	val_out <= 4'hfb4f;
         4'h4b11 	:	val_out <= 4'hfb4f;
         4'h4b12 	:	val_out <= 4'hfb4f;
         4'h4b13 	:	val_out <= 4'hfb4f;
         4'h4b18 	:	val_out <= 4'hfb48;
         4'h4b19 	:	val_out <= 4'hfb48;
         4'h4b1a 	:	val_out <= 4'hfb48;
         4'h4b1b 	:	val_out <= 4'hfb48;
         4'h4b20 	:	val_out <= 4'hfb42;
         4'h4b21 	:	val_out <= 4'hfb42;
         4'h4b22 	:	val_out <= 4'hfb42;
         4'h4b23 	:	val_out <= 4'hfb42;
         4'h4b28 	:	val_out <= 4'hfb3b;
         4'h4b29 	:	val_out <= 4'hfb3b;
         4'h4b2a 	:	val_out <= 4'hfb3b;
         4'h4b2b 	:	val_out <= 4'hfb3b;
         4'h4b30 	:	val_out <= 4'hfb34;
         4'h4b31 	:	val_out <= 4'hfb34;
         4'h4b32 	:	val_out <= 4'hfb34;
         4'h4b33 	:	val_out <= 4'hfb34;
         4'h4b38 	:	val_out <= 4'hfb2d;
         4'h4b39 	:	val_out <= 4'hfb2d;
         4'h4b3a 	:	val_out <= 4'hfb2d;
         4'h4b3b 	:	val_out <= 4'hfb2d;
         4'h4b40 	:	val_out <= 4'hfb26;
         4'h4b41 	:	val_out <= 4'hfb26;
         4'h4b42 	:	val_out <= 4'hfb26;
         4'h4b43 	:	val_out <= 4'hfb26;
         4'h4b48 	:	val_out <= 4'hfb1f;
         4'h4b49 	:	val_out <= 4'hfb1f;
         4'h4b4a 	:	val_out <= 4'hfb1f;
         4'h4b4b 	:	val_out <= 4'hfb1f;
         4'h4b50 	:	val_out <= 4'hfb19;
         4'h4b51 	:	val_out <= 4'hfb19;
         4'h4b52 	:	val_out <= 4'hfb19;
         4'h4b53 	:	val_out <= 4'hfb19;
         4'h4b58 	:	val_out <= 4'hfb12;
         4'h4b59 	:	val_out <= 4'hfb12;
         4'h4b5a 	:	val_out <= 4'hfb12;
         4'h4b5b 	:	val_out <= 4'hfb12;
         4'h4b60 	:	val_out <= 4'hfb0b;
         4'h4b61 	:	val_out <= 4'hfb0b;
         4'h4b62 	:	val_out <= 4'hfb0b;
         4'h4b63 	:	val_out <= 4'hfb0b;
         4'h4b68 	:	val_out <= 4'hfb04;
         4'h4b69 	:	val_out <= 4'hfb04;
         4'h4b6a 	:	val_out <= 4'hfb04;
         4'h4b6b 	:	val_out <= 4'hfb04;
         4'h4b70 	:	val_out <= 4'hfafd;
         4'h4b71 	:	val_out <= 4'hfafd;
         4'h4b72 	:	val_out <= 4'hfafd;
         4'h4b73 	:	val_out <= 4'hfafd;
         4'h4b78 	:	val_out <= 4'hfaf6;
         4'h4b79 	:	val_out <= 4'hfaf6;
         4'h4b7a 	:	val_out <= 4'hfaf6;
         4'h4b7b 	:	val_out <= 4'hfaf6;
         4'h4b80 	:	val_out <= 4'hfaef;
         4'h4b81 	:	val_out <= 4'hfaef;
         4'h4b82 	:	val_out <= 4'hfaef;
         4'h4b83 	:	val_out <= 4'hfaef;
         4'h4b88 	:	val_out <= 4'hfae8;
         4'h4b89 	:	val_out <= 4'hfae8;
         4'h4b8a 	:	val_out <= 4'hfae8;
         4'h4b8b 	:	val_out <= 4'hfae8;
         4'h4b90 	:	val_out <= 4'hfae1;
         4'h4b91 	:	val_out <= 4'hfae1;
         4'h4b92 	:	val_out <= 4'hfae1;
         4'h4b93 	:	val_out <= 4'hfae1;
         4'h4b98 	:	val_out <= 4'hfada;
         4'h4b99 	:	val_out <= 4'hfada;
         4'h4b9a 	:	val_out <= 4'hfada;
         4'h4b9b 	:	val_out <= 4'hfada;
         4'h4ba0 	:	val_out <= 4'hfad3;
         4'h4ba1 	:	val_out <= 4'hfad3;
         4'h4ba2 	:	val_out <= 4'hfad3;
         4'h4ba3 	:	val_out <= 4'hfad3;
         4'h4ba8 	:	val_out <= 4'hfacc;
         4'h4ba9 	:	val_out <= 4'hfacc;
         4'h4baa 	:	val_out <= 4'hfacc;
         4'h4bab 	:	val_out <= 4'hfacc;
         4'h4bb0 	:	val_out <= 4'hfac5;
         4'h4bb1 	:	val_out <= 4'hfac5;
         4'h4bb2 	:	val_out <= 4'hfac5;
         4'h4bb3 	:	val_out <= 4'hfac5;
         4'h4bb8 	:	val_out <= 4'hfabd;
         4'h4bb9 	:	val_out <= 4'hfabd;
         4'h4bba 	:	val_out <= 4'hfabd;
         4'h4bbb 	:	val_out <= 4'hfabd;
         4'h4bc0 	:	val_out <= 4'hfab6;
         4'h4bc1 	:	val_out <= 4'hfab6;
         4'h4bc2 	:	val_out <= 4'hfab6;
         4'h4bc3 	:	val_out <= 4'hfab6;
         4'h4bc8 	:	val_out <= 4'hfaaf;
         4'h4bc9 	:	val_out <= 4'hfaaf;
         4'h4bca 	:	val_out <= 4'hfaaf;
         4'h4bcb 	:	val_out <= 4'hfaaf;
         4'h4bd0 	:	val_out <= 4'hfaa8;
         4'h4bd1 	:	val_out <= 4'hfaa8;
         4'h4bd2 	:	val_out <= 4'hfaa8;
         4'h4bd3 	:	val_out <= 4'hfaa8;
         4'h4bd8 	:	val_out <= 4'hfaa1;
         4'h4bd9 	:	val_out <= 4'hfaa1;
         4'h4bda 	:	val_out <= 4'hfaa1;
         4'h4bdb 	:	val_out <= 4'hfaa1;
         4'h4be0 	:	val_out <= 4'hfa9a;
         4'h4be1 	:	val_out <= 4'hfa9a;
         4'h4be2 	:	val_out <= 4'hfa9a;
         4'h4be3 	:	val_out <= 4'hfa9a;
         4'h4be8 	:	val_out <= 4'hfa92;
         4'h4be9 	:	val_out <= 4'hfa92;
         4'h4bea 	:	val_out <= 4'hfa92;
         4'h4beb 	:	val_out <= 4'hfa92;
         4'h4bf0 	:	val_out <= 4'hfa8b;
         4'h4bf1 	:	val_out <= 4'hfa8b;
         4'h4bf2 	:	val_out <= 4'hfa8b;
         4'h4bf3 	:	val_out <= 4'hfa8b;
         4'h4bf8 	:	val_out <= 4'hfa84;
         4'h4bf9 	:	val_out <= 4'hfa84;
         4'h4bfa 	:	val_out <= 4'hfa84;
         4'h4bfb 	:	val_out <= 4'hfa84;
         4'h4c00 	:	val_out <= 4'hfa7d;
         4'h4c01 	:	val_out <= 4'hfa7d;
         4'h4c02 	:	val_out <= 4'hfa7d;
         4'h4c03 	:	val_out <= 4'hfa7d;
         4'h4c08 	:	val_out <= 4'hfa75;
         4'h4c09 	:	val_out <= 4'hfa75;
         4'h4c0a 	:	val_out <= 4'hfa75;
         4'h4c0b 	:	val_out <= 4'hfa75;
         4'h4c10 	:	val_out <= 4'hfa6e;
         4'h4c11 	:	val_out <= 4'hfa6e;
         4'h4c12 	:	val_out <= 4'hfa6e;
         4'h4c13 	:	val_out <= 4'hfa6e;
         4'h4c18 	:	val_out <= 4'hfa67;
         4'h4c19 	:	val_out <= 4'hfa67;
         4'h4c1a 	:	val_out <= 4'hfa67;
         4'h4c1b 	:	val_out <= 4'hfa67;
         4'h4c20 	:	val_out <= 4'hfa5f;
         4'h4c21 	:	val_out <= 4'hfa5f;
         4'h4c22 	:	val_out <= 4'hfa5f;
         4'h4c23 	:	val_out <= 4'hfa5f;
         4'h4c28 	:	val_out <= 4'hfa58;
         4'h4c29 	:	val_out <= 4'hfa58;
         4'h4c2a 	:	val_out <= 4'hfa58;
         4'h4c2b 	:	val_out <= 4'hfa58;
         4'h4c30 	:	val_out <= 4'hfa50;
         4'h4c31 	:	val_out <= 4'hfa50;
         4'h4c32 	:	val_out <= 4'hfa50;
         4'h4c33 	:	val_out <= 4'hfa50;
         4'h4c38 	:	val_out <= 4'hfa49;
         4'h4c39 	:	val_out <= 4'hfa49;
         4'h4c3a 	:	val_out <= 4'hfa49;
         4'h4c3b 	:	val_out <= 4'hfa49;
         4'h4c40 	:	val_out <= 4'hfa42;
         4'h4c41 	:	val_out <= 4'hfa42;
         4'h4c42 	:	val_out <= 4'hfa42;
         4'h4c43 	:	val_out <= 4'hfa42;
         4'h4c48 	:	val_out <= 4'hfa3a;
         4'h4c49 	:	val_out <= 4'hfa3a;
         4'h4c4a 	:	val_out <= 4'hfa3a;
         4'h4c4b 	:	val_out <= 4'hfa3a;
         4'h4c50 	:	val_out <= 4'hfa33;
         4'h4c51 	:	val_out <= 4'hfa33;
         4'h4c52 	:	val_out <= 4'hfa33;
         4'h4c53 	:	val_out <= 4'hfa33;
         4'h4c58 	:	val_out <= 4'hfa2b;
         4'h4c59 	:	val_out <= 4'hfa2b;
         4'h4c5a 	:	val_out <= 4'hfa2b;
         4'h4c5b 	:	val_out <= 4'hfa2b;
         4'h4c60 	:	val_out <= 4'hfa24;
         4'h4c61 	:	val_out <= 4'hfa24;
         4'h4c62 	:	val_out <= 4'hfa24;
         4'h4c63 	:	val_out <= 4'hfa24;
         4'h4c68 	:	val_out <= 4'hfa1c;
         4'h4c69 	:	val_out <= 4'hfa1c;
         4'h4c6a 	:	val_out <= 4'hfa1c;
         4'h4c6b 	:	val_out <= 4'hfa1c;
         4'h4c70 	:	val_out <= 4'hfa15;
         4'h4c71 	:	val_out <= 4'hfa15;
         4'h4c72 	:	val_out <= 4'hfa15;
         4'h4c73 	:	val_out <= 4'hfa15;
         4'h4c78 	:	val_out <= 4'hfa0d;
         4'h4c79 	:	val_out <= 4'hfa0d;
         4'h4c7a 	:	val_out <= 4'hfa0d;
         4'h4c7b 	:	val_out <= 4'hfa0d;
         4'h4c80 	:	val_out <= 4'hfa05;
         4'h4c81 	:	val_out <= 4'hfa05;
         4'h4c82 	:	val_out <= 4'hfa05;
         4'h4c83 	:	val_out <= 4'hfa05;
         4'h4c88 	:	val_out <= 4'hf9fe;
         4'h4c89 	:	val_out <= 4'hf9fe;
         4'h4c8a 	:	val_out <= 4'hf9fe;
         4'h4c8b 	:	val_out <= 4'hf9fe;
         4'h4c90 	:	val_out <= 4'hf9f6;
         4'h4c91 	:	val_out <= 4'hf9f6;
         4'h4c92 	:	val_out <= 4'hf9f6;
         4'h4c93 	:	val_out <= 4'hf9f6;
         4'h4c98 	:	val_out <= 4'hf9ef;
         4'h4c99 	:	val_out <= 4'hf9ef;
         4'h4c9a 	:	val_out <= 4'hf9ef;
         4'h4c9b 	:	val_out <= 4'hf9ef;
         4'h4ca0 	:	val_out <= 4'hf9e7;
         4'h4ca1 	:	val_out <= 4'hf9e7;
         4'h4ca2 	:	val_out <= 4'hf9e7;
         4'h4ca3 	:	val_out <= 4'hf9e7;
         4'h4ca8 	:	val_out <= 4'hf9df;
         4'h4ca9 	:	val_out <= 4'hf9df;
         4'h4caa 	:	val_out <= 4'hf9df;
         4'h4cab 	:	val_out <= 4'hf9df;
         4'h4cb0 	:	val_out <= 4'hf9d8;
         4'h4cb1 	:	val_out <= 4'hf9d8;
         4'h4cb2 	:	val_out <= 4'hf9d8;
         4'h4cb3 	:	val_out <= 4'hf9d8;
         4'h4cb8 	:	val_out <= 4'hf9d0;
         4'h4cb9 	:	val_out <= 4'hf9d0;
         4'h4cba 	:	val_out <= 4'hf9d0;
         4'h4cbb 	:	val_out <= 4'hf9d0;
         4'h4cc0 	:	val_out <= 4'hf9c8;
         4'h4cc1 	:	val_out <= 4'hf9c8;
         4'h4cc2 	:	val_out <= 4'hf9c8;
         4'h4cc3 	:	val_out <= 4'hf9c8;
         4'h4cc8 	:	val_out <= 4'hf9c0;
         4'h4cc9 	:	val_out <= 4'hf9c0;
         4'h4cca 	:	val_out <= 4'hf9c0;
         4'h4ccb 	:	val_out <= 4'hf9c0;
         4'h4cd0 	:	val_out <= 4'hf9b9;
         4'h4cd1 	:	val_out <= 4'hf9b9;
         4'h4cd2 	:	val_out <= 4'hf9b9;
         4'h4cd3 	:	val_out <= 4'hf9b9;
         4'h4cd8 	:	val_out <= 4'hf9b1;
         4'h4cd9 	:	val_out <= 4'hf9b1;
         4'h4cda 	:	val_out <= 4'hf9b1;
         4'h4cdb 	:	val_out <= 4'hf9b1;
         4'h4ce0 	:	val_out <= 4'hf9a9;
         4'h4ce1 	:	val_out <= 4'hf9a9;
         4'h4ce2 	:	val_out <= 4'hf9a9;
         4'h4ce3 	:	val_out <= 4'hf9a9;
         4'h4ce8 	:	val_out <= 4'hf9a1;
         4'h4ce9 	:	val_out <= 4'hf9a1;
         4'h4cea 	:	val_out <= 4'hf9a1;
         4'h4ceb 	:	val_out <= 4'hf9a1;
         4'h4cf0 	:	val_out <= 4'hf999;
         4'h4cf1 	:	val_out <= 4'hf999;
         4'h4cf2 	:	val_out <= 4'hf999;
         4'h4cf3 	:	val_out <= 4'hf999;
         4'h4cf8 	:	val_out <= 4'hf992;
         4'h4cf9 	:	val_out <= 4'hf992;
         4'h4cfa 	:	val_out <= 4'hf992;
         4'h4cfb 	:	val_out <= 4'hf992;
         4'h4d00 	:	val_out <= 4'hf98a;
         4'h4d01 	:	val_out <= 4'hf98a;
         4'h4d02 	:	val_out <= 4'hf98a;
         4'h4d03 	:	val_out <= 4'hf98a;
         4'h4d08 	:	val_out <= 4'hf982;
         4'h4d09 	:	val_out <= 4'hf982;
         4'h4d0a 	:	val_out <= 4'hf982;
         4'h4d0b 	:	val_out <= 4'hf982;
         4'h4d10 	:	val_out <= 4'hf97a;
         4'h4d11 	:	val_out <= 4'hf97a;
         4'h4d12 	:	val_out <= 4'hf97a;
         4'h4d13 	:	val_out <= 4'hf97a;
         4'h4d18 	:	val_out <= 4'hf972;
         4'h4d19 	:	val_out <= 4'hf972;
         4'h4d1a 	:	val_out <= 4'hf972;
         4'h4d1b 	:	val_out <= 4'hf972;
         4'h4d20 	:	val_out <= 4'hf96a;
         4'h4d21 	:	val_out <= 4'hf96a;
         4'h4d22 	:	val_out <= 4'hf96a;
         4'h4d23 	:	val_out <= 4'hf96a;
         4'h4d28 	:	val_out <= 4'hf962;
         4'h4d29 	:	val_out <= 4'hf962;
         4'h4d2a 	:	val_out <= 4'hf962;
         4'h4d2b 	:	val_out <= 4'hf962;
         4'h4d30 	:	val_out <= 4'hf95a;
         4'h4d31 	:	val_out <= 4'hf95a;
         4'h4d32 	:	val_out <= 4'hf95a;
         4'h4d33 	:	val_out <= 4'hf95a;
         4'h4d38 	:	val_out <= 4'hf952;
         4'h4d39 	:	val_out <= 4'hf952;
         4'h4d3a 	:	val_out <= 4'hf952;
         4'h4d3b 	:	val_out <= 4'hf952;
         4'h4d40 	:	val_out <= 4'hf94a;
         4'h4d41 	:	val_out <= 4'hf94a;
         4'h4d42 	:	val_out <= 4'hf94a;
         4'h4d43 	:	val_out <= 4'hf94a;
         4'h4d48 	:	val_out <= 4'hf942;
         4'h4d49 	:	val_out <= 4'hf942;
         4'h4d4a 	:	val_out <= 4'hf942;
         4'h4d4b 	:	val_out <= 4'hf942;
         4'h4d50 	:	val_out <= 4'hf93a;
         4'h4d51 	:	val_out <= 4'hf93a;
         4'h4d52 	:	val_out <= 4'hf93a;
         4'h4d53 	:	val_out <= 4'hf93a;
         4'h4d58 	:	val_out <= 4'hf932;
         4'h4d59 	:	val_out <= 4'hf932;
         4'h4d5a 	:	val_out <= 4'hf932;
         4'h4d5b 	:	val_out <= 4'hf932;
         4'h4d60 	:	val_out <= 4'hf92a;
         4'h4d61 	:	val_out <= 4'hf92a;
         4'h4d62 	:	val_out <= 4'hf92a;
         4'h4d63 	:	val_out <= 4'hf92a;
         4'h4d68 	:	val_out <= 4'hf922;
         4'h4d69 	:	val_out <= 4'hf922;
         4'h4d6a 	:	val_out <= 4'hf922;
         4'h4d6b 	:	val_out <= 4'hf922;
         4'h4d70 	:	val_out <= 4'hf919;
         4'h4d71 	:	val_out <= 4'hf919;
         4'h4d72 	:	val_out <= 4'hf919;
         4'h4d73 	:	val_out <= 4'hf919;
         4'h4d78 	:	val_out <= 4'hf911;
         4'h4d79 	:	val_out <= 4'hf911;
         4'h4d7a 	:	val_out <= 4'hf911;
         4'h4d7b 	:	val_out <= 4'hf911;
         4'h4d80 	:	val_out <= 4'hf909;
         4'h4d81 	:	val_out <= 4'hf909;
         4'h4d82 	:	val_out <= 4'hf909;
         4'h4d83 	:	val_out <= 4'hf909;
         4'h4d88 	:	val_out <= 4'hf901;
         4'h4d89 	:	val_out <= 4'hf901;
         4'h4d8a 	:	val_out <= 4'hf901;
         4'h4d8b 	:	val_out <= 4'hf901;
         4'h4d90 	:	val_out <= 4'hf8f9;
         4'h4d91 	:	val_out <= 4'hf8f9;
         4'h4d92 	:	val_out <= 4'hf8f9;
         4'h4d93 	:	val_out <= 4'hf8f9;
         4'h4d98 	:	val_out <= 4'hf8f1;
         4'h4d99 	:	val_out <= 4'hf8f1;
         4'h4d9a 	:	val_out <= 4'hf8f1;
         4'h4d9b 	:	val_out <= 4'hf8f1;
         4'h4da0 	:	val_out <= 4'hf8e8;
         4'h4da1 	:	val_out <= 4'hf8e8;
         4'h4da2 	:	val_out <= 4'hf8e8;
         4'h4da3 	:	val_out <= 4'hf8e8;
         4'h4da8 	:	val_out <= 4'hf8e0;
         4'h4da9 	:	val_out <= 4'hf8e0;
         4'h4daa 	:	val_out <= 4'hf8e0;
         4'h4dab 	:	val_out <= 4'hf8e0;
         4'h4db0 	:	val_out <= 4'hf8d8;
         4'h4db1 	:	val_out <= 4'hf8d8;
         4'h4db2 	:	val_out <= 4'hf8d8;
         4'h4db3 	:	val_out <= 4'hf8d8;
         4'h4db8 	:	val_out <= 4'hf8cf;
         4'h4db9 	:	val_out <= 4'hf8cf;
         4'h4dba 	:	val_out <= 4'hf8cf;
         4'h4dbb 	:	val_out <= 4'hf8cf;
         4'h4dc0 	:	val_out <= 4'hf8c7;
         4'h4dc1 	:	val_out <= 4'hf8c7;
         4'h4dc2 	:	val_out <= 4'hf8c7;
         4'h4dc3 	:	val_out <= 4'hf8c7;
         4'h4dc8 	:	val_out <= 4'hf8bf;
         4'h4dc9 	:	val_out <= 4'hf8bf;
         4'h4dca 	:	val_out <= 4'hf8bf;
         4'h4dcb 	:	val_out <= 4'hf8bf;
         4'h4dd0 	:	val_out <= 4'hf8b6;
         4'h4dd1 	:	val_out <= 4'hf8b6;
         4'h4dd2 	:	val_out <= 4'hf8b6;
         4'h4dd3 	:	val_out <= 4'hf8b6;
         4'h4dd8 	:	val_out <= 4'hf8ae;
         4'h4dd9 	:	val_out <= 4'hf8ae;
         4'h4dda 	:	val_out <= 4'hf8ae;
         4'h4ddb 	:	val_out <= 4'hf8ae;
         4'h4de0 	:	val_out <= 4'hf8a6;
         4'h4de1 	:	val_out <= 4'hf8a6;
         4'h4de2 	:	val_out <= 4'hf8a6;
         4'h4de3 	:	val_out <= 4'hf8a6;
         4'h4de8 	:	val_out <= 4'hf89d;
         4'h4de9 	:	val_out <= 4'hf89d;
         4'h4dea 	:	val_out <= 4'hf89d;
         4'h4deb 	:	val_out <= 4'hf89d;
         4'h4df0 	:	val_out <= 4'hf895;
         4'h4df1 	:	val_out <= 4'hf895;
         4'h4df2 	:	val_out <= 4'hf895;
         4'h4df3 	:	val_out <= 4'hf895;
         4'h4df8 	:	val_out <= 4'hf88c;
         4'h4df9 	:	val_out <= 4'hf88c;
         4'h4dfa 	:	val_out <= 4'hf88c;
         4'h4dfb 	:	val_out <= 4'hf88c;
         4'h4e00 	:	val_out <= 4'hf884;
         4'h4e01 	:	val_out <= 4'hf884;
         4'h4e02 	:	val_out <= 4'hf884;
         4'h4e03 	:	val_out <= 4'hf884;
         4'h4e08 	:	val_out <= 4'hf87c;
         4'h4e09 	:	val_out <= 4'hf87c;
         4'h4e0a 	:	val_out <= 4'hf87c;
         4'h4e0b 	:	val_out <= 4'hf87c;
         4'h4e10 	:	val_out <= 4'hf873;
         4'h4e11 	:	val_out <= 4'hf873;
         4'h4e12 	:	val_out <= 4'hf873;
         4'h4e13 	:	val_out <= 4'hf873;
         4'h4e18 	:	val_out <= 4'hf86b;
         4'h4e19 	:	val_out <= 4'hf86b;
         4'h4e1a 	:	val_out <= 4'hf86b;
         4'h4e1b 	:	val_out <= 4'hf86b;
         4'h4e20 	:	val_out <= 4'hf862;
         4'h4e21 	:	val_out <= 4'hf862;
         4'h4e22 	:	val_out <= 4'hf862;
         4'h4e23 	:	val_out <= 4'hf862;
         4'h4e28 	:	val_out <= 4'hf859;
         4'h4e29 	:	val_out <= 4'hf859;
         4'h4e2a 	:	val_out <= 4'hf859;
         4'h4e2b 	:	val_out <= 4'hf859;
         4'h4e30 	:	val_out <= 4'hf851;
         4'h4e31 	:	val_out <= 4'hf851;
         4'h4e32 	:	val_out <= 4'hf851;
         4'h4e33 	:	val_out <= 4'hf851;
         4'h4e38 	:	val_out <= 4'hf848;
         4'h4e39 	:	val_out <= 4'hf848;
         4'h4e3a 	:	val_out <= 4'hf848;
         4'h4e3b 	:	val_out <= 4'hf848;
         4'h4e40 	:	val_out <= 4'hf840;
         4'h4e41 	:	val_out <= 4'hf840;
         4'h4e42 	:	val_out <= 4'hf840;
         4'h4e43 	:	val_out <= 4'hf840;
         4'h4e48 	:	val_out <= 4'hf837;
         4'h4e49 	:	val_out <= 4'hf837;
         4'h4e4a 	:	val_out <= 4'hf837;
         4'h4e4b 	:	val_out <= 4'hf837;
         4'h4e50 	:	val_out <= 4'hf82e;
         4'h4e51 	:	val_out <= 4'hf82e;
         4'h4e52 	:	val_out <= 4'hf82e;
         4'h4e53 	:	val_out <= 4'hf82e;
         4'h4e58 	:	val_out <= 4'hf826;
         4'h4e59 	:	val_out <= 4'hf826;
         4'h4e5a 	:	val_out <= 4'hf826;
         4'h4e5b 	:	val_out <= 4'hf826;
         4'h4e60 	:	val_out <= 4'hf81d;
         4'h4e61 	:	val_out <= 4'hf81d;
         4'h4e62 	:	val_out <= 4'hf81d;
         4'h4e63 	:	val_out <= 4'hf81d;
         4'h4e68 	:	val_out <= 4'hf814;
         4'h4e69 	:	val_out <= 4'hf814;
         4'h4e6a 	:	val_out <= 4'hf814;
         4'h4e6b 	:	val_out <= 4'hf814;
         4'h4e70 	:	val_out <= 4'hf80c;
         4'h4e71 	:	val_out <= 4'hf80c;
         4'h4e72 	:	val_out <= 4'hf80c;
         4'h4e73 	:	val_out <= 4'hf80c;
         4'h4e78 	:	val_out <= 4'hf803;
         4'h4e79 	:	val_out <= 4'hf803;
         4'h4e7a 	:	val_out <= 4'hf803;
         4'h4e7b 	:	val_out <= 4'hf803;
         4'h4e80 	:	val_out <= 4'hf7fa;
         4'h4e81 	:	val_out <= 4'hf7fa;
         4'h4e82 	:	val_out <= 4'hf7fa;
         4'h4e83 	:	val_out <= 4'hf7fa;
         4'h4e88 	:	val_out <= 4'hf7f1;
         4'h4e89 	:	val_out <= 4'hf7f1;
         4'h4e8a 	:	val_out <= 4'hf7f1;
         4'h4e8b 	:	val_out <= 4'hf7f1;
         4'h4e90 	:	val_out <= 4'hf7e9;
         4'h4e91 	:	val_out <= 4'hf7e9;
         4'h4e92 	:	val_out <= 4'hf7e9;
         4'h4e93 	:	val_out <= 4'hf7e9;
         4'h4e98 	:	val_out <= 4'hf7e0;
         4'h4e99 	:	val_out <= 4'hf7e0;
         4'h4e9a 	:	val_out <= 4'hf7e0;
         4'h4e9b 	:	val_out <= 4'hf7e0;
         4'h4ea0 	:	val_out <= 4'hf7d7;
         4'h4ea1 	:	val_out <= 4'hf7d7;
         4'h4ea2 	:	val_out <= 4'hf7d7;
         4'h4ea3 	:	val_out <= 4'hf7d7;
         4'h4ea8 	:	val_out <= 4'hf7ce;
         4'h4ea9 	:	val_out <= 4'hf7ce;
         4'h4eaa 	:	val_out <= 4'hf7ce;
         4'h4eab 	:	val_out <= 4'hf7ce;
         4'h4eb0 	:	val_out <= 4'hf7c5;
         4'h4eb1 	:	val_out <= 4'hf7c5;
         4'h4eb2 	:	val_out <= 4'hf7c5;
         4'h4eb3 	:	val_out <= 4'hf7c5;
         4'h4eb8 	:	val_out <= 4'hf7bc;
         4'h4eb9 	:	val_out <= 4'hf7bc;
         4'h4eba 	:	val_out <= 4'hf7bc;
         4'h4ebb 	:	val_out <= 4'hf7bc;
         4'h4ec0 	:	val_out <= 4'hf7b4;
         4'h4ec1 	:	val_out <= 4'hf7b4;
         4'h4ec2 	:	val_out <= 4'hf7b4;
         4'h4ec3 	:	val_out <= 4'hf7b4;
         4'h4ec8 	:	val_out <= 4'hf7ab;
         4'h4ec9 	:	val_out <= 4'hf7ab;
         4'h4eca 	:	val_out <= 4'hf7ab;
         4'h4ecb 	:	val_out <= 4'hf7ab;
         4'h4ed0 	:	val_out <= 4'hf7a2;
         4'h4ed1 	:	val_out <= 4'hf7a2;
         4'h4ed2 	:	val_out <= 4'hf7a2;
         4'h4ed3 	:	val_out <= 4'hf7a2;
         4'h4ed8 	:	val_out <= 4'hf799;
         4'h4ed9 	:	val_out <= 4'hf799;
         4'h4eda 	:	val_out <= 4'hf799;
         4'h4edb 	:	val_out <= 4'hf799;
         4'h4ee0 	:	val_out <= 4'hf790;
         4'h4ee1 	:	val_out <= 4'hf790;
         4'h4ee2 	:	val_out <= 4'hf790;
         4'h4ee3 	:	val_out <= 4'hf790;
         4'h4ee8 	:	val_out <= 4'hf787;
         4'h4ee9 	:	val_out <= 4'hf787;
         4'h4eea 	:	val_out <= 4'hf787;
         4'h4eeb 	:	val_out <= 4'hf787;
         4'h4ef0 	:	val_out <= 4'hf77e;
         4'h4ef1 	:	val_out <= 4'hf77e;
         4'h4ef2 	:	val_out <= 4'hf77e;
         4'h4ef3 	:	val_out <= 4'hf77e;
         4'h4ef8 	:	val_out <= 4'hf775;
         4'h4ef9 	:	val_out <= 4'hf775;
         4'h4efa 	:	val_out <= 4'hf775;
         4'h4efb 	:	val_out <= 4'hf775;
         4'h4f00 	:	val_out <= 4'hf76c;
         4'h4f01 	:	val_out <= 4'hf76c;
         4'h4f02 	:	val_out <= 4'hf76c;
         4'h4f03 	:	val_out <= 4'hf76c;
         4'h4f08 	:	val_out <= 4'hf763;
         4'h4f09 	:	val_out <= 4'hf763;
         4'h4f0a 	:	val_out <= 4'hf763;
         4'h4f0b 	:	val_out <= 4'hf763;
         4'h4f10 	:	val_out <= 4'hf75a;
         4'h4f11 	:	val_out <= 4'hf75a;
         4'h4f12 	:	val_out <= 4'hf75a;
         4'h4f13 	:	val_out <= 4'hf75a;
         4'h4f18 	:	val_out <= 4'hf751;
         4'h4f19 	:	val_out <= 4'hf751;
         4'h4f1a 	:	val_out <= 4'hf751;
         4'h4f1b 	:	val_out <= 4'hf751;
         4'h4f20 	:	val_out <= 4'hf747;
         4'h4f21 	:	val_out <= 4'hf747;
         4'h4f22 	:	val_out <= 4'hf747;
         4'h4f23 	:	val_out <= 4'hf747;
         4'h4f28 	:	val_out <= 4'hf73e;
         4'h4f29 	:	val_out <= 4'hf73e;
         4'h4f2a 	:	val_out <= 4'hf73e;
         4'h4f2b 	:	val_out <= 4'hf73e;
         4'h4f30 	:	val_out <= 4'hf735;
         4'h4f31 	:	val_out <= 4'hf735;
         4'h4f32 	:	val_out <= 4'hf735;
         4'h4f33 	:	val_out <= 4'hf735;
         4'h4f38 	:	val_out <= 4'hf72c;
         4'h4f39 	:	val_out <= 4'hf72c;
         4'h4f3a 	:	val_out <= 4'hf72c;
         4'h4f3b 	:	val_out <= 4'hf72c;
         4'h4f40 	:	val_out <= 4'hf723;
         4'h4f41 	:	val_out <= 4'hf723;
         4'h4f42 	:	val_out <= 4'hf723;
         4'h4f43 	:	val_out <= 4'hf723;
         4'h4f48 	:	val_out <= 4'hf71a;
         4'h4f49 	:	val_out <= 4'hf71a;
         4'h4f4a 	:	val_out <= 4'hf71a;
         4'h4f4b 	:	val_out <= 4'hf71a;
         4'h4f50 	:	val_out <= 4'hf710;
         4'h4f51 	:	val_out <= 4'hf710;
         4'h4f52 	:	val_out <= 4'hf710;
         4'h4f53 	:	val_out <= 4'hf710;
         4'h4f58 	:	val_out <= 4'hf707;
         4'h4f59 	:	val_out <= 4'hf707;
         4'h4f5a 	:	val_out <= 4'hf707;
         4'h4f5b 	:	val_out <= 4'hf707;
         4'h4f60 	:	val_out <= 4'hf6fe;
         4'h4f61 	:	val_out <= 4'hf6fe;
         4'h4f62 	:	val_out <= 4'hf6fe;
         4'h4f63 	:	val_out <= 4'hf6fe;
         4'h4f68 	:	val_out <= 4'hf6f5;
         4'h4f69 	:	val_out <= 4'hf6f5;
         4'h4f6a 	:	val_out <= 4'hf6f5;
         4'h4f6b 	:	val_out <= 4'hf6f5;
         4'h4f70 	:	val_out <= 4'hf6eb;
         4'h4f71 	:	val_out <= 4'hf6eb;
         4'h4f72 	:	val_out <= 4'hf6eb;
         4'h4f73 	:	val_out <= 4'hf6eb;
         4'h4f78 	:	val_out <= 4'hf6e2;
         4'h4f79 	:	val_out <= 4'hf6e2;
         4'h4f7a 	:	val_out <= 4'hf6e2;
         4'h4f7b 	:	val_out <= 4'hf6e2;
         4'h4f80 	:	val_out <= 4'hf6d9;
         4'h4f81 	:	val_out <= 4'hf6d9;
         4'h4f82 	:	val_out <= 4'hf6d9;
         4'h4f83 	:	val_out <= 4'hf6d9;
         4'h4f88 	:	val_out <= 4'hf6cf;
         4'h4f89 	:	val_out <= 4'hf6cf;
         4'h4f8a 	:	val_out <= 4'hf6cf;
         4'h4f8b 	:	val_out <= 4'hf6cf;
         4'h4f90 	:	val_out <= 4'hf6c6;
         4'h4f91 	:	val_out <= 4'hf6c6;
         4'h4f92 	:	val_out <= 4'hf6c6;
         4'h4f93 	:	val_out <= 4'hf6c6;
         4'h4f98 	:	val_out <= 4'hf6bd;
         4'h4f99 	:	val_out <= 4'hf6bd;
         4'h4f9a 	:	val_out <= 4'hf6bd;
         4'h4f9b 	:	val_out <= 4'hf6bd;
         4'h4fa0 	:	val_out <= 4'hf6b3;
         4'h4fa1 	:	val_out <= 4'hf6b3;
         4'h4fa2 	:	val_out <= 4'hf6b3;
         4'h4fa3 	:	val_out <= 4'hf6b3;
         4'h4fa8 	:	val_out <= 4'hf6aa;
         4'h4fa9 	:	val_out <= 4'hf6aa;
         4'h4faa 	:	val_out <= 4'hf6aa;
         4'h4fab 	:	val_out <= 4'hf6aa;
         4'h4fb0 	:	val_out <= 4'hf6a0;
         4'h4fb1 	:	val_out <= 4'hf6a0;
         4'h4fb2 	:	val_out <= 4'hf6a0;
         4'h4fb3 	:	val_out <= 4'hf6a0;
         4'h4fb8 	:	val_out <= 4'hf697;
         4'h4fb9 	:	val_out <= 4'hf697;
         4'h4fba 	:	val_out <= 4'hf697;
         4'h4fbb 	:	val_out <= 4'hf697;
         4'h4fc0 	:	val_out <= 4'hf68e;
         4'h4fc1 	:	val_out <= 4'hf68e;
         4'h4fc2 	:	val_out <= 4'hf68e;
         4'h4fc3 	:	val_out <= 4'hf68e;
         4'h4fc8 	:	val_out <= 4'hf684;
         4'h4fc9 	:	val_out <= 4'hf684;
         4'h4fca 	:	val_out <= 4'hf684;
         4'h4fcb 	:	val_out <= 4'hf684;
         4'h4fd0 	:	val_out <= 4'hf67b;
         4'h4fd1 	:	val_out <= 4'hf67b;
         4'h4fd2 	:	val_out <= 4'hf67b;
         4'h4fd3 	:	val_out <= 4'hf67b;
         4'h4fd8 	:	val_out <= 4'hf671;
         4'h4fd9 	:	val_out <= 4'hf671;
         4'h4fda 	:	val_out <= 4'hf671;
         4'h4fdb 	:	val_out <= 4'hf671;
         4'h4fe0 	:	val_out <= 4'hf668;
         4'h4fe1 	:	val_out <= 4'hf668;
         4'h4fe2 	:	val_out <= 4'hf668;
         4'h4fe3 	:	val_out <= 4'hf668;
         4'h4fe8 	:	val_out <= 4'hf65e;
         4'h4fe9 	:	val_out <= 4'hf65e;
         4'h4fea 	:	val_out <= 4'hf65e;
         4'h4feb 	:	val_out <= 4'hf65e;
         4'h4ff0 	:	val_out <= 4'hf654;
         4'h4ff1 	:	val_out <= 4'hf654;
         4'h4ff2 	:	val_out <= 4'hf654;
         4'h4ff3 	:	val_out <= 4'hf654;
         4'h4ff8 	:	val_out <= 4'hf64b;
         4'h4ff9 	:	val_out <= 4'hf64b;
         4'h4ffa 	:	val_out <= 4'hf64b;
         4'h4ffb 	:	val_out <= 4'hf64b;
         4'h5000 	:	val_out <= 4'hf641;
         4'h5001 	:	val_out <= 4'hf641;
         4'h5002 	:	val_out <= 4'hf641;
         4'h5003 	:	val_out <= 4'hf641;
         4'h5008 	:	val_out <= 4'hf638;
         4'h5009 	:	val_out <= 4'hf638;
         4'h500a 	:	val_out <= 4'hf638;
         4'h500b 	:	val_out <= 4'hf638;
         4'h5010 	:	val_out <= 4'hf62e;
         4'h5011 	:	val_out <= 4'hf62e;
         4'h5012 	:	val_out <= 4'hf62e;
         4'h5013 	:	val_out <= 4'hf62e;
         4'h5018 	:	val_out <= 4'hf624;
         4'h5019 	:	val_out <= 4'hf624;
         4'h501a 	:	val_out <= 4'hf624;
         4'h501b 	:	val_out <= 4'hf624;
         4'h5020 	:	val_out <= 4'hf61b;
         4'h5021 	:	val_out <= 4'hf61b;
         4'h5022 	:	val_out <= 4'hf61b;
         4'h5023 	:	val_out <= 4'hf61b;
         4'h5028 	:	val_out <= 4'hf611;
         4'h5029 	:	val_out <= 4'hf611;
         4'h502a 	:	val_out <= 4'hf611;
         4'h502b 	:	val_out <= 4'hf611;
         4'h5030 	:	val_out <= 4'hf607;
         4'h5031 	:	val_out <= 4'hf607;
         4'h5032 	:	val_out <= 4'hf607;
         4'h5033 	:	val_out <= 4'hf607;
         4'h5038 	:	val_out <= 4'hf5fd;
         4'h5039 	:	val_out <= 4'hf5fd;
         4'h503a 	:	val_out <= 4'hf5fd;
         4'h503b 	:	val_out <= 4'hf5fd;
         4'h5040 	:	val_out <= 4'hf5f4;
         4'h5041 	:	val_out <= 4'hf5f4;
         4'h5042 	:	val_out <= 4'hf5f4;
         4'h5043 	:	val_out <= 4'hf5f4;
         4'h5048 	:	val_out <= 4'hf5ea;
         4'h5049 	:	val_out <= 4'hf5ea;
         4'h504a 	:	val_out <= 4'hf5ea;
         4'h504b 	:	val_out <= 4'hf5ea;
         4'h5050 	:	val_out <= 4'hf5e0;
         4'h5051 	:	val_out <= 4'hf5e0;
         4'h5052 	:	val_out <= 4'hf5e0;
         4'h5053 	:	val_out <= 4'hf5e0;
         4'h5058 	:	val_out <= 4'hf5d6;
         4'h5059 	:	val_out <= 4'hf5d6;
         4'h505a 	:	val_out <= 4'hf5d6;
         4'h505b 	:	val_out <= 4'hf5d6;
         4'h5060 	:	val_out <= 4'hf5cc;
         4'h5061 	:	val_out <= 4'hf5cc;
         4'h5062 	:	val_out <= 4'hf5cc;
         4'h5063 	:	val_out <= 4'hf5cc;
         4'h5068 	:	val_out <= 4'hf5c3;
         4'h5069 	:	val_out <= 4'hf5c3;
         4'h506a 	:	val_out <= 4'hf5c3;
         4'h506b 	:	val_out <= 4'hf5c3;
         4'h5070 	:	val_out <= 4'hf5b9;
         4'h5071 	:	val_out <= 4'hf5b9;
         4'h5072 	:	val_out <= 4'hf5b9;
         4'h5073 	:	val_out <= 4'hf5b9;
         4'h5078 	:	val_out <= 4'hf5af;
         4'h5079 	:	val_out <= 4'hf5af;
         4'h507a 	:	val_out <= 4'hf5af;
         4'h507b 	:	val_out <= 4'hf5af;
         4'h5080 	:	val_out <= 4'hf5a5;
         4'h5081 	:	val_out <= 4'hf5a5;
         4'h5082 	:	val_out <= 4'hf5a5;
         4'h5083 	:	val_out <= 4'hf5a5;
         4'h5088 	:	val_out <= 4'hf59b;
         4'h5089 	:	val_out <= 4'hf59b;
         4'h508a 	:	val_out <= 4'hf59b;
         4'h508b 	:	val_out <= 4'hf59b;
         4'h5090 	:	val_out <= 4'hf591;
         4'h5091 	:	val_out <= 4'hf591;
         4'h5092 	:	val_out <= 4'hf591;
         4'h5093 	:	val_out <= 4'hf591;
         4'h5098 	:	val_out <= 4'hf587;
         4'h5099 	:	val_out <= 4'hf587;
         4'h509a 	:	val_out <= 4'hf587;
         4'h509b 	:	val_out <= 4'hf587;
         4'h50a0 	:	val_out <= 4'hf57d;
         4'h50a1 	:	val_out <= 4'hf57d;
         4'h50a2 	:	val_out <= 4'hf57d;
         4'h50a3 	:	val_out <= 4'hf57d;
         4'h50a8 	:	val_out <= 4'hf573;
         4'h50a9 	:	val_out <= 4'hf573;
         4'h50aa 	:	val_out <= 4'hf573;
         4'h50ab 	:	val_out <= 4'hf573;
         4'h50b0 	:	val_out <= 4'hf569;
         4'h50b1 	:	val_out <= 4'hf569;
         4'h50b2 	:	val_out <= 4'hf569;
         4'h50b3 	:	val_out <= 4'hf569;
         4'h50b8 	:	val_out <= 4'hf55f;
         4'h50b9 	:	val_out <= 4'hf55f;
         4'h50ba 	:	val_out <= 4'hf55f;
         4'h50bb 	:	val_out <= 4'hf55f;
         4'h50c0 	:	val_out <= 4'hf555;
         4'h50c1 	:	val_out <= 4'hf555;
         4'h50c2 	:	val_out <= 4'hf555;
         4'h50c3 	:	val_out <= 4'hf555;
         4'h50c8 	:	val_out <= 4'hf54b;
         4'h50c9 	:	val_out <= 4'hf54b;
         4'h50ca 	:	val_out <= 4'hf54b;
         4'h50cb 	:	val_out <= 4'hf54b;
         4'h50d0 	:	val_out <= 4'hf541;
         4'h50d1 	:	val_out <= 4'hf541;
         4'h50d2 	:	val_out <= 4'hf541;
         4'h50d3 	:	val_out <= 4'hf541;
         4'h50d8 	:	val_out <= 4'hf537;
         4'h50d9 	:	val_out <= 4'hf537;
         4'h50da 	:	val_out <= 4'hf537;
         4'h50db 	:	val_out <= 4'hf537;
         4'h50e0 	:	val_out <= 4'hf52d;
         4'h50e1 	:	val_out <= 4'hf52d;
         4'h50e2 	:	val_out <= 4'hf52d;
         4'h50e3 	:	val_out <= 4'hf52d;
         4'h50e8 	:	val_out <= 4'hf523;
         4'h50e9 	:	val_out <= 4'hf523;
         4'h50ea 	:	val_out <= 4'hf523;
         4'h50eb 	:	val_out <= 4'hf523;
         4'h50f0 	:	val_out <= 4'hf519;
         4'h50f1 	:	val_out <= 4'hf519;
         4'h50f2 	:	val_out <= 4'hf519;
         4'h50f3 	:	val_out <= 4'hf519;
         4'h50f8 	:	val_out <= 4'hf50f;
         4'h50f9 	:	val_out <= 4'hf50f;
         4'h50fa 	:	val_out <= 4'hf50f;
         4'h50fb 	:	val_out <= 4'hf50f;
         4'h5100 	:	val_out <= 4'hf504;
         4'h5101 	:	val_out <= 4'hf504;
         4'h5102 	:	val_out <= 4'hf504;
         4'h5103 	:	val_out <= 4'hf504;
         4'h5108 	:	val_out <= 4'hf4fa;
         4'h5109 	:	val_out <= 4'hf4fa;
         4'h510a 	:	val_out <= 4'hf4fa;
         4'h510b 	:	val_out <= 4'hf4fa;
         4'h5110 	:	val_out <= 4'hf4f0;
         4'h5111 	:	val_out <= 4'hf4f0;
         4'h5112 	:	val_out <= 4'hf4f0;
         4'h5113 	:	val_out <= 4'hf4f0;
         4'h5118 	:	val_out <= 4'hf4e6;
         4'h5119 	:	val_out <= 4'hf4e6;
         4'h511a 	:	val_out <= 4'hf4e6;
         4'h511b 	:	val_out <= 4'hf4e6;
         4'h5120 	:	val_out <= 4'hf4db;
         4'h5121 	:	val_out <= 4'hf4db;
         4'h5122 	:	val_out <= 4'hf4db;
         4'h5123 	:	val_out <= 4'hf4db;
         4'h5128 	:	val_out <= 4'hf4d1;
         4'h5129 	:	val_out <= 4'hf4d1;
         4'h512a 	:	val_out <= 4'hf4d1;
         4'h512b 	:	val_out <= 4'hf4d1;
         4'h5130 	:	val_out <= 4'hf4c7;
         4'h5131 	:	val_out <= 4'hf4c7;
         4'h5132 	:	val_out <= 4'hf4c7;
         4'h5133 	:	val_out <= 4'hf4c7;
         4'h5138 	:	val_out <= 4'hf4bd;
         4'h5139 	:	val_out <= 4'hf4bd;
         4'h513a 	:	val_out <= 4'hf4bd;
         4'h513b 	:	val_out <= 4'hf4bd;
         4'h5140 	:	val_out <= 4'hf4b2;
         4'h5141 	:	val_out <= 4'hf4b2;
         4'h5142 	:	val_out <= 4'hf4b2;
         4'h5143 	:	val_out <= 4'hf4b2;
         4'h5148 	:	val_out <= 4'hf4a8;
         4'h5149 	:	val_out <= 4'hf4a8;
         4'h514a 	:	val_out <= 4'hf4a8;
         4'h514b 	:	val_out <= 4'hf4a8;
         4'h5150 	:	val_out <= 4'hf49e;
         4'h5151 	:	val_out <= 4'hf49e;
         4'h5152 	:	val_out <= 4'hf49e;
         4'h5153 	:	val_out <= 4'hf49e;
         4'h5158 	:	val_out <= 4'hf493;
         4'h5159 	:	val_out <= 4'hf493;
         4'h515a 	:	val_out <= 4'hf493;
         4'h515b 	:	val_out <= 4'hf493;
         4'h5160 	:	val_out <= 4'hf489;
         4'h5161 	:	val_out <= 4'hf489;
         4'h5162 	:	val_out <= 4'hf489;
         4'h5163 	:	val_out <= 4'hf489;
         4'h5168 	:	val_out <= 4'hf47e;
         4'h5169 	:	val_out <= 4'hf47e;
         4'h516a 	:	val_out <= 4'hf47e;
         4'h516b 	:	val_out <= 4'hf47e;
         4'h5170 	:	val_out <= 4'hf474;
         4'h5171 	:	val_out <= 4'hf474;
         4'h5172 	:	val_out <= 4'hf474;
         4'h5173 	:	val_out <= 4'hf474;
         4'h5178 	:	val_out <= 4'hf46a;
         4'h5179 	:	val_out <= 4'hf46a;
         4'h517a 	:	val_out <= 4'hf46a;
         4'h517b 	:	val_out <= 4'hf46a;
         4'h5180 	:	val_out <= 4'hf45f;
         4'h5181 	:	val_out <= 4'hf45f;
         4'h5182 	:	val_out <= 4'hf45f;
         4'h5183 	:	val_out <= 4'hf45f;
         4'h5188 	:	val_out <= 4'hf455;
         4'h5189 	:	val_out <= 4'hf455;
         4'h518a 	:	val_out <= 4'hf455;
         4'h518b 	:	val_out <= 4'hf455;
         4'h5190 	:	val_out <= 4'hf44a;
         4'h5191 	:	val_out <= 4'hf44a;
         4'h5192 	:	val_out <= 4'hf44a;
         4'h5193 	:	val_out <= 4'hf44a;
         4'h5198 	:	val_out <= 4'hf440;
         4'h5199 	:	val_out <= 4'hf440;
         4'h519a 	:	val_out <= 4'hf440;
         4'h519b 	:	val_out <= 4'hf440;
         4'h51a0 	:	val_out <= 4'hf435;
         4'h51a1 	:	val_out <= 4'hf435;
         4'h51a2 	:	val_out <= 4'hf435;
         4'h51a3 	:	val_out <= 4'hf435;
         4'h51a8 	:	val_out <= 4'hf42b;
         4'h51a9 	:	val_out <= 4'hf42b;
         4'h51aa 	:	val_out <= 4'hf42b;
         4'h51ab 	:	val_out <= 4'hf42b;
         4'h51b0 	:	val_out <= 4'hf420;
         4'h51b1 	:	val_out <= 4'hf420;
         4'h51b2 	:	val_out <= 4'hf420;
         4'h51b3 	:	val_out <= 4'hf420;
         4'h51b8 	:	val_out <= 4'hf415;
         4'h51b9 	:	val_out <= 4'hf415;
         4'h51ba 	:	val_out <= 4'hf415;
         4'h51bb 	:	val_out <= 4'hf415;
         4'h51c0 	:	val_out <= 4'hf40b;
         4'h51c1 	:	val_out <= 4'hf40b;
         4'h51c2 	:	val_out <= 4'hf40b;
         4'h51c3 	:	val_out <= 4'hf40b;
         4'h51c8 	:	val_out <= 4'hf400;
         4'h51c9 	:	val_out <= 4'hf400;
         4'h51ca 	:	val_out <= 4'hf400;
         4'h51cb 	:	val_out <= 4'hf400;
         4'h51d0 	:	val_out <= 4'hf3f6;
         4'h51d1 	:	val_out <= 4'hf3f6;
         4'h51d2 	:	val_out <= 4'hf3f6;
         4'h51d3 	:	val_out <= 4'hf3f6;
         4'h51d8 	:	val_out <= 4'hf3eb;
         4'h51d9 	:	val_out <= 4'hf3eb;
         4'h51da 	:	val_out <= 4'hf3eb;
         4'h51db 	:	val_out <= 4'hf3eb;
         4'h51e0 	:	val_out <= 4'hf3e0;
         4'h51e1 	:	val_out <= 4'hf3e0;
         4'h51e2 	:	val_out <= 4'hf3e0;
         4'h51e3 	:	val_out <= 4'hf3e0;
         4'h51e8 	:	val_out <= 4'hf3d6;
         4'h51e9 	:	val_out <= 4'hf3d6;
         4'h51ea 	:	val_out <= 4'hf3d6;
         4'h51eb 	:	val_out <= 4'hf3d6;
         4'h51f0 	:	val_out <= 4'hf3cb;
         4'h51f1 	:	val_out <= 4'hf3cb;
         4'h51f2 	:	val_out <= 4'hf3cb;
         4'h51f3 	:	val_out <= 4'hf3cb;
         4'h51f8 	:	val_out <= 4'hf3c0;
         4'h51f9 	:	val_out <= 4'hf3c0;
         4'h51fa 	:	val_out <= 4'hf3c0;
         4'h51fb 	:	val_out <= 4'hf3c0;
         4'h5200 	:	val_out <= 4'hf3b5;
         4'h5201 	:	val_out <= 4'hf3b5;
         4'h5202 	:	val_out <= 4'hf3b5;
         4'h5203 	:	val_out <= 4'hf3b5;
         4'h5208 	:	val_out <= 4'hf3ab;
         4'h5209 	:	val_out <= 4'hf3ab;
         4'h520a 	:	val_out <= 4'hf3ab;
         4'h520b 	:	val_out <= 4'hf3ab;
         4'h5210 	:	val_out <= 4'hf3a0;
         4'h5211 	:	val_out <= 4'hf3a0;
         4'h5212 	:	val_out <= 4'hf3a0;
         4'h5213 	:	val_out <= 4'hf3a0;
         4'h5218 	:	val_out <= 4'hf395;
         4'h5219 	:	val_out <= 4'hf395;
         4'h521a 	:	val_out <= 4'hf395;
         4'h521b 	:	val_out <= 4'hf395;
         4'h5220 	:	val_out <= 4'hf38a;
         4'h5221 	:	val_out <= 4'hf38a;
         4'h5222 	:	val_out <= 4'hf38a;
         4'h5223 	:	val_out <= 4'hf38a;
         4'h5228 	:	val_out <= 4'hf37f;
         4'h5229 	:	val_out <= 4'hf37f;
         4'h522a 	:	val_out <= 4'hf37f;
         4'h522b 	:	val_out <= 4'hf37f;
         4'h5230 	:	val_out <= 4'hf375;
         4'h5231 	:	val_out <= 4'hf375;
         4'h5232 	:	val_out <= 4'hf375;
         4'h5233 	:	val_out <= 4'hf375;
         4'h5238 	:	val_out <= 4'hf36a;
         4'h5239 	:	val_out <= 4'hf36a;
         4'h523a 	:	val_out <= 4'hf36a;
         4'h523b 	:	val_out <= 4'hf36a;
         4'h5240 	:	val_out <= 4'hf35f;
         4'h5241 	:	val_out <= 4'hf35f;
         4'h5242 	:	val_out <= 4'hf35f;
         4'h5243 	:	val_out <= 4'hf35f;
         4'h5248 	:	val_out <= 4'hf354;
         4'h5249 	:	val_out <= 4'hf354;
         4'h524a 	:	val_out <= 4'hf354;
         4'h524b 	:	val_out <= 4'hf354;
         4'h5250 	:	val_out <= 4'hf349;
         4'h5251 	:	val_out <= 4'hf349;
         4'h5252 	:	val_out <= 4'hf349;
         4'h5253 	:	val_out <= 4'hf349;
         4'h5258 	:	val_out <= 4'hf33e;
         4'h5259 	:	val_out <= 4'hf33e;
         4'h525a 	:	val_out <= 4'hf33e;
         4'h525b 	:	val_out <= 4'hf33e;
         4'h5260 	:	val_out <= 4'hf333;
         4'h5261 	:	val_out <= 4'hf333;
         4'h5262 	:	val_out <= 4'hf333;
         4'h5263 	:	val_out <= 4'hf333;
         4'h5268 	:	val_out <= 4'hf328;
         4'h5269 	:	val_out <= 4'hf328;
         4'h526a 	:	val_out <= 4'hf328;
         4'h526b 	:	val_out <= 4'hf328;
         4'h5270 	:	val_out <= 4'hf31d;
         4'h5271 	:	val_out <= 4'hf31d;
         4'h5272 	:	val_out <= 4'hf31d;
         4'h5273 	:	val_out <= 4'hf31d;
         4'h5278 	:	val_out <= 4'hf312;
         4'h5279 	:	val_out <= 4'hf312;
         4'h527a 	:	val_out <= 4'hf312;
         4'h527b 	:	val_out <= 4'hf312;
         4'h5280 	:	val_out <= 4'hf307;
         4'h5281 	:	val_out <= 4'hf307;
         4'h5282 	:	val_out <= 4'hf307;
         4'h5283 	:	val_out <= 4'hf307;
         4'h5288 	:	val_out <= 4'hf2fc;
         4'h5289 	:	val_out <= 4'hf2fc;
         4'h528a 	:	val_out <= 4'hf2fc;
         4'h528b 	:	val_out <= 4'hf2fc;
         4'h5290 	:	val_out <= 4'hf2f1;
         4'h5291 	:	val_out <= 4'hf2f1;
         4'h5292 	:	val_out <= 4'hf2f1;
         4'h5293 	:	val_out <= 4'hf2f1;
         4'h5298 	:	val_out <= 4'hf2e6;
         4'h5299 	:	val_out <= 4'hf2e6;
         4'h529a 	:	val_out <= 4'hf2e6;
         4'h529b 	:	val_out <= 4'hf2e6;
         4'h52a0 	:	val_out <= 4'hf2db;
         4'h52a1 	:	val_out <= 4'hf2db;
         4'h52a2 	:	val_out <= 4'hf2db;
         4'h52a3 	:	val_out <= 4'hf2db;
         4'h52a8 	:	val_out <= 4'hf2d0;
         4'h52a9 	:	val_out <= 4'hf2d0;
         4'h52aa 	:	val_out <= 4'hf2d0;
         4'h52ab 	:	val_out <= 4'hf2d0;
         4'h52b0 	:	val_out <= 4'hf2c5;
         4'h52b1 	:	val_out <= 4'hf2c5;
         4'h52b2 	:	val_out <= 4'hf2c5;
         4'h52b3 	:	val_out <= 4'hf2c5;
         4'h52b8 	:	val_out <= 4'hf2ba;
         4'h52b9 	:	val_out <= 4'hf2ba;
         4'h52ba 	:	val_out <= 4'hf2ba;
         4'h52bb 	:	val_out <= 4'hf2ba;
         4'h52c0 	:	val_out <= 4'hf2af;
         4'h52c1 	:	val_out <= 4'hf2af;
         4'h52c2 	:	val_out <= 4'hf2af;
         4'h52c3 	:	val_out <= 4'hf2af;
         4'h52c8 	:	val_out <= 4'hf2a3;
         4'h52c9 	:	val_out <= 4'hf2a3;
         4'h52ca 	:	val_out <= 4'hf2a3;
         4'h52cb 	:	val_out <= 4'hf2a3;
         4'h52d0 	:	val_out <= 4'hf298;
         4'h52d1 	:	val_out <= 4'hf298;
         4'h52d2 	:	val_out <= 4'hf298;
         4'h52d3 	:	val_out <= 4'hf298;
         4'h52d8 	:	val_out <= 4'hf28d;
         4'h52d9 	:	val_out <= 4'hf28d;
         4'h52da 	:	val_out <= 4'hf28d;
         4'h52db 	:	val_out <= 4'hf28d;
         4'h52e0 	:	val_out <= 4'hf282;
         4'h52e1 	:	val_out <= 4'hf282;
         4'h52e2 	:	val_out <= 4'hf282;
         4'h52e3 	:	val_out <= 4'hf282;
         4'h52e8 	:	val_out <= 4'hf276;
         4'h52e9 	:	val_out <= 4'hf276;
         4'h52ea 	:	val_out <= 4'hf276;
         4'h52eb 	:	val_out <= 4'hf276;
         4'h52f0 	:	val_out <= 4'hf26b;
         4'h52f1 	:	val_out <= 4'hf26b;
         4'h52f2 	:	val_out <= 4'hf26b;
         4'h52f3 	:	val_out <= 4'hf26b;
         4'h52f8 	:	val_out <= 4'hf260;
         4'h52f9 	:	val_out <= 4'hf260;
         4'h52fa 	:	val_out <= 4'hf260;
         4'h52fb 	:	val_out <= 4'hf260;
         4'h5300 	:	val_out <= 4'hf255;
         4'h5301 	:	val_out <= 4'hf255;
         4'h5302 	:	val_out <= 4'hf255;
         4'h5303 	:	val_out <= 4'hf255;
         4'h5308 	:	val_out <= 4'hf249;
         4'h5309 	:	val_out <= 4'hf249;
         4'h530a 	:	val_out <= 4'hf249;
         4'h530b 	:	val_out <= 4'hf249;
         4'h5310 	:	val_out <= 4'hf23e;
         4'h5311 	:	val_out <= 4'hf23e;
         4'h5312 	:	val_out <= 4'hf23e;
         4'h5313 	:	val_out <= 4'hf23e;
         4'h5318 	:	val_out <= 4'hf233;
         4'h5319 	:	val_out <= 4'hf233;
         4'h531a 	:	val_out <= 4'hf233;
         4'h531b 	:	val_out <= 4'hf233;
         4'h5320 	:	val_out <= 4'hf227;
         4'h5321 	:	val_out <= 4'hf227;
         4'h5322 	:	val_out <= 4'hf227;
         4'h5323 	:	val_out <= 4'hf227;
         4'h5328 	:	val_out <= 4'hf21c;
         4'h5329 	:	val_out <= 4'hf21c;
         4'h532a 	:	val_out <= 4'hf21c;
         4'h532b 	:	val_out <= 4'hf21c;
         4'h5330 	:	val_out <= 4'hf211;
         4'h5331 	:	val_out <= 4'hf211;
         4'h5332 	:	val_out <= 4'hf211;
         4'h5333 	:	val_out <= 4'hf211;
         4'h5338 	:	val_out <= 4'hf205;
         4'h5339 	:	val_out <= 4'hf205;
         4'h533a 	:	val_out <= 4'hf205;
         4'h533b 	:	val_out <= 4'hf205;
         4'h5340 	:	val_out <= 4'hf1fa;
         4'h5341 	:	val_out <= 4'hf1fa;
         4'h5342 	:	val_out <= 4'hf1fa;
         4'h5343 	:	val_out <= 4'hf1fa;
         4'h5348 	:	val_out <= 4'hf1ee;
         4'h5349 	:	val_out <= 4'hf1ee;
         4'h534a 	:	val_out <= 4'hf1ee;
         4'h534b 	:	val_out <= 4'hf1ee;
         4'h5350 	:	val_out <= 4'hf1e3;
         4'h5351 	:	val_out <= 4'hf1e3;
         4'h5352 	:	val_out <= 4'hf1e3;
         4'h5353 	:	val_out <= 4'hf1e3;
         4'h5358 	:	val_out <= 4'hf1d7;
         4'h5359 	:	val_out <= 4'hf1d7;
         4'h535a 	:	val_out <= 4'hf1d7;
         4'h535b 	:	val_out <= 4'hf1d7;
         4'h5360 	:	val_out <= 4'hf1cc;
         4'h5361 	:	val_out <= 4'hf1cc;
         4'h5362 	:	val_out <= 4'hf1cc;
         4'h5363 	:	val_out <= 4'hf1cc;
         4'h5368 	:	val_out <= 4'hf1c0;
         4'h5369 	:	val_out <= 4'hf1c0;
         4'h536a 	:	val_out <= 4'hf1c0;
         4'h536b 	:	val_out <= 4'hf1c0;
         4'h5370 	:	val_out <= 4'hf1b5;
         4'h5371 	:	val_out <= 4'hf1b5;
         4'h5372 	:	val_out <= 4'hf1b5;
         4'h5373 	:	val_out <= 4'hf1b5;
         4'h5378 	:	val_out <= 4'hf1a9;
         4'h5379 	:	val_out <= 4'hf1a9;
         4'h537a 	:	val_out <= 4'hf1a9;
         4'h537b 	:	val_out <= 4'hf1a9;
         4'h5380 	:	val_out <= 4'hf19e;
         4'h5381 	:	val_out <= 4'hf19e;
         4'h5382 	:	val_out <= 4'hf19e;
         4'h5383 	:	val_out <= 4'hf19e;
         4'h5388 	:	val_out <= 4'hf192;
         4'h5389 	:	val_out <= 4'hf192;
         4'h538a 	:	val_out <= 4'hf192;
         4'h538b 	:	val_out <= 4'hf192;
         4'h5390 	:	val_out <= 4'hf186;
         4'h5391 	:	val_out <= 4'hf186;
         4'h5392 	:	val_out <= 4'hf186;
         4'h5393 	:	val_out <= 4'hf186;
         4'h5398 	:	val_out <= 4'hf17b;
         4'h5399 	:	val_out <= 4'hf17b;
         4'h539a 	:	val_out <= 4'hf17b;
         4'h539b 	:	val_out <= 4'hf17b;
         4'h53a0 	:	val_out <= 4'hf16f;
         4'h53a1 	:	val_out <= 4'hf16f;
         4'h53a2 	:	val_out <= 4'hf16f;
         4'h53a3 	:	val_out <= 4'hf16f;
         4'h53a8 	:	val_out <= 4'hf164;
         4'h53a9 	:	val_out <= 4'hf164;
         4'h53aa 	:	val_out <= 4'hf164;
         4'h53ab 	:	val_out <= 4'hf164;
         4'h53b0 	:	val_out <= 4'hf158;
         4'h53b1 	:	val_out <= 4'hf158;
         4'h53b2 	:	val_out <= 4'hf158;
         4'h53b3 	:	val_out <= 4'hf158;
         4'h53b8 	:	val_out <= 4'hf14c;
         4'h53b9 	:	val_out <= 4'hf14c;
         4'h53ba 	:	val_out <= 4'hf14c;
         4'h53bb 	:	val_out <= 4'hf14c;
         4'h53c0 	:	val_out <= 4'hf141;
         4'h53c1 	:	val_out <= 4'hf141;
         4'h53c2 	:	val_out <= 4'hf141;
         4'h53c3 	:	val_out <= 4'hf141;
         4'h53c8 	:	val_out <= 4'hf135;
         4'h53c9 	:	val_out <= 4'hf135;
         4'h53ca 	:	val_out <= 4'hf135;
         4'h53cb 	:	val_out <= 4'hf135;
         4'h53d0 	:	val_out <= 4'hf129;
         4'h53d1 	:	val_out <= 4'hf129;
         4'h53d2 	:	val_out <= 4'hf129;
         4'h53d3 	:	val_out <= 4'hf129;
         4'h53d8 	:	val_out <= 4'hf11d;
         4'h53d9 	:	val_out <= 4'hf11d;
         4'h53da 	:	val_out <= 4'hf11d;
         4'h53db 	:	val_out <= 4'hf11d;
         4'h53e0 	:	val_out <= 4'hf112;
         4'h53e1 	:	val_out <= 4'hf112;
         4'h53e2 	:	val_out <= 4'hf112;
         4'h53e3 	:	val_out <= 4'hf112;
         4'h53e8 	:	val_out <= 4'hf106;
         4'h53e9 	:	val_out <= 4'hf106;
         4'h53ea 	:	val_out <= 4'hf106;
         4'h53eb 	:	val_out <= 4'hf106;
         4'h53f0 	:	val_out <= 4'hf0fa;
         4'h53f1 	:	val_out <= 4'hf0fa;
         4'h53f2 	:	val_out <= 4'hf0fa;
         4'h53f3 	:	val_out <= 4'hf0fa;
         4'h53f8 	:	val_out <= 4'hf0ee;
         4'h53f9 	:	val_out <= 4'hf0ee;
         4'h53fa 	:	val_out <= 4'hf0ee;
         4'h53fb 	:	val_out <= 4'hf0ee;
         4'h5400 	:	val_out <= 4'hf0e2;
         4'h5401 	:	val_out <= 4'hf0e2;
         4'h5402 	:	val_out <= 4'hf0e2;
         4'h5403 	:	val_out <= 4'hf0e2;
         4'h5408 	:	val_out <= 4'hf0d6;
         4'h5409 	:	val_out <= 4'hf0d6;
         4'h540a 	:	val_out <= 4'hf0d6;
         4'h540b 	:	val_out <= 4'hf0d6;
         4'h5410 	:	val_out <= 4'hf0cb;
         4'h5411 	:	val_out <= 4'hf0cb;
         4'h5412 	:	val_out <= 4'hf0cb;
         4'h5413 	:	val_out <= 4'hf0cb;
         4'h5418 	:	val_out <= 4'hf0bf;
         4'h5419 	:	val_out <= 4'hf0bf;
         4'h541a 	:	val_out <= 4'hf0bf;
         4'h541b 	:	val_out <= 4'hf0bf;
         4'h5420 	:	val_out <= 4'hf0b3;
         4'h5421 	:	val_out <= 4'hf0b3;
         4'h5422 	:	val_out <= 4'hf0b3;
         4'h5423 	:	val_out <= 4'hf0b3;
         4'h5428 	:	val_out <= 4'hf0a7;
         4'h5429 	:	val_out <= 4'hf0a7;
         4'h542a 	:	val_out <= 4'hf0a7;
         4'h542b 	:	val_out <= 4'hf0a7;
         4'h5430 	:	val_out <= 4'hf09b;
         4'h5431 	:	val_out <= 4'hf09b;
         4'h5432 	:	val_out <= 4'hf09b;
         4'h5433 	:	val_out <= 4'hf09b;
         4'h5438 	:	val_out <= 4'hf08f;
         4'h5439 	:	val_out <= 4'hf08f;
         4'h543a 	:	val_out <= 4'hf08f;
         4'h543b 	:	val_out <= 4'hf08f;
         4'h5440 	:	val_out <= 4'hf083;
         4'h5441 	:	val_out <= 4'hf083;
         4'h5442 	:	val_out <= 4'hf083;
         4'h5443 	:	val_out <= 4'hf083;
         4'h5448 	:	val_out <= 4'hf077;
         4'h5449 	:	val_out <= 4'hf077;
         4'h544a 	:	val_out <= 4'hf077;
         4'h544b 	:	val_out <= 4'hf077;
         4'h5450 	:	val_out <= 4'hf06b;
         4'h5451 	:	val_out <= 4'hf06b;
         4'h5452 	:	val_out <= 4'hf06b;
         4'h5453 	:	val_out <= 4'hf06b;
         4'h5458 	:	val_out <= 4'hf05f;
         4'h5459 	:	val_out <= 4'hf05f;
         4'h545a 	:	val_out <= 4'hf05f;
         4'h545b 	:	val_out <= 4'hf05f;
         4'h5460 	:	val_out <= 4'hf053;
         4'h5461 	:	val_out <= 4'hf053;
         4'h5462 	:	val_out <= 4'hf053;
         4'h5463 	:	val_out <= 4'hf053;
         4'h5468 	:	val_out <= 4'hf047;
         4'h5469 	:	val_out <= 4'hf047;
         4'h546a 	:	val_out <= 4'hf047;
         4'h546b 	:	val_out <= 4'hf047;
         4'h5470 	:	val_out <= 4'hf03b;
         4'h5471 	:	val_out <= 4'hf03b;
         4'h5472 	:	val_out <= 4'hf03b;
         4'h5473 	:	val_out <= 4'hf03b;
         4'h5478 	:	val_out <= 4'hf02f;
         4'h5479 	:	val_out <= 4'hf02f;
         4'h547a 	:	val_out <= 4'hf02f;
         4'h547b 	:	val_out <= 4'hf02f;
         4'h5480 	:	val_out <= 4'hf023;
         4'h5481 	:	val_out <= 4'hf023;
         4'h5482 	:	val_out <= 4'hf023;
         4'h5483 	:	val_out <= 4'hf023;
         4'h5488 	:	val_out <= 4'hf016;
         4'h5489 	:	val_out <= 4'hf016;
         4'h548a 	:	val_out <= 4'hf016;
         4'h548b 	:	val_out <= 4'hf016;
         4'h5490 	:	val_out <= 4'hf00a;
         4'h5491 	:	val_out <= 4'hf00a;
         4'h5492 	:	val_out <= 4'hf00a;
         4'h5493 	:	val_out <= 4'hf00a;
         4'h5498 	:	val_out <= 4'heffe;
         4'h5499 	:	val_out <= 4'heffe;
         4'h549a 	:	val_out <= 4'heffe;
         4'h549b 	:	val_out <= 4'heffe;
         4'h54a0 	:	val_out <= 4'heff2;
         4'h54a1 	:	val_out <= 4'heff2;
         4'h54a2 	:	val_out <= 4'heff2;
         4'h54a3 	:	val_out <= 4'heff2;
         4'h54a8 	:	val_out <= 4'hefe6;
         4'h54a9 	:	val_out <= 4'hefe6;
         4'h54aa 	:	val_out <= 4'hefe6;
         4'h54ab 	:	val_out <= 4'hefe6;
         4'h54b0 	:	val_out <= 4'hefda;
         4'h54b1 	:	val_out <= 4'hefda;
         4'h54b2 	:	val_out <= 4'hefda;
         4'h54b3 	:	val_out <= 4'hefda;
         4'h54b8 	:	val_out <= 4'hefcd;
         4'h54b9 	:	val_out <= 4'hefcd;
         4'h54ba 	:	val_out <= 4'hefcd;
         4'h54bb 	:	val_out <= 4'hefcd;
         4'h54c0 	:	val_out <= 4'hefc1;
         4'h54c1 	:	val_out <= 4'hefc1;
         4'h54c2 	:	val_out <= 4'hefc1;
         4'h54c3 	:	val_out <= 4'hefc1;
         4'h54c8 	:	val_out <= 4'hefb5;
         4'h54c9 	:	val_out <= 4'hefb5;
         4'h54ca 	:	val_out <= 4'hefb5;
         4'h54cb 	:	val_out <= 4'hefb5;
         4'h54d0 	:	val_out <= 4'hefa9;
         4'h54d1 	:	val_out <= 4'hefa9;
         4'h54d2 	:	val_out <= 4'hefa9;
         4'h54d3 	:	val_out <= 4'hefa9;
         4'h54d8 	:	val_out <= 4'hef9c;
         4'h54d9 	:	val_out <= 4'hef9c;
         4'h54da 	:	val_out <= 4'hef9c;
         4'h54db 	:	val_out <= 4'hef9c;
         4'h54e0 	:	val_out <= 4'hef90;
         4'h54e1 	:	val_out <= 4'hef90;
         4'h54e2 	:	val_out <= 4'hef90;
         4'h54e3 	:	val_out <= 4'hef90;
         4'h54e8 	:	val_out <= 4'hef84;
         4'h54e9 	:	val_out <= 4'hef84;
         4'h54ea 	:	val_out <= 4'hef84;
         4'h54eb 	:	val_out <= 4'hef84;
         4'h54f0 	:	val_out <= 4'hef77;
         4'h54f1 	:	val_out <= 4'hef77;
         4'h54f2 	:	val_out <= 4'hef77;
         4'h54f3 	:	val_out <= 4'hef77;
         4'h54f8 	:	val_out <= 4'hef6b;
         4'h54f9 	:	val_out <= 4'hef6b;
         4'h54fa 	:	val_out <= 4'hef6b;
         4'h54fb 	:	val_out <= 4'hef6b;
         4'h5500 	:	val_out <= 4'hef5f;
         4'h5501 	:	val_out <= 4'hef5f;
         4'h5502 	:	val_out <= 4'hef5f;
         4'h5503 	:	val_out <= 4'hef5f;
         4'h5508 	:	val_out <= 4'hef52;
         4'h5509 	:	val_out <= 4'hef52;
         4'h550a 	:	val_out <= 4'hef52;
         4'h550b 	:	val_out <= 4'hef52;
         4'h5510 	:	val_out <= 4'hef46;
         4'h5511 	:	val_out <= 4'hef46;
         4'h5512 	:	val_out <= 4'hef46;
         4'h5513 	:	val_out <= 4'hef46;
         4'h5518 	:	val_out <= 4'hef39;
         4'h5519 	:	val_out <= 4'hef39;
         4'h551a 	:	val_out <= 4'hef39;
         4'h551b 	:	val_out <= 4'hef39;
         4'h5520 	:	val_out <= 4'hef2d;
         4'h5521 	:	val_out <= 4'hef2d;
         4'h5522 	:	val_out <= 4'hef2d;
         4'h5523 	:	val_out <= 4'hef2d;
         4'h5528 	:	val_out <= 4'hef20;
         4'h5529 	:	val_out <= 4'hef20;
         4'h552a 	:	val_out <= 4'hef20;
         4'h552b 	:	val_out <= 4'hef20;
         4'h5530 	:	val_out <= 4'hef14;
         4'h5531 	:	val_out <= 4'hef14;
         4'h5532 	:	val_out <= 4'hef14;
         4'h5533 	:	val_out <= 4'hef14;
         4'h5538 	:	val_out <= 4'hef07;
         4'h5539 	:	val_out <= 4'hef07;
         4'h553a 	:	val_out <= 4'hef07;
         4'h553b 	:	val_out <= 4'hef07;
         4'h5540 	:	val_out <= 4'heefb;
         4'h5541 	:	val_out <= 4'heefb;
         4'h5542 	:	val_out <= 4'heefb;
         4'h5543 	:	val_out <= 4'heefb;
         4'h5548 	:	val_out <= 4'heeee;
         4'h5549 	:	val_out <= 4'heeee;
         4'h554a 	:	val_out <= 4'heeee;
         4'h554b 	:	val_out <= 4'heeee;
         4'h5550 	:	val_out <= 4'heee2;
         4'h5551 	:	val_out <= 4'heee2;
         4'h5552 	:	val_out <= 4'heee2;
         4'h5553 	:	val_out <= 4'heee2;
         4'h5558 	:	val_out <= 4'heed5;
         4'h5559 	:	val_out <= 4'heed5;
         4'h555a 	:	val_out <= 4'heed5;
         4'h555b 	:	val_out <= 4'heed5;
         4'h5560 	:	val_out <= 4'heec9;
         4'h5561 	:	val_out <= 4'heec9;
         4'h5562 	:	val_out <= 4'heec9;
         4'h5563 	:	val_out <= 4'heec9;
         4'h5568 	:	val_out <= 4'heebc;
         4'h5569 	:	val_out <= 4'heebc;
         4'h556a 	:	val_out <= 4'heebc;
         4'h556b 	:	val_out <= 4'heebc;
         4'h5570 	:	val_out <= 4'heeaf;
         4'h5571 	:	val_out <= 4'heeaf;
         4'h5572 	:	val_out <= 4'heeaf;
         4'h5573 	:	val_out <= 4'heeaf;
         4'h5578 	:	val_out <= 4'heea3;
         4'h5579 	:	val_out <= 4'heea3;
         4'h557a 	:	val_out <= 4'heea3;
         4'h557b 	:	val_out <= 4'heea3;
         4'h5580 	:	val_out <= 4'hee96;
         4'h5581 	:	val_out <= 4'hee96;
         4'h5582 	:	val_out <= 4'hee96;
         4'h5583 	:	val_out <= 4'hee96;
         4'h5588 	:	val_out <= 4'hee89;
         4'h5589 	:	val_out <= 4'hee89;
         4'h558a 	:	val_out <= 4'hee89;
         4'h558b 	:	val_out <= 4'hee89;
         4'h5590 	:	val_out <= 4'hee7d;
         4'h5591 	:	val_out <= 4'hee7d;
         4'h5592 	:	val_out <= 4'hee7d;
         4'h5593 	:	val_out <= 4'hee7d;
         4'h5598 	:	val_out <= 4'hee70;
         4'h5599 	:	val_out <= 4'hee70;
         4'h559a 	:	val_out <= 4'hee70;
         4'h559b 	:	val_out <= 4'hee70;
         4'h55a0 	:	val_out <= 4'hee63;
         4'h55a1 	:	val_out <= 4'hee63;
         4'h55a2 	:	val_out <= 4'hee63;
         4'h55a3 	:	val_out <= 4'hee63;
         4'h55a8 	:	val_out <= 4'hee57;
         4'h55a9 	:	val_out <= 4'hee57;
         4'h55aa 	:	val_out <= 4'hee57;
         4'h55ab 	:	val_out <= 4'hee57;
         4'h55b0 	:	val_out <= 4'hee4a;
         4'h55b1 	:	val_out <= 4'hee4a;
         4'h55b2 	:	val_out <= 4'hee4a;
         4'h55b3 	:	val_out <= 4'hee4a;
         4'h55b8 	:	val_out <= 4'hee3d;
         4'h55b9 	:	val_out <= 4'hee3d;
         4'h55ba 	:	val_out <= 4'hee3d;
         4'h55bb 	:	val_out <= 4'hee3d;
         4'h55c0 	:	val_out <= 4'hee30;
         4'h55c1 	:	val_out <= 4'hee30;
         4'h55c2 	:	val_out <= 4'hee30;
         4'h55c3 	:	val_out <= 4'hee30;
         4'h55c8 	:	val_out <= 4'hee24;
         4'h55c9 	:	val_out <= 4'hee24;
         4'h55ca 	:	val_out <= 4'hee24;
         4'h55cb 	:	val_out <= 4'hee24;
         4'h55d0 	:	val_out <= 4'hee17;
         4'h55d1 	:	val_out <= 4'hee17;
         4'h55d2 	:	val_out <= 4'hee17;
         4'h55d3 	:	val_out <= 4'hee17;
         4'h55d8 	:	val_out <= 4'hee0a;
         4'h55d9 	:	val_out <= 4'hee0a;
         4'h55da 	:	val_out <= 4'hee0a;
         4'h55db 	:	val_out <= 4'hee0a;
         4'h55e0 	:	val_out <= 4'hedfd;
         4'h55e1 	:	val_out <= 4'hedfd;
         4'h55e2 	:	val_out <= 4'hedfd;
         4'h55e3 	:	val_out <= 4'hedfd;
         4'h55e8 	:	val_out <= 4'hedf0;
         4'h55e9 	:	val_out <= 4'hedf0;
         4'h55ea 	:	val_out <= 4'hedf0;
         4'h55eb 	:	val_out <= 4'hedf0;
         4'h55f0 	:	val_out <= 4'hede3;
         4'h55f1 	:	val_out <= 4'hede3;
         4'h55f2 	:	val_out <= 4'hede3;
         4'h55f3 	:	val_out <= 4'hede3;
         4'h55f8 	:	val_out <= 4'hedd6;
         4'h55f9 	:	val_out <= 4'hedd6;
         4'h55fa 	:	val_out <= 4'hedd6;
         4'h55fb 	:	val_out <= 4'hedd6;
         4'h5600 	:	val_out <= 4'hedca;
         4'h5601 	:	val_out <= 4'hedca;
         4'h5602 	:	val_out <= 4'hedca;
         4'h5603 	:	val_out <= 4'hedca;
         4'h5608 	:	val_out <= 4'hedbd;
         4'h5609 	:	val_out <= 4'hedbd;
         4'h560a 	:	val_out <= 4'hedbd;
         4'h560b 	:	val_out <= 4'hedbd;
         4'h5610 	:	val_out <= 4'hedb0;
         4'h5611 	:	val_out <= 4'hedb0;
         4'h5612 	:	val_out <= 4'hedb0;
         4'h5613 	:	val_out <= 4'hedb0;
         4'h5618 	:	val_out <= 4'heda3;
         4'h5619 	:	val_out <= 4'heda3;
         4'h561a 	:	val_out <= 4'heda3;
         4'h561b 	:	val_out <= 4'heda3;
         4'h5620 	:	val_out <= 4'hed96;
         4'h5621 	:	val_out <= 4'hed96;
         4'h5622 	:	val_out <= 4'hed96;
         4'h5623 	:	val_out <= 4'hed96;
         4'h5628 	:	val_out <= 4'hed89;
         4'h5629 	:	val_out <= 4'hed89;
         4'h562a 	:	val_out <= 4'hed89;
         4'h562b 	:	val_out <= 4'hed89;
         4'h5630 	:	val_out <= 4'hed7c;
         4'h5631 	:	val_out <= 4'hed7c;
         4'h5632 	:	val_out <= 4'hed7c;
         4'h5633 	:	val_out <= 4'hed7c;
         4'h5638 	:	val_out <= 4'hed6f;
         4'h5639 	:	val_out <= 4'hed6f;
         4'h563a 	:	val_out <= 4'hed6f;
         4'h563b 	:	val_out <= 4'hed6f;
         4'h5640 	:	val_out <= 4'hed62;
         4'h5641 	:	val_out <= 4'hed62;
         4'h5642 	:	val_out <= 4'hed62;
         4'h5643 	:	val_out <= 4'hed62;
         4'h5648 	:	val_out <= 4'hed55;
         4'h5649 	:	val_out <= 4'hed55;
         4'h564a 	:	val_out <= 4'hed55;
         4'h564b 	:	val_out <= 4'hed55;
         4'h5650 	:	val_out <= 4'hed48;
         4'h5651 	:	val_out <= 4'hed48;
         4'h5652 	:	val_out <= 4'hed48;
         4'h5653 	:	val_out <= 4'hed48;
         4'h5658 	:	val_out <= 4'hed3a;
         4'h5659 	:	val_out <= 4'hed3a;
         4'h565a 	:	val_out <= 4'hed3a;
         4'h565b 	:	val_out <= 4'hed3a;
         4'h5660 	:	val_out <= 4'hed2d;
         4'h5661 	:	val_out <= 4'hed2d;
         4'h5662 	:	val_out <= 4'hed2d;
         4'h5663 	:	val_out <= 4'hed2d;
         4'h5668 	:	val_out <= 4'hed20;
         4'h5669 	:	val_out <= 4'hed20;
         4'h566a 	:	val_out <= 4'hed20;
         4'h566b 	:	val_out <= 4'hed20;
         4'h5670 	:	val_out <= 4'hed13;
         4'h5671 	:	val_out <= 4'hed13;
         4'h5672 	:	val_out <= 4'hed13;
         4'h5673 	:	val_out <= 4'hed13;
         4'h5678 	:	val_out <= 4'hed06;
         4'h5679 	:	val_out <= 4'hed06;
         4'h567a 	:	val_out <= 4'hed06;
         4'h567b 	:	val_out <= 4'hed06;
         4'h5680 	:	val_out <= 4'hecf9;
         4'h5681 	:	val_out <= 4'hecf9;
         4'h5682 	:	val_out <= 4'hecf9;
         4'h5683 	:	val_out <= 4'hecf9;
         4'h5688 	:	val_out <= 4'hecec;
         4'h5689 	:	val_out <= 4'hecec;
         4'h568a 	:	val_out <= 4'hecec;
         4'h568b 	:	val_out <= 4'hecec;
         4'h5690 	:	val_out <= 4'hecde;
         4'h5691 	:	val_out <= 4'hecde;
         4'h5692 	:	val_out <= 4'hecde;
         4'h5693 	:	val_out <= 4'hecde;
         4'h5698 	:	val_out <= 4'hecd1;
         4'h5699 	:	val_out <= 4'hecd1;
         4'h569a 	:	val_out <= 4'hecd1;
         4'h569b 	:	val_out <= 4'hecd1;
         4'h56a0 	:	val_out <= 4'hecc4;
         4'h56a1 	:	val_out <= 4'hecc4;
         4'h56a2 	:	val_out <= 4'hecc4;
         4'h56a3 	:	val_out <= 4'hecc4;
         4'h56a8 	:	val_out <= 4'hecb7;
         4'h56a9 	:	val_out <= 4'hecb7;
         4'h56aa 	:	val_out <= 4'hecb7;
         4'h56ab 	:	val_out <= 4'hecb7;
         4'h56b0 	:	val_out <= 4'heca9;
         4'h56b1 	:	val_out <= 4'heca9;
         4'h56b2 	:	val_out <= 4'heca9;
         4'h56b3 	:	val_out <= 4'heca9;
         4'h56b8 	:	val_out <= 4'hec9c;
         4'h56b9 	:	val_out <= 4'hec9c;
         4'h56ba 	:	val_out <= 4'hec9c;
         4'h56bb 	:	val_out <= 4'hec9c;
         4'h56c0 	:	val_out <= 4'hec8f;
         4'h56c1 	:	val_out <= 4'hec8f;
         4'h56c2 	:	val_out <= 4'hec8f;
         4'h56c3 	:	val_out <= 4'hec8f;
         4'h56c8 	:	val_out <= 4'hec81;
         4'h56c9 	:	val_out <= 4'hec81;
         4'h56ca 	:	val_out <= 4'hec81;
         4'h56cb 	:	val_out <= 4'hec81;
         4'h56d0 	:	val_out <= 4'hec74;
         4'h56d1 	:	val_out <= 4'hec74;
         4'h56d2 	:	val_out <= 4'hec74;
         4'h56d3 	:	val_out <= 4'hec74;
         4'h56d8 	:	val_out <= 4'hec67;
         4'h56d9 	:	val_out <= 4'hec67;
         4'h56da 	:	val_out <= 4'hec67;
         4'h56db 	:	val_out <= 4'hec67;
         4'h56e0 	:	val_out <= 4'hec59;
         4'h56e1 	:	val_out <= 4'hec59;
         4'h56e2 	:	val_out <= 4'hec59;
         4'h56e3 	:	val_out <= 4'hec59;
         4'h56e8 	:	val_out <= 4'hec4c;
         4'h56e9 	:	val_out <= 4'hec4c;
         4'h56ea 	:	val_out <= 4'hec4c;
         4'h56eb 	:	val_out <= 4'hec4c;
         4'h56f0 	:	val_out <= 4'hec3f;
         4'h56f1 	:	val_out <= 4'hec3f;
         4'h56f2 	:	val_out <= 4'hec3f;
         4'h56f3 	:	val_out <= 4'hec3f;
         4'h56f8 	:	val_out <= 4'hec31;
         4'h56f9 	:	val_out <= 4'hec31;
         4'h56fa 	:	val_out <= 4'hec31;
         4'h56fb 	:	val_out <= 4'hec31;
         4'h5700 	:	val_out <= 4'hec24;
         4'h5701 	:	val_out <= 4'hec24;
         4'h5702 	:	val_out <= 4'hec24;
         4'h5703 	:	val_out <= 4'hec24;
         4'h5708 	:	val_out <= 4'hec16;
         4'h5709 	:	val_out <= 4'hec16;
         4'h570a 	:	val_out <= 4'hec16;
         4'h570b 	:	val_out <= 4'hec16;
         4'h5710 	:	val_out <= 4'hec09;
         4'h5711 	:	val_out <= 4'hec09;
         4'h5712 	:	val_out <= 4'hec09;
         4'h5713 	:	val_out <= 4'hec09;
         4'h5718 	:	val_out <= 4'hebfb;
         4'h5719 	:	val_out <= 4'hebfb;
         4'h571a 	:	val_out <= 4'hebfb;
         4'h571b 	:	val_out <= 4'hebfb;
         4'h5720 	:	val_out <= 4'hebee;
         4'h5721 	:	val_out <= 4'hebee;
         4'h5722 	:	val_out <= 4'hebee;
         4'h5723 	:	val_out <= 4'hebee;
         4'h5728 	:	val_out <= 4'hebe0;
         4'h5729 	:	val_out <= 4'hebe0;
         4'h572a 	:	val_out <= 4'hebe0;
         4'h572b 	:	val_out <= 4'hebe0;
         4'h5730 	:	val_out <= 4'hebd3;
         4'h5731 	:	val_out <= 4'hebd3;
         4'h5732 	:	val_out <= 4'hebd3;
         4'h5733 	:	val_out <= 4'hebd3;
         4'h5738 	:	val_out <= 4'hebc5;
         4'h5739 	:	val_out <= 4'hebc5;
         4'h573a 	:	val_out <= 4'hebc5;
         4'h573b 	:	val_out <= 4'hebc5;
         4'h5740 	:	val_out <= 4'hebb8;
         4'h5741 	:	val_out <= 4'hebb8;
         4'h5742 	:	val_out <= 4'hebb8;
         4'h5743 	:	val_out <= 4'hebb8;
         4'h5748 	:	val_out <= 4'hebaa;
         4'h5749 	:	val_out <= 4'hebaa;
         4'h574a 	:	val_out <= 4'hebaa;
         4'h574b 	:	val_out <= 4'hebaa;
         4'h5750 	:	val_out <= 4'heb9c;
         4'h5751 	:	val_out <= 4'heb9c;
         4'h5752 	:	val_out <= 4'heb9c;
         4'h5753 	:	val_out <= 4'heb9c;
         4'h5758 	:	val_out <= 4'heb8f;
         4'h5759 	:	val_out <= 4'heb8f;
         4'h575a 	:	val_out <= 4'heb8f;
         4'h575b 	:	val_out <= 4'heb8f;
         4'h5760 	:	val_out <= 4'heb81;
         4'h5761 	:	val_out <= 4'heb81;
         4'h5762 	:	val_out <= 4'heb81;
         4'h5763 	:	val_out <= 4'heb81;
         4'h5768 	:	val_out <= 4'heb73;
         4'h5769 	:	val_out <= 4'heb73;
         4'h576a 	:	val_out <= 4'heb73;
         4'h576b 	:	val_out <= 4'heb73;
         4'h5770 	:	val_out <= 4'heb66;
         4'h5771 	:	val_out <= 4'heb66;
         4'h5772 	:	val_out <= 4'heb66;
         4'h5773 	:	val_out <= 4'heb66;
         4'h5778 	:	val_out <= 4'heb58;
         4'h5779 	:	val_out <= 4'heb58;
         4'h577a 	:	val_out <= 4'heb58;
         4'h577b 	:	val_out <= 4'heb58;
         4'h5780 	:	val_out <= 4'heb4a;
         4'h5781 	:	val_out <= 4'heb4a;
         4'h5782 	:	val_out <= 4'heb4a;
         4'h5783 	:	val_out <= 4'heb4a;
         4'h5788 	:	val_out <= 4'heb3d;
         4'h5789 	:	val_out <= 4'heb3d;
         4'h578a 	:	val_out <= 4'heb3d;
         4'h578b 	:	val_out <= 4'heb3d;
         4'h5790 	:	val_out <= 4'heb2f;
         4'h5791 	:	val_out <= 4'heb2f;
         4'h5792 	:	val_out <= 4'heb2f;
         4'h5793 	:	val_out <= 4'heb2f;
         4'h5798 	:	val_out <= 4'heb21;
         4'h5799 	:	val_out <= 4'heb21;
         4'h579a 	:	val_out <= 4'heb21;
         4'h579b 	:	val_out <= 4'heb21;
         4'h57a0 	:	val_out <= 4'heb13;
         4'h57a1 	:	val_out <= 4'heb13;
         4'h57a2 	:	val_out <= 4'heb13;
         4'h57a3 	:	val_out <= 4'heb13;
         4'h57a8 	:	val_out <= 4'heb06;
         4'h57a9 	:	val_out <= 4'heb06;
         4'h57aa 	:	val_out <= 4'heb06;
         4'h57ab 	:	val_out <= 4'heb06;
         4'h57b0 	:	val_out <= 4'heaf8;
         4'h57b1 	:	val_out <= 4'heaf8;
         4'h57b2 	:	val_out <= 4'heaf8;
         4'h57b3 	:	val_out <= 4'heaf8;
         4'h57b8 	:	val_out <= 4'heaea;
         4'h57b9 	:	val_out <= 4'heaea;
         4'h57ba 	:	val_out <= 4'heaea;
         4'h57bb 	:	val_out <= 4'heaea;
         4'h57c0 	:	val_out <= 4'headc;
         4'h57c1 	:	val_out <= 4'headc;
         4'h57c2 	:	val_out <= 4'headc;
         4'h57c3 	:	val_out <= 4'headc;
         4'h57c8 	:	val_out <= 4'heace;
         4'h57c9 	:	val_out <= 4'heace;
         4'h57ca 	:	val_out <= 4'heace;
         4'h57cb 	:	val_out <= 4'heace;
         4'h57d0 	:	val_out <= 4'heac1;
         4'h57d1 	:	val_out <= 4'heac1;
         4'h57d2 	:	val_out <= 4'heac1;
         4'h57d3 	:	val_out <= 4'heac1;
         4'h57d8 	:	val_out <= 4'heab3;
         4'h57d9 	:	val_out <= 4'heab3;
         4'h57da 	:	val_out <= 4'heab3;
         4'h57db 	:	val_out <= 4'heab3;
         4'h57e0 	:	val_out <= 4'heaa5;
         4'h57e1 	:	val_out <= 4'heaa5;
         4'h57e2 	:	val_out <= 4'heaa5;
         4'h57e3 	:	val_out <= 4'heaa5;
         4'h57e8 	:	val_out <= 4'hea97;
         4'h57e9 	:	val_out <= 4'hea97;
         4'h57ea 	:	val_out <= 4'hea97;
         4'h57eb 	:	val_out <= 4'hea97;
         4'h57f0 	:	val_out <= 4'hea89;
         4'h57f1 	:	val_out <= 4'hea89;
         4'h57f2 	:	val_out <= 4'hea89;
         4'h57f3 	:	val_out <= 4'hea89;
         4'h57f8 	:	val_out <= 4'hea7b;
         4'h57f9 	:	val_out <= 4'hea7b;
         4'h57fa 	:	val_out <= 4'hea7b;
         4'h57fb 	:	val_out <= 4'hea7b;
         4'h5800 	:	val_out <= 4'hea6d;
         4'h5801 	:	val_out <= 4'hea6d;
         4'h5802 	:	val_out <= 4'hea6d;
         4'h5803 	:	val_out <= 4'hea6d;
         4'h5808 	:	val_out <= 4'hea5f;
         4'h5809 	:	val_out <= 4'hea5f;
         4'h580a 	:	val_out <= 4'hea5f;
         4'h580b 	:	val_out <= 4'hea5f;
         4'h5810 	:	val_out <= 4'hea51;
         4'h5811 	:	val_out <= 4'hea51;
         4'h5812 	:	val_out <= 4'hea51;
         4'h5813 	:	val_out <= 4'hea51;
         4'h5818 	:	val_out <= 4'hea43;
         4'h5819 	:	val_out <= 4'hea43;
         4'h581a 	:	val_out <= 4'hea43;
         4'h581b 	:	val_out <= 4'hea43;
         4'h5820 	:	val_out <= 4'hea35;
         4'h5821 	:	val_out <= 4'hea35;
         4'h5822 	:	val_out <= 4'hea35;
         4'h5823 	:	val_out <= 4'hea35;
         4'h5828 	:	val_out <= 4'hea27;
         4'h5829 	:	val_out <= 4'hea27;
         4'h582a 	:	val_out <= 4'hea27;
         4'h582b 	:	val_out <= 4'hea27;
         4'h5830 	:	val_out <= 4'hea19;
         4'h5831 	:	val_out <= 4'hea19;
         4'h5832 	:	val_out <= 4'hea19;
         4'h5833 	:	val_out <= 4'hea19;
         4'h5838 	:	val_out <= 4'hea0b;
         4'h5839 	:	val_out <= 4'hea0b;
         4'h583a 	:	val_out <= 4'hea0b;
         4'h583b 	:	val_out <= 4'hea0b;
         4'h5840 	:	val_out <= 4'he9fd;
         4'h5841 	:	val_out <= 4'he9fd;
         4'h5842 	:	val_out <= 4'he9fd;
         4'h5843 	:	val_out <= 4'he9fd;
         4'h5848 	:	val_out <= 4'he9ef;
         4'h5849 	:	val_out <= 4'he9ef;
         4'h584a 	:	val_out <= 4'he9ef;
         4'h584b 	:	val_out <= 4'he9ef;
         4'h5850 	:	val_out <= 4'he9e1;
         4'h5851 	:	val_out <= 4'he9e1;
         4'h5852 	:	val_out <= 4'he9e1;
         4'h5853 	:	val_out <= 4'he9e1;
         4'h5858 	:	val_out <= 4'he9d3;
         4'h5859 	:	val_out <= 4'he9d3;
         4'h585a 	:	val_out <= 4'he9d3;
         4'h585b 	:	val_out <= 4'he9d3;
         4'h5860 	:	val_out <= 4'he9c4;
         4'h5861 	:	val_out <= 4'he9c4;
         4'h5862 	:	val_out <= 4'he9c4;
         4'h5863 	:	val_out <= 4'he9c4;
         4'h5868 	:	val_out <= 4'he9b6;
         4'h5869 	:	val_out <= 4'he9b6;
         4'h586a 	:	val_out <= 4'he9b6;
         4'h586b 	:	val_out <= 4'he9b6;
         4'h5870 	:	val_out <= 4'he9a8;
         4'h5871 	:	val_out <= 4'he9a8;
         4'h5872 	:	val_out <= 4'he9a8;
         4'h5873 	:	val_out <= 4'he9a8;
         4'h5878 	:	val_out <= 4'he99a;
         4'h5879 	:	val_out <= 4'he99a;
         4'h587a 	:	val_out <= 4'he99a;
         4'h587b 	:	val_out <= 4'he99a;
         4'h5880 	:	val_out <= 4'he98c;
         4'h5881 	:	val_out <= 4'he98c;
         4'h5882 	:	val_out <= 4'he98c;
         4'h5883 	:	val_out <= 4'he98c;
         4'h5888 	:	val_out <= 4'he97d;
         4'h5889 	:	val_out <= 4'he97d;
         4'h588a 	:	val_out <= 4'he97d;
         4'h588b 	:	val_out <= 4'he97d;
         4'h5890 	:	val_out <= 4'he96f;
         4'h5891 	:	val_out <= 4'he96f;
         4'h5892 	:	val_out <= 4'he96f;
         4'h5893 	:	val_out <= 4'he96f;
         4'h5898 	:	val_out <= 4'he961;
         4'h5899 	:	val_out <= 4'he961;
         4'h589a 	:	val_out <= 4'he961;
         4'h589b 	:	val_out <= 4'he961;
         4'h58a0 	:	val_out <= 4'he953;
         4'h58a1 	:	val_out <= 4'he953;
         4'h58a2 	:	val_out <= 4'he953;
         4'h58a3 	:	val_out <= 4'he953;
         4'h58a8 	:	val_out <= 4'he944;
         4'h58a9 	:	val_out <= 4'he944;
         4'h58aa 	:	val_out <= 4'he944;
         4'h58ab 	:	val_out <= 4'he944;
         4'h58b0 	:	val_out <= 4'he936;
         4'h58b1 	:	val_out <= 4'he936;
         4'h58b2 	:	val_out <= 4'he936;
         4'h58b3 	:	val_out <= 4'he936;
         4'h58b8 	:	val_out <= 4'he928;
         4'h58b9 	:	val_out <= 4'he928;
         4'h58ba 	:	val_out <= 4'he928;
         4'h58bb 	:	val_out <= 4'he928;
         4'h58c0 	:	val_out <= 4'he919;
         4'h58c1 	:	val_out <= 4'he919;
         4'h58c2 	:	val_out <= 4'he919;
         4'h58c3 	:	val_out <= 4'he919;
         4'h58c8 	:	val_out <= 4'he90b;
         4'h58c9 	:	val_out <= 4'he90b;
         4'h58ca 	:	val_out <= 4'he90b;
         4'h58cb 	:	val_out <= 4'he90b;
         4'h58d0 	:	val_out <= 4'he8fd;
         4'h58d1 	:	val_out <= 4'he8fd;
         4'h58d2 	:	val_out <= 4'he8fd;
         4'h58d3 	:	val_out <= 4'he8fd;
         4'h58d8 	:	val_out <= 4'he8ee;
         4'h58d9 	:	val_out <= 4'he8ee;
         4'h58da 	:	val_out <= 4'he8ee;
         4'h58db 	:	val_out <= 4'he8ee;
         4'h58e0 	:	val_out <= 4'he8e0;
         4'h58e1 	:	val_out <= 4'he8e0;
         4'h58e2 	:	val_out <= 4'he8e0;
         4'h58e3 	:	val_out <= 4'he8e0;
         4'h58e8 	:	val_out <= 4'he8d1;
         4'h58e9 	:	val_out <= 4'he8d1;
         4'h58ea 	:	val_out <= 4'he8d1;
         4'h58eb 	:	val_out <= 4'he8d1;
         4'h58f0 	:	val_out <= 4'he8c3;
         4'h58f1 	:	val_out <= 4'he8c3;
         4'h58f2 	:	val_out <= 4'he8c3;
         4'h58f3 	:	val_out <= 4'he8c3;
         4'h58f8 	:	val_out <= 4'he8b5;
         4'h58f9 	:	val_out <= 4'he8b5;
         4'h58fa 	:	val_out <= 4'he8b5;
         4'h58fb 	:	val_out <= 4'he8b5;
         4'h5900 	:	val_out <= 4'he8a6;
         4'h5901 	:	val_out <= 4'he8a6;
         4'h5902 	:	val_out <= 4'he8a6;
         4'h5903 	:	val_out <= 4'he8a6;
         4'h5908 	:	val_out <= 4'he898;
         4'h5909 	:	val_out <= 4'he898;
         4'h590a 	:	val_out <= 4'he898;
         4'h590b 	:	val_out <= 4'he898;
         4'h5910 	:	val_out <= 4'he889;
         4'h5911 	:	val_out <= 4'he889;
         4'h5912 	:	val_out <= 4'he889;
         4'h5913 	:	val_out <= 4'he889;
         4'h5918 	:	val_out <= 4'he87b;
         4'h5919 	:	val_out <= 4'he87b;
         4'h591a 	:	val_out <= 4'he87b;
         4'h591b 	:	val_out <= 4'he87b;
         4'h5920 	:	val_out <= 4'he86c;
         4'h5921 	:	val_out <= 4'he86c;
         4'h5922 	:	val_out <= 4'he86c;
         4'h5923 	:	val_out <= 4'he86c;
         4'h5928 	:	val_out <= 4'he85e;
         4'h5929 	:	val_out <= 4'he85e;
         4'h592a 	:	val_out <= 4'he85e;
         4'h592b 	:	val_out <= 4'he85e;
         4'h5930 	:	val_out <= 4'he84f;
         4'h5931 	:	val_out <= 4'he84f;
         4'h5932 	:	val_out <= 4'he84f;
         4'h5933 	:	val_out <= 4'he84f;
         4'h5938 	:	val_out <= 4'he840;
         4'h5939 	:	val_out <= 4'he840;
         4'h593a 	:	val_out <= 4'he840;
         4'h593b 	:	val_out <= 4'he840;
         4'h5940 	:	val_out <= 4'he832;
         4'h5941 	:	val_out <= 4'he832;
         4'h5942 	:	val_out <= 4'he832;
         4'h5943 	:	val_out <= 4'he832;
         4'h5948 	:	val_out <= 4'he823;
         4'h5949 	:	val_out <= 4'he823;
         4'h594a 	:	val_out <= 4'he823;
         4'h594b 	:	val_out <= 4'he823;
         4'h5950 	:	val_out <= 4'he815;
         4'h5951 	:	val_out <= 4'he815;
         4'h5952 	:	val_out <= 4'he815;
         4'h5953 	:	val_out <= 4'he815;
         4'h5958 	:	val_out <= 4'he806;
         4'h5959 	:	val_out <= 4'he806;
         4'h595a 	:	val_out <= 4'he806;
         4'h595b 	:	val_out <= 4'he806;
         4'h5960 	:	val_out <= 4'he7f7;
         4'h5961 	:	val_out <= 4'he7f7;
         4'h5962 	:	val_out <= 4'he7f7;
         4'h5963 	:	val_out <= 4'he7f7;
         4'h5968 	:	val_out <= 4'he7e9;
         4'h5969 	:	val_out <= 4'he7e9;
         4'h596a 	:	val_out <= 4'he7e9;
         4'h596b 	:	val_out <= 4'he7e9;
         4'h5970 	:	val_out <= 4'he7da;
         4'h5971 	:	val_out <= 4'he7da;
         4'h5972 	:	val_out <= 4'he7da;
         4'h5973 	:	val_out <= 4'he7da;
         4'h5978 	:	val_out <= 4'he7cb;
         4'h5979 	:	val_out <= 4'he7cb;
         4'h597a 	:	val_out <= 4'he7cb;
         4'h597b 	:	val_out <= 4'he7cb;
         4'h5980 	:	val_out <= 4'he7bd;
         4'h5981 	:	val_out <= 4'he7bd;
         4'h5982 	:	val_out <= 4'he7bd;
         4'h5983 	:	val_out <= 4'he7bd;
         4'h5988 	:	val_out <= 4'he7ae;
         4'h5989 	:	val_out <= 4'he7ae;
         4'h598a 	:	val_out <= 4'he7ae;
         4'h598b 	:	val_out <= 4'he7ae;
         4'h5990 	:	val_out <= 4'he79f;
         4'h5991 	:	val_out <= 4'he79f;
         4'h5992 	:	val_out <= 4'he79f;
         4'h5993 	:	val_out <= 4'he79f;
         4'h5998 	:	val_out <= 4'he790;
         4'h5999 	:	val_out <= 4'he790;
         4'h599a 	:	val_out <= 4'he790;
         4'h599b 	:	val_out <= 4'he790;
         4'h59a0 	:	val_out <= 4'he782;
         4'h59a1 	:	val_out <= 4'he782;
         4'h59a2 	:	val_out <= 4'he782;
         4'h59a3 	:	val_out <= 4'he782;
         4'h59a8 	:	val_out <= 4'he773;
         4'h59a9 	:	val_out <= 4'he773;
         4'h59aa 	:	val_out <= 4'he773;
         4'h59ab 	:	val_out <= 4'he773;
         4'h59b0 	:	val_out <= 4'he764;
         4'h59b1 	:	val_out <= 4'he764;
         4'h59b2 	:	val_out <= 4'he764;
         4'h59b3 	:	val_out <= 4'he764;
         4'h59b8 	:	val_out <= 4'he755;
         4'h59b9 	:	val_out <= 4'he755;
         4'h59ba 	:	val_out <= 4'he755;
         4'h59bb 	:	val_out <= 4'he755;
         4'h59c0 	:	val_out <= 4'he746;
         4'h59c1 	:	val_out <= 4'he746;
         4'h59c2 	:	val_out <= 4'he746;
         4'h59c3 	:	val_out <= 4'he746;
         4'h59c8 	:	val_out <= 4'he737;
         4'h59c9 	:	val_out <= 4'he737;
         4'h59ca 	:	val_out <= 4'he737;
         4'h59cb 	:	val_out <= 4'he737;
         4'h59d0 	:	val_out <= 4'he729;
         4'h59d1 	:	val_out <= 4'he729;
         4'h59d2 	:	val_out <= 4'he729;
         4'h59d3 	:	val_out <= 4'he729;
         4'h59d8 	:	val_out <= 4'he71a;
         4'h59d9 	:	val_out <= 4'he71a;
         4'h59da 	:	val_out <= 4'he71a;
         4'h59db 	:	val_out <= 4'he71a;
         4'h59e0 	:	val_out <= 4'he70b;
         4'h59e1 	:	val_out <= 4'he70b;
         4'h59e2 	:	val_out <= 4'he70b;
         4'h59e3 	:	val_out <= 4'he70b;
         4'h59e8 	:	val_out <= 4'he6fc;
         4'h59e9 	:	val_out <= 4'he6fc;
         4'h59ea 	:	val_out <= 4'he6fc;
         4'h59eb 	:	val_out <= 4'he6fc;
         4'h59f0 	:	val_out <= 4'he6ed;
         4'h59f1 	:	val_out <= 4'he6ed;
         4'h59f2 	:	val_out <= 4'he6ed;
         4'h59f3 	:	val_out <= 4'he6ed;
         4'h59f8 	:	val_out <= 4'he6de;
         4'h59f9 	:	val_out <= 4'he6de;
         4'h59fa 	:	val_out <= 4'he6de;
         4'h59fb 	:	val_out <= 4'he6de;
         4'h5a00 	:	val_out <= 4'he6cf;
         4'h5a01 	:	val_out <= 4'he6cf;
         4'h5a02 	:	val_out <= 4'he6cf;
         4'h5a03 	:	val_out <= 4'he6cf;
         4'h5a08 	:	val_out <= 4'he6c0;
         4'h5a09 	:	val_out <= 4'he6c0;
         4'h5a0a 	:	val_out <= 4'he6c0;
         4'h5a0b 	:	val_out <= 4'he6c0;
         4'h5a10 	:	val_out <= 4'he6b1;
         4'h5a11 	:	val_out <= 4'he6b1;
         4'h5a12 	:	val_out <= 4'he6b1;
         4'h5a13 	:	val_out <= 4'he6b1;
         4'h5a18 	:	val_out <= 4'he6a2;
         4'h5a19 	:	val_out <= 4'he6a2;
         4'h5a1a 	:	val_out <= 4'he6a2;
         4'h5a1b 	:	val_out <= 4'he6a2;
         4'h5a20 	:	val_out <= 4'he693;
         4'h5a21 	:	val_out <= 4'he693;
         4'h5a22 	:	val_out <= 4'he693;
         4'h5a23 	:	val_out <= 4'he693;
         4'h5a28 	:	val_out <= 4'he684;
         4'h5a29 	:	val_out <= 4'he684;
         4'h5a2a 	:	val_out <= 4'he684;
         4'h5a2b 	:	val_out <= 4'he684;
         4'h5a30 	:	val_out <= 4'he675;
         4'h5a31 	:	val_out <= 4'he675;
         4'h5a32 	:	val_out <= 4'he675;
         4'h5a33 	:	val_out <= 4'he675;
         4'h5a38 	:	val_out <= 4'he666;
         4'h5a39 	:	val_out <= 4'he666;
         4'h5a3a 	:	val_out <= 4'he666;
         4'h5a3b 	:	val_out <= 4'he666;
         4'h5a40 	:	val_out <= 4'he657;
         4'h5a41 	:	val_out <= 4'he657;
         4'h5a42 	:	val_out <= 4'he657;
         4'h5a43 	:	val_out <= 4'he657;
         4'h5a48 	:	val_out <= 4'he648;
         4'h5a49 	:	val_out <= 4'he648;
         4'h5a4a 	:	val_out <= 4'he648;
         4'h5a4b 	:	val_out <= 4'he648;
         4'h5a50 	:	val_out <= 4'he639;
         4'h5a51 	:	val_out <= 4'he639;
         4'h5a52 	:	val_out <= 4'he639;
         4'h5a53 	:	val_out <= 4'he639;
         4'h5a58 	:	val_out <= 4'he629;
         4'h5a59 	:	val_out <= 4'he629;
         4'h5a5a 	:	val_out <= 4'he629;
         4'h5a5b 	:	val_out <= 4'he629;
         4'h5a60 	:	val_out <= 4'he61a;
         4'h5a61 	:	val_out <= 4'he61a;
         4'h5a62 	:	val_out <= 4'he61a;
         4'h5a63 	:	val_out <= 4'he61a;
         4'h5a68 	:	val_out <= 4'he60b;
         4'h5a69 	:	val_out <= 4'he60b;
         4'h5a6a 	:	val_out <= 4'he60b;
         4'h5a6b 	:	val_out <= 4'he60b;
         4'h5a70 	:	val_out <= 4'he5fc;
         4'h5a71 	:	val_out <= 4'he5fc;
         4'h5a72 	:	val_out <= 4'he5fc;
         4'h5a73 	:	val_out <= 4'he5fc;
         4'h5a78 	:	val_out <= 4'he5ed;
         4'h5a79 	:	val_out <= 4'he5ed;
         4'h5a7a 	:	val_out <= 4'he5ed;
         4'h5a7b 	:	val_out <= 4'he5ed;
         4'h5a80 	:	val_out <= 4'he5dd;
         4'h5a81 	:	val_out <= 4'he5dd;
         4'h5a82 	:	val_out <= 4'he5dd;
         4'h5a83 	:	val_out <= 4'he5dd;
         4'h5a88 	:	val_out <= 4'he5ce;
         4'h5a89 	:	val_out <= 4'he5ce;
         4'h5a8a 	:	val_out <= 4'he5ce;
         4'h5a8b 	:	val_out <= 4'he5ce;
         4'h5a90 	:	val_out <= 4'he5bf;
         4'h5a91 	:	val_out <= 4'he5bf;
         4'h5a92 	:	val_out <= 4'he5bf;
         4'h5a93 	:	val_out <= 4'he5bf;
         4'h5a98 	:	val_out <= 4'he5b0;
         4'h5a99 	:	val_out <= 4'he5b0;
         4'h5a9a 	:	val_out <= 4'he5b0;
         4'h5a9b 	:	val_out <= 4'he5b0;
         4'h5aa0 	:	val_out <= 4'he5a0;
         4'h5aa1 	:	val_out <= 4'he5a0;
         4'h5aa2 	:	val_out <= 4'he5a0;
         4'h5aa3 	:	val_out <= 4'he5a0;
         4'h5aa8 	:	val_out <= 4'he591;
         4'h5aa9 	:	val_out <= 4'he591;
         4'h5aaa 	:	val_out <= 4'he591;
         4'h5aab 	:	val_out <= 4'he591;
         4'h5ab0 	:	val_out <= 4'he582;
         4'h5ab1 	:	val_out <= 4'he582;
         4'h5ab2 	:	val_out <= 4'he582;
         4'h5ab3 	:	val_out <= 4'he582;
         4'h5ab8 	:	val_out <= 4'he573;
         4'h5ab9 	:	val_out <= 4'he573;
         4'h5aba 	:	val_out <= 4'he573;
         4'h5abb 	:	val_out <= 4'he573;
         4'h5ac0 	:	val_out <= 4'he563;
         4'h5ac1 	:	val_out <= 4'he563;
         4'h5ac2 	:	val_out <= 4'he563;
         4'h5ac3 	:	val_out <= 4'he563;
         4'h5ac8 	:	val_out <= 4'he554;
         4'h5ac9 	:	val_out <= 4'he554;
         4'h5aca 	:	val_out <= 4'he554;
         4'h5acb 	:	val_out <= 4'he554;
         4'h5ad0 	:	val_out <= 4'he545;
         4'h5ad1 	:	val_out <= 4'he545;
         4'h5ad2 	:	val_out <= 4'he545;
         4'h5ad3 	:	val_out <= 4'he545;
         4'h5ad8 	:	val_out <= 4'he535;
         4'h5ad9 	:	val_out <= 4'he535;
         4'h5ada 	:	val_out <= 4'he535;
         4'h5adb 	:	val_out <= 4'he535;
         4'h5ae0 	:	val_out <= 4'he526;
         4'h5ae1 	:	val_out <= 4'he526;
         4'h5ae2 	:	val_out <= 4'he526;
         4'h5ae3 	:	val_out <= 4'he526;
         4'h5ae8 	:	val_out <= 4'he516;
         4'h5ae9 	:	val_out <= 4'he516;
         4'h5aea 	:	val_out <= 4'he516;
         4'h5aeb 	:	val_out <= 4'he516;
         4'h5af0 	:	val_out <= 4'he507;
         4'h5af1 	:	val_out <= 4'he507;
         4'h5af2 	:	val_out <= 4'he507;
         4'h5af3 	:	val_out <= 4'he507;
         4'h5af8 	:	val_out <= 4'he4f7;
         4'h5af9 	:	val_out <= 4'he4f7;
         4'h5afa 	:	val_out <= 4'he4f7;
         4'h5afb 	:	val_out <= 4'he4f7;
         4'h5b00 	:	val_out <= 4'he4e8;
         4'h5b01 	:	val_out <= 4'he4e8;
         4'h5b02 	:	val_out <= 4'he4e8;
         4'h5b03 	:	val_out <= 4'he4e8;
         4'h5b08 	:	val_out <= 4'he4d9;
         4'h5b09 	:	val_out <= 4'he4d9;
         4'h5b0a 	:	val_out <= 4'he4d9;
         4'h5b0b 	:	val_out <= 4'he4d9;
         4'h5b10 	:	val_out <= 4'he4c9;
         4'h5b11 	:	val_out <= 4'he4c9;
         4'h5b12 	:	val_out <= 4'he4c9;
         4'h5b13 	:	val_out <= 4'he4c9;
         4'h5b18 	:	val_out <= 4'he4ba;
         4'h5b19 	:	val_out <= 4'he4ba;
         4'h5b1a 	:	val_out <= 4'he4ba;
         4'h5b1b 	:	val_out <= 4'he4ba;
         4'h5b20 	:	val_out <= 4'he4aa;
         4'h5b21 	:	val_out <= 4'he4aa;
         4'h5b22 	:	val_out <= 4'he4aa;
         4'h5b23 	:	val_out <= 4'he4aa;
         4'h5b28 	:	val_out <= 4'he49b;
         4'h5b29 	:	val_out <= 4'he49b;
         4'h5b2a 	:	val_out <= 4'he49b;
         4'h5b2b 	:	val_out <= 4'he49b;
         4'h5b30 	:	val_out <= 4'he48b;
         4'h5b31 	:	val_out <= 4'he48b;
         4'h5b32 	:	val_out <= 4'he48b;
         4'h5b33 	:	val_out <= 4'he48b;
         4'h5b38 	:	val_out <= 4'he47b;
         4'h5b39 	:	val_out <= 4'he47b;
         4'h5b3a 	:	val_out <= 4'he47b;
         4'h5b3b 	:	val_out <= 4'he47b;
         4'h5b40 	:	val_out <= 4'he46c;
         4'h5b41 	:	val_out <= 4'he46c;
         4'h5b42 	:	val_out <= 4'he46c;
         4'h5b43 	:	val_out <= 4'he46c;
         4'h5b48 	:	val_out <= 4'he45c;
         4'h5b49 	:	val_out <= 4'he45c;
         4'h5b4a 	:	val_out <= 4'he45c;
         4'h5b4b 	:	val_out <= 4'he45c;
         4'h5b50 	:	val_out <= 4'he44d;
         4'h5b51 	:	val_out <= 4'he44d;
         4'h5b52 	:	val_out <= 4'he44d;
         4'h5b53 	:	val_out <= 4'he44d;
         4'h5b58 	:	val_out <= 4'he43d;
         4'h5b59 	:	val_out <= 4'he43d;
         4'h5b5a 	:	val_out <= 4'he43d;
         4'h5b5b 	:	val_out <= 4'he43d;
         4'h5b60 	:	val_out <= 4'he42d;
         4'h5b61 	:	val_out <= 4'he42d;
         4'h5b62 	:	val_out <= 4'he42d;
         4'h5b63 	:	val_out <= 4'he42d;
         4'h5b68 	:	val_out <= 4'he41e;
         4'h5b69 	:	val_out <= 4'he41e;
         4'h5b6a 	:	val_out <= 4'he41e;
         4'h5b6b 	:	val_out <= 4'he41e;
         4'h5b70 	:	val_out <= 4'he40e;
         4'h5b71 	:	val_out <= 4'he40e;
         4'h5b72 	:	val_out <= 4'he40e;
         4'h5b73 	:	val_out <= 4'he40e;
         4'h5b78 	:	val_out <= 4'he3fe;
         4'h5b79 	:	val_out <= 4'he3fe;
         4'h5b7a 	:	val_out <= 4'he3fe;
         4'h5b7b 	:	val_out <= 4'he3fe;
         4'h5b80 	:	val_out <= 4'he3ef;
         4'h5b81 	:	val_out <= 4'he3ef;
         4'h5b82 	:	val_out <= 4'he3ef;
         4'h5b83 	:	val_out <= 4'he3ef;
         4'h5b88 	:	val_out <= 4'he3df;
         4'h5b89 	:	val_out <= 4'he3df;
         4'h5b8a 	:	val_out <= 4'he3df;
         4'h5b8b 	:	val_out <= 4'he3df;
         4'h5b90 	:	val_out <= 4'he3cf;
         4'h5b91 	:	val_out <= 4'he3cf;
         4'h5b92 	:	val_out <= 4'he3cf;
         4'h5b93 	:	val_out <= 4'he3cf;
         4'h5b98 	:	val_out <= 4'he3c0;
         4'h5b99 	:	val_out <= 4'he3c0;
         4'h5b9a 	:	val_out <= 4'he3c0;
         4'h5b9b 	:	val_out <= 4'he3c0;
         4'h5ba0 	:	val_out <= 4'he3b0;
         4'h5ba1 	:	val_out <= 4'he3b0;
         4'h5ba2 	:	val_out <= 4'he3b0;
         4'h5ba3 	:	val_out <= 4'he3b0;
         4'h5ba8 	:	val_out <= 4'he3a0;
         4'h5ba9 	:	val_out <= 4'he3a0;
         4'h5baa 	:	val_out <= 4'he3a0;
         4'h5bab 	:	val_out <= 4'he3a0;
         4'h5bb0 	:	val_out <= 4'he390;
         4'h5bb1 	:	val_out <= 4'he390;
         4'h5bb2 	:	val_out <= 4'he390;
         4'h5bb3 	:	val_out <= 4'he390;
         4'h5bb8 	:	val_out <= 4'he380;
         4'h5bb9 	:	val_out <= 4'he380;
         4'h5bba 	:	val_out <= 4'he380;
         4'h5bbb 	:	val_out <= 4'he380;
         4'h5bc0 	:	val_out <= 4'he371;
         4'h5bc1 	:	val_out <= 4'he371;
         4'h5bc2 	:	val_out <= 4'he371;
         4'h5bc3 	:	val_out <= 4'he371;
         4'h5bc8 	:	val_out <= 4'he361;
         4'h5bc9 	:	val_out <= 4'he361;
         4'h5bca 	:	val_out <= 4'he361;
         4'h5bcb 	:	val_out <= 4'he361;
         4'h5bd0 	:	val_out <= 4'he351;
         4'h5bd1 	:	val_out <= 4'he351;
         4'h5bd2 	:	val_out <= 4'he351;
         4'h5bd3 	:	val_out <= 4'he351;
         4'h5bd8 	:	val_out <= 4'he341;
         4'h5bd9 	:	val_out <= 4'he341;
         4'h5bda 	:	val_out <= 4'he341;
         4'h5bdb 	:	val_out <= 4'he341;
         4'h5be0 	:	val_out <= 4'he331;
         4'h5be1 	:	val_out <= 4'he331;
         4'h5be2 	:	val_out <= 4'he331;
         4'h5be3 	:	val_out <= 4'he331;
         4'h5be8 	:	val_out <= 4'he321;
         4'h5be9 	:	val_out <= 4'he321;
         4'h5bea 	:	val_out <= 4'he321;
         4'h5beb 	:	val_out <= 4'he321;
         4'h5bf0 	:	val_out <= 4'he311;
         4'h5bf1 	:	val_out <= 4'he311;
         4'h5bf2 	:	val_out <= 4'he311;
         4'h5bf3 	:	val_out <= 4'he311;
         4'h5bf8 	:	val_out <= 4'he301;
         4'h5bf9 	:	val_out <= 4'he301;
         4'h5bfa 	:	val_out <= 4'he301;
         4'h5bfb 	:	val_out <= 4'he301;
         4'h5c00 	:	val_out <= 4'he2f2;
         4'h5c01 	:	val_out <= 4'he2f2;
         4'h5c02 	:	val_out <= 4'he2f2;
         4'h5c03 	:	val_out <= 4'he2f2;
         4'h5c08 	:	val_out <= 4'he2e2;
         4'h5c09 	:	val_out <= 4'he2e2;
         4'h5c0a 	:	val_out <= 4'he2e2;
         4'h5c0b 	:	val_out <= 4'he2e2;
         4'h5c10 	:	val_out <= 4'he2d2;
         4'h5c11 	:	val_out <= 4'he2d2;
         4'h5c12 	:	val_out <= 4'he2d2;
         4'h5c13 	:	val_out <= 4'he2d2;
         4'h5c18 	:	val_out <= 4'he2c2;
         4'h5c19 	:	val_out <= 4'he2c2;
         4'h5c1a 	:	val_out <= 4'he2c2;
         4'h5c1b 	:	val_out <= 4'he2c2;
         4'h5c20 	:	val_out <= 4'he2b2;
         4'h5c21 	:	val_out <= 4'he2b2;
         4'h5c22 	:	val_out <= 4'he2b2;
         4'h5c23 	:	val_out <= 4'he2b2;
         4'h5c28 	:	val_out <= 4'he2a2;
         4'h5c29 	:	val_out <= 4'he2a2;
         4'h5c2a 	:	val_out <= 4'he2a2;
         4'h5c2b 	:	val_out <= 4'he2a2;
         4'h5c30 	:	val_out <= 4'he292;
         4'h5c31 	:	val_out <= 4'he292;
         4'h5c32 	:	val_out <= 4'he292;
         4'h5c33 	:	val_out <= 4'he292;
         4'h5c38 	:	val_out <= 4'he282;
         4'h5c39 	:	val_out <= 4'he282;
         4'h5c3a 	:	val_out <= 4'he282;
         4'h5c3b 	:	val_out <= 4'he282;
         4'h5c40 	:	val_out <= 4'he271;
         4'h5c41 	:	val_out <= 4'he271;
         4'h5c42 	:	val_out <= 4'he271;
         4'h5c43 	:	val_out <= 4'he271;
         4'h5c48 	:	val_out <= 4'he261;
         4'h5c49 	:	val_out <= 4'he261;
         4'h5c4a 	:	val_out <= 4'he261;
         4'h5c4b 	:	val_out <= 4'he261;
         4'h5c50 	:	val_out <= 4'he251;
         4'h5c51 	:	val_out <= 4'he251;
         4'h5c52 	:	val_out <= 4'he251;
         4'h5c53 	:	val_out <= 4'he251;
         4'h5c58 	:	val_out <= 4'he241;
         4'h5c59 	:	val_out <= 4'he241;
         4'h5c5a 	:	val_out <= 4'he241;
         4'h5c5b 	:	val_out <= 4'he241;
         4'h5c60 	:	val_out <= 4'he231;
         4'h5c61 	:	val_out <= 4'he231;
         4'h5c62 	:	val_out <= 4'he231;
         4'h5c63 	:	val_out <= 4'he231;
         4'h5c68 	:	val_out <= 4'he221;
         4'h5c69 	:	val_out <= 4'he221;
         4'h5c6a 	:	val_out <= 4'he221;
         4'h5c6b 	:	val_out <= 4'he221;
         4'h5c70 	:	val_out <= 4'he211;
         4'h5c71 	:	val_out <= 4'he211;
         4'h5c72 	:	val_out <= 4'he211;
         4'h5c73 	:	val_out <= 4'he211;
         4'h5c78 	:	val_out <= 4'he201;
         4'h5c79 	:	val_out <= 4'he201;
         4'h5c7a 	:	val_out <= 4'he201;
         4'h5c7b 	:	val_out <= 4'he201;
         4'h5c80 	:	val_out <= 4'he1f1;
         4'h5c81 	:	val_out <= 4'he1f1;
         4'h5c82 	:	val_out <= 4'he1f1;
         4'h5c83 	:	val_out <= 4'he1f1;
         4'h5c88 	:	val_out <= 4'he1e0;
         4'h5c89 	:	val_out <= 4'he1e0;
         4'h5c8a 	:	val_out <= 4'he1e0;
         4'h5c8b 	:	val_out <= 4'he1e0;
         4'h5c90 	:	val_out <= 4'he1d0;
         4'h5c91 	:	val_out <= 4'he1d0;
         4'h5c92 	:	val_out <= 4'he1d0;
         4'h5c93 	:	val_out <= 4'he1d0;
         4'h5c98 	:	val_out <= 4'he1c0;
         4'h5c99 	:	val_out <= 4'he1c0;
         4'h5c9a 	:	val_out <= 4'he1c0;
         4'h5c9b 	:	val_out <= 4'he1c0;
         4'h5ca0 	:	val_out <= 4'he1b0;
         4'h5ca1 	:	val_out <= 4'he1b0;
         4'h5ca2 	:	val_out <= 4'he1b0;
         4'h5ca3 	:	val_out <= 4'he1b0;
         4'h5ca8 	:	val_out <= 4'he19f;
         4'h5ca9 	:	val_out <= 4'he19f;
         4'h5caa 	:	val_out <= 4'he19f;
         4'h5cab 	:	val_out <= 4'he19f;
         4'h5cb0 	:	val_out <= 4'he18f;
         4'h5cb1 	:	val_out <= 4'he18f;
         4'h5cb2 	:	val_out <= 4'he18f;
         4'h5cb3 	:	val_out <= 4'he18f;
         4'h5cb8 	:	val_out <= 4'he17f;
         4'h5cb9 	:	val_out <= 4'he17f;
         4'h5cba 	:	val_out <= 4'he17f;
         4'h5cbb 	:	val_out <= 4'he17f;
         4'h5cc0 	:	val_out <= 4'he16f;
         4'h5cc1 	:	val_out <= 4'he16f;
         4'h5cc2 	:	val_out <= 4'he16f;
         4'h5cc3 	:	val_out <= 4'he16f;
         4'h5cc8 	:	val_out <= 4'he15e;
         4'h5cc9 	:	val_out <= 4'he15e;
         4'h5cca 	:	val_out <= 4'he15e;
         4'h5ccb 	:	val_out <= 4'he15e;
         4'h5cd0 	:	val_out <= 4'he14e;
         4'h5cd1 	:	val_out <= 4'he14e;
         4'h5cd2 	:	val_out <= 4'he14e;
         4'h5cd3 	:	val_out <= 4'he14e;
         4'h5cd8 	:	val_out <= 4'he13e;
         4'h5cd9 	:	val_out <= 4'he13e;
         4'h5cda 	:	val_out <= 4'he13e;
         4'h5cdb 	:	val_out <= 4'he13e;
         4'h5ce0 	:	val_out <= 4'he12d;
         4'h5ce1 	:	val_out <= 4'he12d;
         4'h5ce2 	:	val_out <= 4'he12d;
         4'h5ce3 	:	val_out <= 4'he12d;
         4'h5ce8 	:	val_out <= 4'he11d;
         4'h5ce9 	:	val_out <= 4'he11d;
         4'h5cea 	:	val_out <= 4'he11d;
         4'h5ceb 	:	val_out <= 4'he11d;
         4'h5cf0 	:	val_out <= 4'he10d;
         4'h5cf1 	:	val_out <= 4'he10d;
         4'h5cf2 	:	val_out <= 4'he10d;
         4'h5cf3 	:	val_out <= 4'he10d;
         4'h5cf8 	:	val_out <= 4'he0fc;
         4'h5cf9 	:	val_out <= 4'he0fc;
         4'h5cfa 	:	val_out <= 4'he0fc;
         4'h5cfb 	:	val_out <= 4'he0fc;
         4'h5d00 	:	val_out <= 4'he0ec;
         4'h5d01 	:	val_out <= 4'he0ec;
         4'h5d02 	:	val_out <= 4'he0ec;
         4'h5d03 	:	val_out <= 4'he0ec;
         4'h5d08 	:	val_out <= 4'he0db;
         4'h5d09 	:	val_out <= 4'he0db;
         4'h5d0a 	:	val_out <= 4'he0db;
         4'h5d0b 	:	val_out <= 4'he0db;
         4'h5d10 	:	val_out <= 4'he0cb;
         4'h5d11 	:	val_out <= 4'he0cb;
         4'h5d12 	:	val_out <= 4'he0cb;
         4'h5d13 	:	val_out <= 4'he0cb;
         4'h5d18 	:	val_out <= 4'he0ba;
         4'h5d19 	:	val_out <= 4'he0ba;
         4'h5d1a 	:	val_out <= 4'he0ba;
         4'h5d1b 	:	val_out <= 4'he0ba;
         4'h5d20 	:	val_out <= 4'he0aa;
         4'h5d21 	:	val_out <= 4'he0aa;
         4'h5d22 	:	val_out <= 4'he0aa;
         4'h5d23 	:	val_out <= 4'he0aa;
         4'h5d28 	:	val_out <= 4'he099;
         4'h5d29 	:	val_out <= 4'he099;
         4'h5d2a 	:	val_out <= 4'he099;
         4'h5d2b 	:	val_out <= 4'he099;
         4'h5d30 	:	val_out <= 4'he089;
         4'h5d31 	:	val_out <= 4'he089;
         4'h5d32 	:	val_out <= 4'he089;
         4'h5d33 	:	val_out <= 4'he089;
         4'h5d38 	:	val_out <= 4'he078;
         4'h5d39 	:	val_out <= 4'he078;
         4'h5d3a 	:	val_out <= 4'he078;
         4'h5d3b 	:	val_out <= 4'he078;
         4'h5d40 	:	val_out <= 4'he068;
         4'h5d41 	:	val_out <= 4'he068;
         4'h5d42 	:	val_out <= 4'he068;
         4'h5d43 	:	val_out <= 4'he068;
         4'h5d48 	:	val_out <= 4'he057;
         4'h5d49 	:	val_out <= 4'he057;
         4'h5d4a 	:	val_out <= 4'he057;
         4'h5d4b 	:	val_out <= 4'he057;
         4'h5d50 	:	val_out <= 4'he047;
         4'h5d51 	:	val_out <= 4'he047;
         4'h5d52 	:	val_out <= 4'he047;
         4'h5d53 	:	val_out <= 4'he047;
         4'h5d58 	:	val_out <= 4'he036;
         4'h5d59 	:	val_out <= 4'he036;
         4'h5d5a 	:	val_out <= 4'he036;
         4'h5d5b 	:	val_out <= 4'he036;
         4'h5d60 	:	val_out <= 4'he026;
         4'h5d61 	:	val_out <= 4'he026;
         4'h5d62 	:	val_out <= 4'he026;
         4'h5d63 	:	val_out <= 4'he026;
         4'h5d68 	:	val_out <= 4'he015;
         4'h5d69 	:	val_out <= 4'he015;
         4'h5d6a 	:	val_out <= 4'he015;
         4'h5d6b 	:	val_out <= 4'he015;
         4'h5d70 	:	val_out <= 4'he004;
         4'h5d71 	:	val_out <= 4'he004;
         4'h5d72 	:	val_out <= 4'he004;
         4'h5d73 	:	val_out <= 4'he004;
         4'h5d78 	:	val_out <= 4'hdff4;
         4'h5d79 	:	val_out <= 4'hdff4;
         4'h5d7a 	:	val_out <= 4'hdff4;
         4'h5d7b 	:	val_out <= 4'hdff4;
         4'h5d80 	:	val_out <= 4'hdfe3;
         4'h5d81 	:	val_out <= 4'hdfe3;
         4'h5d82 	:	val_out <= 4'hdfe3;
         4'h5d83 	:	val_out <= 4'hdfe3;
         4'h5d88 	:	val_out <= 4'hdfd3;
         4'h5d89 	:	val_out <= 4'hdfd3;
         4'h5d8a 	:	val_out <= 4'hdfd3;
         4'h5d8b 	:	val_out <= 4'hdfd3;
         4'h5d90 	:	val_out <= 4'hdfc2;
         4'h5d91 	:	val_out <= 4'hdfc2;
         4'h5d92 	:	val_out <= 4'hdfc2;
         4'h5d93 	:	val_out <= 4'hdfc2;
         4'h5d98 	:	val_out <= 4'hdfb1;
         4'h5d99 	:	val_out <= 4'hdfb1;
         4'h5d9a 	:	val_out <= 4'hdfb1;
         4'h5d9b 	:	val_out <= 4'hdfb1;
         4'h5da0 	:	val_out <= 4'hdfa0;
         4'h5da1 	:	val_out <= 4'hdfa0;
         4'h5da2 	:	val_out <= 4'hdfa0;
         4'h5da3 	:	val_out <= 4'hdfa0;
         4'h5da8 	:	val_out <= 4'hdf90;
         4'h5da9 	:	val_out <= 4'hdf90;
         4'h5daa 	:	val_out <= 4'hdf90;
         4'h5dab 	:	val_out <= 4'hdf90;
         4'h5db0 	:	val_out <= 4'hdf7f;
         4'h5db1 	:	val_out <= 4'hdf7f;
         4'h5db2 	:	val_out <= 4'hdf7f;
         4'h5db3 	:	val_out <= 4'hdf7f;
         4'h5db8 	:	val_out <= 4'hdf6e;
         4'h5db9 	:	val_out <= 4'hdf6e;
         4'h5dba 	:	val_out <= 4'hdf6e;
         4'h5dbb 	:	val_out <= 4'hdf6e;
         4'h5dc0 	:	val_out <= 4'hdf5e;
         4'h5dc1 	:	val_out <= 4'hdf5e;
         4'h5dc2 	:	val_out <= 4'hdf5e;
         4'h5dc3 	:	val_out <= 4'hdf5e;
         4'h5dc8 	:	val_out <= 4'hdf4d;
         4'h5dc9 	:	val_out <= 4'hdf4d;
         4'h5dca 	:	val_out <= 4'hdf4d;
         4'h5dcb 	:	val_out <= 4'hdf4d;
         4'h5dd0 	:	val_out <= 4'hdf3c;
         4'h5dd1 	:	val_out <= 4'hdf3c;
         4'h5dd2 	:	val_out <= 4'hdf3c;
         4'h5dd3 	:	val_out <= 4'hdf3c;
         4'h5dd8 	:	val_out <= 4'hdf2b;
         4'h5dd9 	:	val_out <= 4'hdf2b;
         4'h5dda 	:	val_out <= 4'hdf2b;
         4'h5ddb 	:	val_out <= 4'hdf2b;
         4'h5de0 	:	val_out <= 4'hdf1a;
         4'h5de1 	:	val_out <= 4'hdf1a;
         4'h5de2 	:	val_out <= 4'hdf1a;
         4'h5de3 	:	val_out <= 4'hdf1a;
         4'h5de8 	:	val_out <= 4'hdf0a;
         4'h5de9 	:	val_out <= 4'hdf0a;
         4'h5dea 	:	val_out <= 4'hdf0a;
         4'h5deb 	:	val_out <= 4'hdf0a;
         4'h5df0 	:	val_out <= 4'hdef9;
         4'h5df1 	:	val_out <= 4'hdef9;
         4'h5df2 	:	val_out <= 4'hdef9;
         4'h5df3 	:	val_out <= 4'hdef9;
         4'h5df8 	:	val_out <= 4'hdee8;
         4'h5df9 	:	val_out <= 4'hdee8;
         4'h5dfa 	:	val_out <= 4'hdee8;
         4'h5dfb 	:	val_out <= 4'hdee8;
         4'h5e00 	:	val_out <= 4'hded7;
         4'h5e01 	:	val_out <= 4'hded7;
         4'h5e02 	:	val_out <= 4'hded7;
         4'h5e03 	:	val_out <= 4'hded7;
         4'h5e08 	:	val_out <= 4'hdec6;
         4'h5e09 	:	val_out <= 4'hdec6;
         4'h5e0a 	:	val_out <= 4'hdec6;
         4'h5e0b 	:	val_out <= 4'hdec6;
         4'h5e10 	:	val_out <= 4'hdeb5;
         4'h5e11 	:	val_out <= 4'hdeb5;
         4'h5e12 	:	val_out <= 4'hdeb5;
         4'h5e13 	:	val_out <= 4'hdeb5;
         4'h5e18 	:	val_out <= 4'hdea4;
         4'h5e19 	:	val_out <= 4'hdea4;
         4'h5e1a 	:	val_out <= 4'hdea4;
         4'h5e1b 	:	val_out <= 4'hdea4;
         4'h5e20 	:	val_out <= 4'hde93;
         4'h5e21 	:	val_out <= 4'hde93;
         4'h5e22 	:	val_out <= 4'hde93;
         4'h5e23 	:	val_out <= 4'hde93;
         4'h5e28 	:	val_out <= 4'hde82;
         4'h5e29 	:	val_out <= 4'hde82;
         4'h5e2a 	:	val_out <= 4'hde82;
         4'h5e2b 	:	val_out <= 4'hde82;
         4'h5e30 	:	val_out <= 4'hde71;
         4'h5e31 	:	val_out <= 4'hde71;
         4'h5e32 	:	val_out <= 4'hde71;
         4'h5e33 	:	val_out <= 4'hde71;
         4'h5e38 	:	val_out <= 4'hde60;
         4'h5e39 	:	val_out <= 4'hde60;
         4'h5e3a 	:	val_out <= 4'hde60;
         4'h5e3b 	:	val_out <= 4'hde60;
         4'h5e40 	:	val_out <= 4'hde50;
         4'h5e41 	:	val_out <= 4'hde50;
         4'h5e42 	:	val_out <= 4'hde50;
         4'h5e43 	:	val_out <= 4'hde50;
         4'h5e48 	:	val_out <= 4'hde3f;
         4'h5e49 	:	val_out <= 4'hde3f;
         4'h5e4a 	:	val_out <= 4'hde3f;
         4'h5e4b 	:	val_out <= 4'hde3f;
         4'h5e50 	:	val_out <= 4'hde2d;
         4'h5e51 	:	val_out <= 4'hde2d;
         4'h5e52 	:	val_out <= 4'hde2d;
         4'h5e53 	:	val_out <= 4'hde2d;
         4'h5e58 	:	val_out <= 4'hde1c;
         4'h5e59 	:	val_out <= 4'hde1c;
         4'h5e5a 	:	val_out <= 4'hde1c;
         4'h5e5b 	:	val_out <= 4'hde1c;
         4'h5e60 	:	val_out <= 4'hde0b;
         4'h5e61 	:	val_out <= 4'hde0b;
         4'h5e62 	:	val_out <= 4'hde0b;
         4'h5e63 	:	val_out <= 4'hde0b;
         4'h5e68 	:	val_out <= 4'hddfa;
         4'h5e69 	:	val_out <= 4'hddfa;
         4'h5e6a 	:	val_out <= 4'hddfa;
         4'h5e6b 	:	val_out <= 4'hddfa;
         4'h5e70 	:	val_out <= 4'hdde9;
         4'h5e71 	:	val_out <= 4'hdde9;
         4'h5e72 	:	val_out <= 4'hdde9;
         4'h5e73 	:	val_out <= 4'hdde9;
         4'h5e78 	:	val_out <= 4'hddd8;
         4'h5e79 	:	val_out <= 4'hddd8;
         4'h5e7a 	:	val_out <= 4'hddd8;
         4'h5e7b 	:	val_out <= 4'hddd8;
         4'h5e80 	:	val_out <= 4'hddc7;
         4'h5e81 	:	val_out <= 4'hddc7;
         4'h5e82 	:	val_out <= 4'hddc7;
         4'h5e83 	:	val_out <= 4'hddc7;
         4'h5e88 	:	val_out <= 4'hddb6;
         4'h5e89 	:	val_out <= 4'hddb6;
         4'h5e8a 	:	val_out <= 4'hddb6;
         4'h5e8b 	:	val_out <= 4'hddb6;
         4'h5e90 	:	val_out <= 4'hdda5;
         4'h5e91 	:	val_out <= 4'hdda5;
         4'h5e92 	:	val_out <= 4'hdda5;
         4'h5e93 	:	val_out <= 4'hdda5;
         4'h5e98 	:	val_out <= 4'hdd94;
         4'h5e99 	:	val_out <= 4'hdd94;
         4'h5e9a 	:	val_out <= 4'hdd94;
         4'h5e9b 	:	val_out <= 4'hdd94;
         4'h5ea0 	:	val_out <= 4'hdd83;
         4'h5ea1 	:	val_out <= 4'hdd83;
         4'h5ea2 	:	val_out <= 4'hdd83;
         4'h5ea3 	:	val_out <= 4'hdd83;
         4'h5ea8 	:	val_out <= 4'hdd71;
         4'h5ea9 	:	val_out <= 4'hdd71;
         4'h5eaa 	:	val_out <= 4'hdd71;
         4'h5eab 	:	val_out <= 4'hdd71;
         4'h5eb0 	:	val_out <= 4'hdd60;
         4'h5eb1 	:	val_out <= 4'hdd60;
         4'h5eb2 	:	val_out <= 4'hdd60;
         4'h5eb3 	:	val_out <= 4'hdd60;
         4'h5eb8 	:	val_out <= 4'hdd4f;
         4'h5eb9 	:	val_out <= 4'hdd4f;
         4'h5eba 	:	val_out <= 4'hdd4f;
         4'h5ebb 	:	val_out <= 4'hdd4f;
         4'h5ec0 	:	val_out <= 4'hdd3e;
         4'h5ec1 	:	val_out <= 4'hdd3e;
         4'h5ec2 	:	val_out <= 4'hdd3e;
         4'h5ec3 	:	val_out <= 4'hdd3e;
         4'h5ec8 	:	val_out <= 4'hdd2d;
         4'h5ec9 	:	val_out <= 4'hdd2d;
         4'h5eca 	:	val_out <= 4'hdd2d;
         4'h5ecb 	:	val_out <= 4'hdd2d;
         4'h5ed0 	:	val_out <= 4'hdd1b;
         4'h5ed1 	:	val_out <= 4'hdd1b;
         4'h5ed2 	:	val_out <= 4'hdd1b;
         4'h5ed3 	:	val_out <= 4'hdd1b;
         4'h5ed8 	:	val_out <= 4'hdd0a;
         4'h5ed9 	:	val_out <= 4'hdd0a;
         4'h5eda 	:	val_out <= 4'hdd0a;
         4'h5edb 	:	val_out <= 4'hdd0a;
         4'h5ee0 	:	val_out <= 4'hdcf9;
         4'h5ee1 	:	val_out <= 4'hdcf9;
         4'h5ee2 	:	val_out <= 4'hdcf9;
         4'h5ee3 	:	val_out <= 4'hdcf9;
         4'h5ee8 	:	val_out <= 4'hdce8;
         4'h5ee9 	:	val_out <= 4'hdce8;
         4'h5eea 	:	val_out <= 4'hdce8;
         4'h5eeb 	:	val_out <= 4'hdce8;
         4'h5ef0 	:	val_out <= 4'hdcd6;
         4'h5ef1 	:	val_out <= 4'hdcd6;
         4'h5ef2 	:	val_out <= 4'hdcd6;
         4'h5ef3 	:	val_out <= 4'hdcd6;
         4'h5ef8 	:	val_out <= 4'hdcc5;
         4'h5ef9 	:	val_out <= 4'hdcc5;
         4'h5efa 	:	val_out <= 4'hdcc5;
         4'h5efb 	:	val_out <= 4'hdcc5;
         4'h5f00 	:	val_out <= 4'hdcb4;
         4'h5f01 	:	val_out <= 4'hdcb4;
         4'h5f02 	:	val_out <= 4'hdcb4;
         4'h5f03 	:	val_out <= 4'hdcb4;
         4'h5f08 	:	val_out <= 4'hdca2;
         4'h5f09 	:	val_out <= 4'hdca2;
         4'h5f0a 	:	val_out <= 4'hdca2;
         4'h5f0b 	:	val_out <= 4'hdca2;
         4'h5f10 	:	val_out <= 4'hdc91;
         4'h5f11 	:	val_out <= 4'hdc91;
         4'h5f12 	:	val_out <= 4'hdc91;
         4'h5f13 	:	val_out <= 4'hdc91;
         4'h5f18 	:	val_out <= 4'hdc80;
         4'h5f19 	:	val_out <= 4'hdc80;
         4'h5f1a 	:	val_out <= 4'hdc80;
         4'h5f1b 	:	val_out <= 4'hdc80;
         4'h5f20 	:	val_out <= 4'hdc6e;
         4'h5f21 	:	val_out <= 4'hdc6e;
         4'h5f22 	:	val_out <= 4'hdc6e;
         4'h5f23 	:	val_out <= 4'hdc6e;
         4'h5f28 	:	val_out <= 4'hdc5d;
         4'h5f29 	:	val_out <= 4'hdc5d;
         4'h5f2a 	:	val_out <= 4'hdc5d;
         4'h5f2b 	:	val_out <= 4'hdc5d;
         4'h5f30 	:	val_out <= 4'hdc4b;
         4'h5f31 	:	val_out <= 4'hdc4b;
         4'h5f32 	:	val_out <= 4'hdc4b;
         4'h5f33 	:	val_out <= 4'hdc4b;
         4'h5f38 	:	val_out <= 4'hdc3a;
         4'h5f39 	:	val_out <= 4'hdc3a;
         4'h5f3a 	:	val_out <= 4'hdc3a;
         4'h5f3b 	:	val_out <= 4'hdc3a;
         4'h5f40 	:	val_out <= 4'hdc29;
         4'h5f41 	:	val_out <= 4'hdc29;
         4'h5f42 	:	val_out <= 4'hdc29;
         4'h5f43 	:	val_out <= 4'hdc29;
         4'h5f48 	:	val_out <= 4'hdc17;
         4'h5f49 	:	val_out <= 4'hdc17;
         4'h5f4a 	:	val_out <= 4'hdc17;
         4'h5f4b 	:	val_out <= 4'hdc17;
         4'h5f50 	:	val_out <= 4'hdc06;
         4'h5f51 	:	val_out <= 4'hdc06;
         4'h5f52 	:	val_out <= 4'hdc06;
         4'h5f53 	:	val_out <= 4'hdc06;
         4'h5f58 	:	val_out <= 4'hdbf4;
         4'h5f59 	:	val_out <= 4'hdbf4;
         4'h5f5a 	:	val_out <= 4'hdbf4;
         4'h5f5b 	:	val_out <= 4'hdbf4;
         4'h5f60 	:	val_out <= 4'hdbe3;
         4'h5f61 	:	val_out <= 4'hdbe3;
         4'h5f62 	:	val_out <= 4'hdbe3;
         4'h5f63 	:	val_out <= 4'hdbe3;
         4'h5f68 	:	val_out <= 4'hdbd1;
         4'h5f69 	:	val_out <= 4'hdbd1;
         4'h5f6a 	:	val_out <= 4'hdbd1;
         4'h5f6b 	:	val_out <= 4'hdbd1;
         4'h5f70 	:	val_out <= 4'hdbc0;
         4'h5f71 	:	val_out <= 4'hdbc0;
         4'h5f72 	:	val_out <= 4'hdbc0;
         4'h5f73 	:	val_out <= 4'hdbc0;
         4'h5f78 	:	val_out <= 4'hdbae;
         4'h5f79 	:	val_out <= 4'hdbae;
         4'h5f7a 	:	val_out <= 4'hdbae;
         4'h5f7b 	:	val_out <= 4'hdbae;
         4'h5f80 	:	val_out <= 4'hdb9d;
         4'h5f81 	:	val_out <= 4'hdb9d;
         4'h5f82 	:	val_out <= 4'hdb9d;
         4'h5f83 	:	val_out <= 4'hdb9d;
         4'h5f88 	:	val_out <= 4'hdb8b;
         4'h5f89 	:	val_out <= 4'hdb8b;
         4'h5f8a 	:	val_out <= 4'hdb8b;
         4'h5f8b 	:	val_out <= 4'hdb8b;
         4'h5f90 	:	val_out <= 4'hdb79;
         4'h5f91 	:	val_out <= 4'hdb79;
         4'h5f92 	:	val_out <= 4'hdb79;
         4'h5f93 	:	val_out <= 4'hdb79;
         4'h5f98 	:	val_out <= 4'hdb68;
         4'h5f99 	:	val_out <= 4'hdb68;
         4'h5f9a 	:	val_out <= 4'hdb68;
         4'h5f9b 	:	val_out <= 4'hdb68;
         4'h5fa0 	:	val_out <= 4'hdb56;
         4'h5fa1 	:	val_out <= 4'hdb56;
         4'h5fa2 	:	val_out <= 4'hdb56;
         4'h5fa3 	:	val_out <= 4'hdb56;
         4'h5fa8 	:	val_out <= 4'hdb45;
         4'h5fa9 	:	val_out <= 4'hdb45;
         4'h5faa 	:	val_out <= 4'hdb45;
         4'h5fab 	:	val_out <= 4'hdb45;
         4'h5fb0 	:	val_out <= 4'hdb33;
         4'h5fb1 	:	val_out <= 4'hdb33;
         4'h5fb2 	:	val_out <= 4'hdb33;
         4'h5fb3 	:	val_out <= 4'hdb33;
         4'h5fb8 	:	val_out <= 4'hdb21;
         4'h5fb9 	:	val_out <= 4'hdb21;
         4'h5fba 	:	val_out <= 4'hdb21;
         4'h5fbb 	:	val_out <= 4'hdb21;
         4'h5fc0 	:	val_out <= 4'hdb10;
         4'h5fc1 	:	val_out <= 4'hdb10;
         4'h5fc2 	:	val_out <= 4'hdb10;
         4'h5fc3 	:	val_out <= 4'hdb10;
         4'h5fc8 	:	val_out <= 4'hdafe;
         4'h5fc9 	:	val_out <= 4'hdafe;
         4'h5fca 	:	val_out <= 4'hdafe;
         4'h5fcb 	:	val_out <= 4'hdafe;
         4'h5fd0 	:	val_out <= 4'hdaec;
         4'h5fd1 	:	val_out <= 4'hdaec;
         4'h5fd2 	:	val_out <= 4'hdaec;
         4'h5fd3 	:	val_out <= 4'hdaec;
         4'h5fd8 	:	val_out <= 4'hdadb;
         4'h5fd9 	:	val_out <= 4'hdadb;
         4'h5fda 	:	val_out <= 4'hdadb;
         4'h5fdb 	:	val_out <= 4'hdadb;
         4'h5fe0 	:	val_out <= 4'hdac9;
         4'h5fe1 	:	val_out <= 4'hdac9;
         4'h5fe2 	:	val_out <= 4'hdac9;
         4'h5fe3 	:	val_out <= 4'hdac9;
         4'h5fe8 	:	val_out <= 4'hdab7;
         4'h5fe9 	:	val_out <= 4'hdab7;
         4'h5fea 	:	val_out <= 4'hdab7;
         4'h5feb 	:	val_out <= 4'hdab7;
         4'h5ff0 	:	val_out <= 4'hdaa5;
         4'h5ff1 	:	val_out <= 4'hdaa5;
         4'h5ff2 	:	val_out <= 4'hdaa5;
         4'h5ff3 	:	val_out <= 4'hdaa5;
         4'h5ff8 	:	val_out <= 4'hda94;
         4'h5ff9 	:	val_out <= 4'hda94;
         4'h5ffa 	:	val_out <= 4'hda94;
         4'h5ffb 	:	val_out <= 4'hda94;
         4'h6000 	:	val_out <= 4'hda82;
         4'h6001 	:	val_out <= 4'hda82;
         4'h6002 	:	val_out <= 4'hda82;
         4'h6003 	:	val_out <= 4'hda82;
         4'h6008 	:	val_out <= 4'hda70;
         4'h6009 	:	val_out <= 4'hda70;
         4'h600a 	:	val_out <= 4'hda70;
         4'h600b 	:	val_out <= 4'hda70;
         4'h6010 	:	val_out <= 4'hda5e;
         4'h6011 	:	val_out <= 4'hda5e;
         4'h6012 	:	val_out <= 4'hda5e;
         4'h6013 	:	val_out <= 4'hda5e;
         4'h6018 	:	val_out <= 4'hda4d;
         4'h6019 	:	val_out <= 4'hda4d;
         4'h601a 	:	val_out <= 4'hda4d;
         4'h601b 	:	val_out <= 4'hda4d;
         4'h6020 	:	val_out <= 4'hda3b;
         4'h6021 	:	val_out <= 4'hda3b;
         4'h6022 	:	val_out <= 4'hda3b;
         4'h6023 	:	val_out <= 4'hda3b;
         4'h6028 	:	val_out <= 4'hda29;
         4'h6029 	:	val_out <= 4'hda29;
         4'h602a 	:	val_out <= 4'hda29;
         4'h602b 	:	val_out <= 4'hda29;
         4'h6030 	:	val_out <= 4'hda17;
         4'h6031 	:	val_out <= 4'hda17;
         4'h6032 	:	val_out <= 4'hda17;
         4'h6033 	:	val_out <= 4'hda17;
         4'h6038 	:	val_out <= 4'hda05;
         4'h6039 	:	val_out <= 4'hda05;
         4'h603a 	:	val_out <= 4'hda05;
         4'h603b 	:	val_out <= 4'hda05;
         4'h6040 	:	val_out <= 4'hd9f3;
         4'h6041 	:	val_out <= 4'hd9f3;
         4'h6042 	:	val_out <= 4'hd9f3;
         4'h6043 	:	val_out <= 4'hd9f3;
         4'h6048 	:	val_out <= 4'hd9e1;
         4'h6049 	:	val_out <= 4'hd9e1;
         4'h604a 	:	val_out <= 4'hd9e1;
         4'h604b 	:	val_out <= 4'hd9e1;
         4'h6050 	:	val_out <= 4'hd9d0;
         4'h6051 	:	val_out <= 4'hd9d0;
         4'h6052 	:	val_out <= 4'hd9d0;
         4'h6053 	:	val_out <= 4'hd9d0;
         4'h6058 	:	val_out <= 4'hd9be;
         4'h6059 	:	val_out <= 4'hd9be;
         4'h605a 	:	val_out <= 4'hd9be;
         4'h605b 	:	val_out <= 4'hd9be;
         4'h6060 	:	val_out <= 4'hd9ac;
         4'h6061 	:	val_out <= 4'hd9ac;
         4'h6062 	:	val_out <= 4'hd9ac;
         4'h6063 	:	val_out <= 4'hd9ac;
         4'h6068 	:	val_out <= 4'hd99a;
         4'h6069 	:	val_out <= 4'hd99a;
         4'h606a 	:	val_out <= 4'hd99a;
         4'h606b 	:	val_out <= 4'hd99a;
         4'h6070 	:	val_out <= 4'hd988;
         4'h6071 	:	val_out <= 4'hd988;
         4'h6072 	:	val_out <= 4'hd988;
         4'h6073 	:	val_out <= 4'hd988;
         4'h6078 	:	val_out <= 4'hd976;
         4'h6079 	:	val_out <= 4'hd976;
         4'h607a 	:	val_out <= 4'hd976;
         4'h607b 	:	val_out <= 4'hd976;
         4'h6080 	:	val_out <= 4'hd964;
         4'h6081 	:	val_out <= 4'hd964;
         4'h6082 	:	val_out <= 4'hd964;
         4'h6083 	:	val_out <= 4'hd964;
         4'h6088 	:	val_out <= 4'hd952;
         4'h6089 	:	val_out <= 4'hd952;
         4'h608a 	:	val_out <= 4'hd952;
         4'h608b 	:	val_out <= 4'hd952;
         4'h6090 	:	val_out <= 4'hd940;
         4'h6091 	:	val_out <= 4'hd940;
         4'h6092 	:	val_out <= 4'hd940;
         4'h6093 	:	val_out <= 4'hd940;
         4'h6098 	:	val_out <= 4'hd92e;
         4'h6099 	:	val_out <= 4'hd92e;
         4'h609a 	:	val_out <= 4'hd92e;
         4'h609b 	:	val_out <= 4'hd92e;
         4'h60a0 	:	val_out <= 4'hd91c;
         4'h60a1 	:	val_out <= 4'hd91c;
         4'h60a2 	:	val_out <= 4'hd91c;
         4'h60a3 	:	val_out <= 4'hd91c;
         4'h60a8 	:	val_out <= 4'hd90a;
         4'h60a9 	:	val_out <= 4'hd90a;
         4'h60aa 	:	val_out <= 4'hd90a;
         4'h60ab 	:	val_out <= 4'hd90a;
         4'h60b0 	:	val_out <= 4'hd8f8;
         4'h60b1 	:	val_out <= 4'hd8f8;
         4'h60b2 	:	val_out <= 4'hd8f8;
         4'h60b3 	:	val_out <= 4'hd8f8;
         4'h60b8 	:	val_out <= 4'hd8e6;
         4'h60b9 	:	val_out <= 4'hd8e6;
         4'h60ba 	:	val_out <= 4'hd8e6;
         4'h60bb 	:	val_out <= 4'hd8e6;
         4'h60c0 	:	val_out <= 4'hd8d4;
         4'h60c1 	:	val_out <= 4'hd8d4;
         4'h60c2 	:	val_out <= 4'hd8d4;
         4'h60c3 	:	val_out <= 4'hd8d4;
         4'h60c8 	:	val_out <= 4'hd8c1;
         4'h60c9 	:	val_out <= 4'hd8c1;
         4'h60ca 	:	val_out <= 4'hd8c1;
         4'h60cb 	:	val_out <= 4'hd8c1;
         4'h60d0 	:	val_out <= 4'hd8af;
         4'h60d1 	:	val_out <= 4'hd8af;
         4'h60d2 	:	val_out <= 4'hd8af;
         4'h60d3 	:	val_out <= 4'hd8af;
         4'h60d8 	:	val_out <= 4'hd89d;
         4'h60d9 	:	val_out <= 4'hd89d;
         4'h60da 	:	val_out <= 4'hd89d;
         4'h60db 	:	val_out <= 4'hd89d;
         4'h60e0 	:	val_out <= 4'hd88b;
         4'h60e1 	:	val_out <= 4'hd88b;
         4'h60e2 	:	val_out <= 4'hd88b;
         4'h60e3 	:	val_out <= 4'hd88b;
         4'h60e8 	:	val_out <= 4'hd879;
         4'h60e9 	:	val_out <= 4'hd879;
         4'h60ea 	:	val_out <= 4'hd879;
         4'h60eb 	:	val_out <= 4'hd879;
         4'h60f0 	:	val_out <= 4'hd867;
         4'h60f1 	:	val_out <= 4'hd867;
         4'h60f2 	:	val_out <= 4'hd867;
         4'h60f3 	:	val_out <= 4'hd867;
         4'h60f8 	:	val_out <= 4'hd855;
         4'h60f9 	:	val_out <= 4'hd855;
         4'h60fa 	:	val_out <= 4'hd855;
         4'h60fb 	:	val_out <= 4'hd855;
         4'h6100 	:	val_out <= 4'hd842;
         4'h6101 	:	val_out <= 4'hd842;
         4'h6102 	:	val_out <= 4'hd842;
         4'h6103 	:	val_out <= 4'hd842;
         4'h6108 	:	val_out <= 4'hd830;
         4'h6109 	:	val_out <= 4'hd830;
         4'h610a 	:	val_out <= 4'hd830;
         4'h610b 	:	val_out <= 4'hd830;
         4'h6110 	:	val_out <= 4'hd81e;
         4'h6111 	:	val_out <= 4'hd81e;
         4'h6112 	:	val_out <= 4'hd81e;
         4'h6113 	:	val_out <= 4'hd81e;
         4'h6118 	:	val_out <= 4'hd80c;
         4'h6119 	:	val_out <= 4'hd80c;
         4'h611a 	:	val_out <= 4'hd80c;
         4'h611b 	:	val_out <= 4'hd80c;
         4'h6120 	:	val_out <= 4'hd7f9;
         4'h6121 	:	val_out <= 4'hd7f9;
         4'h6122 	:	val_out <= 4'hd7f9;
         4'h6123 	:	val_out <= 4'hd7f9;
         4'h6128 	:	val_out <= 4'hd7e7;
         4'h6129 	:	val_out <= 4'hd7e7;
         4'h612a 	:	val_out <= 4'hd7e7;
         4'h612b 	:	val_out <= 4'hd7e7;
         4'h6130 	:	val_out <= 4'hd7d5;
         4'h6131 	:	val_out <= 4'hd7d5;
         4'h6132 	:	val_out <= 4'hd7d5;
         4'h6133 	:	val_out <= 4'hd7d5;
         4'h6138 	:	val_out <= 4'hd7c3;
         4'h6139 	:	val_out <= 4'hd7c3;
         4'h613a 	:	val_out <= 4'hd7c3;
         4'h613b 	:	val_out <= 4'hd7c3;
         4'h6140 	:	val_out <= 4'hd7b0;
         4'h6141 	:	val_out <= 4'hd7b0;
         4'h6142 	:	val_out <= 4'hd7b0;
         4'h6143 	:	val_out <= 4'hd7b0;
         4'h6148 	:	val_out <= 4'hd79e;
         4'h6149 	:	val_out <= 4'hd79e;
         4'h614a 	:	val_out <= 4'hd79e;
         4'h614b 	:	val_out <= 4'hd79e;
         4'h6150 	:	val_out <= 4'hd78c;
         4'h6151 	:	val_out <= 4'hd78c;
         4'h6152 	:	val_out <= 4'hd78c;
         4'h6153 	:	val_out <= 4'hd78c;
         4'h6158 	:	val_out <= 4'hd779;
         4'h6159 	:	val_out <= 4'hd779;
         4'h615a 	:	val_out <= 4'hd779;
         4'h615b 	:	val_out <= 4'hd779;
         4'h6160 	:	val_out <= 4'hd767;
         4'h6161 	:	val_out <= 4'hd767;
         4'h6162 	:	val_out <= 4'hd767;
         4'h6163 	:	val_out <= 4'hd767;
         4'h6168 	:	val_out <= 4'hd755;
         4'h6169 	:	val_out <= 4'hd755;
         4'h616a 	:	val_out <= 4'hd755;
         4'h616b 	:	val_out <= 4'hd755;
         4'h6170 	:	val_out <= 4'hd742;
         4'h6171 	:	val_out <= 4'hd742;
         4'h6172 	:	val_out <= 4'hd742;
         4'h6173 	:	val_out <= 4'hd742;
         4'h6178 	:	val_out <= 4'hd730;
         4'h6179 	:	val_out <= 4'hd730;
         4'h617a 	:	val_out <= 4'hd730;
         4'h617b 	:	val_out <= 4'hd730;
         4'h6180 	:	val_out <= 4'hd71d;
         4'h6181 	:	val_out <= 4'hd71d;
         4'h6182 	:	val_out <= 4'hd71d;
         4'h6183 	:	val_out <= 4'hd71d;
         4'h6188 	:	val_out <= 4'hd70b;
         4'h6189 	:	val_out <= 4'hd70b;
         4'h618a 	:	val_out <= 4'hd70b;
         4'h618b 	:	val_out <= 4'hd70b;
         4'h6190 	:	val_out <= 4'hd6f9;
         4'h6191 	:	val_out <= 4'hd6f9;
         4'h6192 	:	val_out <= 4'hd6f9;
         4'h6193 	:	val_out <= 4'hd6f9;
         4'h6198 	:	val_out <= 4'hd6e6;
         4'h6199 	:	val_out <= 4'hd6e6;
         4'h619a 	:	val_out <= 4'hd6e6;
         4'h619b 	:	val_out <= 4'hd6e6;
         4'h61a0 	:	val_out <= 4'hd6d4;
         4'h61a1 	:	val_out <= 4'hd6d4;
         4'h61a2 	:	val_out <= 4'hd6d4;
         4'h61a3 	:	val_out <= 4'hd6d4;
         4'h61a8 	:	val_out <= 4'hd6c1;
         4'h61a9 	:	val_out <= 4'hd6c1;
         4'h61aa 	:	val_out <= 4'hd6c1;
         4'h61ab 	:	val_out <= 4'hd6c1;
         4'h61b0 	:	val_out <= 4'hd6af;
         4'h61b1 	:	val_out <= 4'hd6af;
         4'h61b2 	:	val_out <= 4'hd6af;
         4'h61b3 	:	val_out <= 4'hd6af;
         4'h61b8 	:	val_out <= 4'hd69c;
         4'h61b9 	:	val_out <= 4'hd69c;
         4'h61ba 	:	val_out <= 4'hd69c;
         4'h61bb 	:	val_out <= 4'hd69c;
         4'h61c0 	:	val_out <= 4'hd68a;
         4'h61c1 	:	val_out <= 4'hd68a;
         4'h61c2 	:	val_out <= 4'hd68a;
         4'h61c3 	:	val_out <= 4'hd68a;
         4'h61c8 	:	val_out <= 4'hd677;
         4'h61c9 	:	val_out <= 4'hd677;
         4'h61ca 	:	val_out <= 4'hd677;
         4'h61cb 	:	val_out <= 4'hd677;
         4'h61d0 	:	val_out <= 4'hd665;
         4'h61d1 	:	val_out <= 4'hd665;
         4'h61d2 	:	val_out <= 4'hd665;
         4'h61d3 	:	val_out <= 4'hd665;
         4'h61d8 	:	val_out <= 4'hd652;
         4'h61d9 	:	val_out <= 4'hd652;
         4'h61da 	:	val_out <= 4'hd652;
         4'h61db 	:	val_out <= 4'hd652;
         4'h61e0 	:	val_out <= 4'hd640;
         4'h61e1 	:	val_out <= 4'hd640;
         4'h61e2 	:	val_out <= 4'hd640;
         4'h61e3 	:	val_out <= 4'hd640;
         4'h61e8 	:	val_out <= 4'hd62d;
         4'h61e9 	:	val_out <= 4'hd62d;
         4'h61ea 	:	val_out <= 4'hd62d;
         4'h61eb 	:	val_out <= 4'hd62d;
         4'h61f0 	:	val_out <= 4'hd61a;
         4'h61f1 	:	val_out <= 4'hd61a;
         4'h61f2 	:	val_out <= 4'hd61a;
         4'h61f3 	:	val_out <= 4'hd61a;
         4'h61f8 	:	val_out <= 4'hd608;
         4'h61f9 	:	val_out <= 4'hd608;
         4'h61fa 	:	val_out <= 4'hd608;
         4'h61fb 	:	val_out <= 4'hd608;
         4'h6200 	:	val_out <= 4'hd5f5;
         4'h6201 	:	val_out <= 4'hd5f5;
         4'h6202 	:	val_out <= 4'hd5f5;
         4'h6203 	:	val_out <= 4'hd5f5;
         4'h6208 	:	val_out <= 4'hd5e3;
         4'h6209 	:	val_out <= 4'hd5e3;
         4'h620a 	:	val_out <= 4'hd5e3;
         4'h620b 	:	val_out <= 4'hd5e3;
         4'h6210 	:	val_out <= 4'hd5d0;
         4'h6211 	:	val_out <= 4'hd5d0;
         4'h6212 	:	val_out <= 4'hd5d0;
         4'h6213 	:	val_out <= 4'hd5d0;
         4'h6218 	:	val_out <= 4'hd5bd;
         4'h6219 	:	val_out <= 4'hd5bd;
         4'h621a 	:	val_out <= 4'hd5bd;
         4'h621b 	:	val_out <= 4'hd5bd;
         4'h6220 	:	val_out <= 4'hd5ab;
         4'h6221 	:	val_out <= 4'hd5ab;
         4'h6222 	:	val_out <= 4'hd5ab;
         4'h6223 	:	val_out <= 4'hd5ab;
         4'h6228 	:	val_out <= 4'hd598;
         4'h6229 	:	val_out <= 4'hd598;
         4'h622a 	:	val_out <= 4'hd598;
         4'h622b 	:	val_out <= 4'hd598;
         4'h6230 	:	val_out <= 4'hd585;
         4'h6231 	:	val_out <= 4'hd585;
         4'h6232 	:	val_out <= 4'hd585;
         4'h6233 	:	val_out <= 4'hd585;
         4'h6238 	:	val_out <= 4'hd572;
         4'h6239 	:	val_out <= 4'hd572;
         4'h623a 	:	val_out <= 4'hd572;
         4'h623b 	:	val_out <= 4'hd572;
         4'h6240 	:	val_out <= 4'hd560;
         4'h6241 	:	val_out <= 4'hd560;
         4'h6242 	:	val_out <= 4'hd560;
         4'h6243 	:	val_out <= 4'hd560;
         4'h6248 	:	val_out <= 4'hd54d;
         4'h6249 	:	val_out <= 4'hd54d;
         4'h624a 	:	val_out <= 4'hd54d;
         4'h624b 	:	val_out <= 4'hd54d;
         4'h6250 	:	val_out <= 4'hd53a;
         4'h6251 	:	val_out <= 4'hd53a;
         4'h6252 	:	val_out <= 4'hd53a;
         4'h6253 	:	val_out <= 4'hd53a;
         4'h6258 	:	val_out <= 4'hd528;
         4'h6259 	:	val_out <= 4'hd528;
         4'h625a 	:	val_out <= 4'hd528;
         4'h625b 	:	val_out <= 4'hd528;
         4'h6260 	:	val_out <= 4'hd515;
         4'h6261 	:	val_out <= 4'hd515;
         4'h6262 	:	val_out <= 4'hd515;
         4'h6263 	:	val_out <= 4'hd515;
         4'h6268 	:	val_out <= 4'hd502;
         4'h6269 	:	val_out <= 4'hd502;
         4'h626a 	:	val_out <= 4'hd502;
         4'h626b 	:	val_out <= 4'hd502;
         4'h6270 	:	val_out <= 4'hd4ef;
         4'h6271 	:	val_out <= 4'hd4ef;
         4'h6272 	:	val_out <= 4'hd4ef;
         4'h6273 	:	val_out <= 4'hd4ef;
         4'h6278 	:	val_out <= 4'hd4dc;
         4'h6279 	:	val_out <= 4'hd4dc;
         4'h627a 	:	val_out <= 4'hd4dc;
         4'h627b 	:	val_out <= 4'hd4dc;
         4'h6280 	:	val_out <= 4'hd4ca;
         4'h6281 	:	val_out <= 4'hd4ca;
         4'h6282 	:	val_out <= 4'hd4ca;
         4'h6283 	:	val_out <= 4'hd4ca;
         4'h6288 	:	val_out <= 4'hd4b7;
         4'h6289 	:	val_out <= 4'hd4b7;
         4'h628a 	:	val_out <= 4'hd4b7;
         4'h628b 	:	val_out <= 4'hd4b7;
         4'h6290 	:	val_out <= 4'hd4a4;
         4'h6291 	:	val_out <= 4'hd4a4;
         4'h6292 	:	val_out <= 4'hd4a4;
         4'h6293 	:	val_out <= 4'hd4a4;
         4'h6298 	:	val_out <= 4'hd491;
         4'h6299 	:	val_out <= 4'hd491;
         4'h629a 	:	val_out <= 4'hd491;
         4'h629b 	:	val_out <= 4'hd491;
         4'h62a0 	:	val_out <= 4'hd47e;
         4'h62a1 	:	val_out <= 4'hd47e;
         4'h62a2 	:	val_out <= 4'hd47e;
         4'h62a3 	:	val_out <= 4'hd47e;
         4'h62a8 	:	val_out <= 4'hd46b;
         4'h62a9 	:	val_out <= 4'hd46b;
         4'h62aa 	:	val_out <= 4'hd46b;
         4'h62ab 	:	val_out <= 4'hd46b;
         4'h62b0 	:	val_out <= 4'hd458;
         4'h62b1 	:	val_out <= 4'hd458;
         4'h62b2 	:	val_out <= 4'hd458;
         4'h62b3 	:	val_out <= 4'hd458;
         4'h62b8 	:	val_out <= 4'hd445;
         4'h62b9 	:	val_out <= 4'hd445;
         4'h62ba 	:	val_out <= 4'hd445;
         4'h62bb 	:	val_out <= 4'hd445;
         4'h62c0 	:	val_out <= 4'hd433;
         4'h62c1 	:	val_out <= 4'hd433;
         4'h62c2 	:	val_out <= 4'hd433;
         4'h62c3 	:	val_out <= 4'hd433;
         4'h62c8 	:	val_out <= 4'hd420;
         4'h62c9 	:	val_out <= 4'hd420;
         4'h62ca 	:	val_out <= 4'hd420;
         4'h62cb 	:	val_out <= 4'hd420;
         4'h62d0 	:	val_out <= 4'hd40d;
         4'h62d1 	:	val_out <= 4'hd40d;
         4'h62d2 	:	val_out <= 4'hd40d;
         4'h62d3 	:	val_out <= 4'hd40d;
         4'h62d8 	:	val_out <= 4'hd3fa;
         4'h62d9 	:	val_out <= 4'hd3fa;
         4'h62da 	:	val_out <= 4'hd3fa;
         4'h62db 	:	val_out <= 4'hd3fa;
         4'h62e0 	:	val_out <= 4'hd3e7;
         4'h62e1 	:	val_out <= 4'hd3e7;
         4'h62e2 	:	val_out <= 4'hd3e7;
         4'h62e3 	:	val_out <= 4'hd3e7;
         4'h62e8 	:	val_out <= 4'hd3d4;
         4'h62e9 	:	val_out <= 4'hd3d4;
         4'h62ea 	:	val_out <= 4'hd3d4;
         4'h62eb 	:	val_out <= 4'hd3d4;
         4'h62f0 	:	val_out <= 4'hd3c1;
         4'h62f1 	:	val_out <= 4'hd3c1;
         4'h62f2 	:	val_out <= 4'hd3c1;
         4'h62f3 	:	val_out <= 4'hd3c1;
         4'h62f8 	:	val_out <= 4'hd3ae;
         4'h62f9 	:	val_out <= 4'hd3ae;
         4'h62fa 	:	val_out <= 4'hd3ae;
         4'h62fb 	:	val_out <= 4'hd3ae;
         4'h6300 	:	val_out <= 4'hd39b;
         4'h6301 	:	val_out <= 4'hd39b;
         4'h6302 	:	val_out <= 4'hd39b;
         4'h6303 	:	val_out <= 4'hd39b;
         4'h6308 	:	val_out <= 4'hd388;
         4'h6309 	:	val_out <= 4'hd388;
         4'h630a 	:	val_out <= 4'hd388;
         4'h630b 	:	val_out <= 4'hd388;
         4'h6310 	:	val_out <= 4'hd375;
         4'h6311 	:	val_out <= 4'hd375;
         4'h6312 	:	val_out <= 4'hd375;
         4'h6313 	:	val_out <= 4'hd375;
         4'h6318 	:	val_out <= 4'hd362;
         4'h6319 	:	val_out <= 4'hd362;
         4'h631a 	:	val_out <= 4'hd362;
         4'h631b 	:	val_out <= 4'hd362;
         4'h6320 	:	val_out <= 4'hd34e;
         4'h6321 	:	val_out <= 4'hd34e;
         4'h6322 	:	val_out <= 4'hd34e;
         4'h6323 	:	val_out <= 4'hd34e;
         4'h6328 	:	val_out <= 4'hd33b;
         4'h6329 	:	val_out <= 4'hd33b;
         4'h632a 	:	val_out <= 4'hd33b;
         4'h632b 	:	val_out <= 4'hd33b;
         4'h6330 	:	val_out <= 4'hd328;
         4'h6331 	:	val_out <= 4'hd328;
         4'h6332 	:	val_out <= 4'hd328;
         4'h6333 	:	val_out <= 4'hd328;
         4'h6338 	:	val_out <= 4'hd315;
         4'h6339 	:	val_out <= 4'hd315;
         4'h633a 	:	val_out <= 4'hd315;
         4'h633b 	:	val_out <= 4'hd315;
         4'h6340 	:	val_out <= 4'hd302;
         4'h6341 	:	val_out <= 4'hd302;
         4'h6342 	:	val_out <= 4'hd302;
         4'h6343 	:	val_out <= 4'hd302;
         4'h6348 	:	val_out <= 4'hd2ef;
         4'h6349 	:	val_out <= 4'hd2ef;
         4'h634a 	:	val_out <= 4'hd2ef;
         4'h634b 	:	val_out <= 4'hd2ef;
         4'h6350 	:	val_out <= 4'hd2dc;
         4'h6351 	:	val_out <= 4'hd2dc;
         4'h6352 	:	val_out <= 4'hd2dc;
         4'h6353 	:	val_out <= 4'hd2dc;
         4'h6358 	:	val_out <= 4'hd2c9;
         4'h6359 	:	val_out <= 4'hd2c9;
         4'h635a 	:	val_out <= 4'hd2c9;
         4'h635b 	:	val_out <= 4'hd2c9;
         4'h6360 	:	val_out <= 4'hd2b5;
         4'h6361 	:	val_out <= 4'hd2b5;
         4'h6362 	:	val_out <= 4'hd2b5;
         4'h6363 	:	val_out <= 4'hd2b5;
         4'h6368 	:	val_out <= 4'hd2a2;
         4'h6369 	:	val_out <= 4'hd2a2;
         4'h636a 	:	val_out <= 4'hd2a2;
         4'h636b 	:	val_out <= 4'hd2a2;
         4'h6370 	:	val_out <= 4'hd28f;
         4'h6371 	:	val_out <= 4'hd28f;
         4'h6372 	:	val_out <= 4'hd28f;
         4'h6373 	:	val_out <= 4'hd28f;
         4'h6378 	:	val_out <= 4'hd27c;
         4'h6379 	:	val_out <= 4'hd27c;
         4'h637a 	:	val_out <= 4'hd27c;
         4'h637b 	:	val_out <= 4'hd27c;
         4'h6380 	:	val_out <= 4'hd269;
         4'h6381 	:	val_out <= 4'hd269;
         4'h6382 	:	val_out <= 4'hd269;
         4'h6383 	:	val_out <= 4'hd269;
         4'h6388 	:	val_out <= 4'hd255;
         4'h6389 	:	val_out <= 4'hd255;
         4'h638a 	:	val_out <= 4'hd255;
         4'h638b 	:	val_out <= 4'hd255;
         4'h6390 	:	val_out <= 4'hd242;
         4'h6391 	:	val_out <= 4'hd242;
         4'h6392 	:	val_out <= 4'hd242;
         4'h6393 	:	val_out <= 4'hd242;
         4'h6398 	:	val_out <= 4'hd22f;
         4'h6399 	:	val_out <= 4'hd22f;
         4'h639a 	:	val_out <= 4'hd22f;
         4'h639b 	:	val_out <= 4'hd22f;
         4'h63a0 	:	val_out <= 4'hd21c;
         4'h63a1 	:	val_out <= 4'hd21c;
         4'h63a2 	:	val_out <= 4'hd21c;
         4'h63a3 	:	val_out <= 4'hd21c;
         4'h63a8 	:	val_out <= 4'hd208;
         4'h63a9 	:	val_out <= 4'hd208;
         4'h63aa 	:	val_out <= 4'hd208;
         4'h63ab 	:	val_out <= 4'hd208;
         4'h63b0 	:	val_out <= 4'hd1f5;
         4'h63b1 	:	val_out <= 4'hd1f5;
         4'h63b2 	:	val_out <= 4'hd1f5;
         4'h63b3 	:	val_out <= 4'hd1f5;
         4'h63b8 	:	val_out <= 4'hd1e2;
         4'h63b9 	:	val_out <= 4'hd1e2;
         4'h63ba 	:	val_out <= 4'hd1e2;
         4'h63bb 	:	val_out <= 4'hd1e2;
         4'h63c0 	:	val_out <= 4'hd1ce;
         4'h63c1 	:	val_out <= 4'hd1ce;
         4'h63c2 	:	val_out <= 4'hd1ce;
         4'h63c3 	:	val_out <= 4'hd1ce;
         4'h63c8 	:	val_out <= 4'hd1bb;
         4'h63c9 	:	val_out <= 4'hd1bb;
         4'h63ca 	:	val_out <= 4'hd1bb;
         4'h63cb 	:	val_out <= 4'hd1bb;
         4'h63d0 	:	val_out <= 4'hd1a8;
         4'h63d1 	:	val_out <= 4'hd1a8;
         4'h63d2 	:	val_out <= 4'hd1a8;
         4'h63d3 	:	val_out <= 4'hd1a8;
         4'h63d8 	:	val_out <= 4'hd194;
         4'h63d9 	:	val_out <= 4'hd194;
         4'h63da 	:	val_out <= 4'hd194;
         4'h63db 	:	val_out <= 4'hd194;
         4'h63e0 	:	val_out <= 4'hd181;
         4'h63e1 	:	val_out <= 4'hd181;
         4'h63e2 	:	val_out <= 4'hd181;
         4'h63e3 	:	val_out <= 4'hd181;
         4'h63e8 	:	val_out <= 4'hd16e;
         4'h63e9 	:	val_out <= 4'hd16e;
         4'h63ea 	:	val_out <= 4'hd16e;
         4'h63eb 	:	val_out <= 4'hd16e;
         4'h63f0 	:	val_out <= 4'hd15a;
         4'h63f1 	:	val_out <= 4'hd15a;
         4'h63f2 	:	val_out <= 4'hd15a;
         4'h63f3 	:	val_out <= 4'hd15a;
         4'h63f8 	:	val_out <= 4'hd147;
         4'h63f9 	:	val_out <= 4'hd147;
         4'h63fa 	:	val_out <= 4'hd147;
         4'h63fb 	:	val_out <= 4'hd147;
         4'h6400 	:	val_out <= 4'hd133;
         4'h6401 	:	val_out <= 4'hd133;
         4'h6402 	:	val_out <= 4'hd133;
         4'h6403 	:	val_out <= 4'hd133;
         4'h6408 	:	val_out <= 4'hd120;
         4'h6409 	:	val_out <= 4'hd120;
         4'h640a 	:	val_out <= 4'hd120;
         4'h640b 	:	val_out <= 4'hd120;
         4'h6410 	:	val_out <= 4'hd10c;
         4'h6411 	:	val_out <= 4'hd10c;
         4'h6412 	:	val_out <= 4'hd10c;
         4'h6413 	:	val_out <= 4'hd10c;
         4'h6418 	:	val_out <= 4'hd0f9;
         4'h6419 	:	val_out <= 4'hd0f9;
         4'h641a 	:	val_out <= 4'hd0f9;
         4'h641b 	:	val_out <= 4'hd0f9;
         4'h6420 	:	val_out <= 4'hd0e5;
         4'h6421 	:	val_out <= 4'hd0e5;
         4'h6422 	:	val_out <= 4'hd0e5;
         4'h6423 	:	val_out <= 4'hd0e5;
         4'h6428 	:	val_out <= 4'hd0d2;
         4'h6429 	:	val_out <= 4'hd0d2;
         4'h642a 	:	val_out <= 4'hd0d2;
         4'h642b 	:	val_out <= 4'hd0d2;
         4'h6430 	:	val_out <= 4'hd0bf;
         4'h6431 	:	val_out <= 4'hd0bf;
         4'h6432 	:	val_out <= 4'hd0bf;
         4'h6433 	:	val_out <= 4'hd0bf;
         4'h6438 	:	val_out <= 4'hd0ab;
         4'h6439 	:	val_out <= 4'hd0ab;
         4'h643a 	:	val_out <= 4'hd0ab;
         4'h643b 	:	val_out <= 4'hd0ab;
         4'h6440 	:	val_out <= 4'hd097;
         4'h6441 	:	val_out <= 4'hd097;
         4'h6442 	:	val_out <= 4'hd097;
         4'h6443 	:	val_out <= 4'hd097;
         4'h6448 	:	val_out <= 4'hd084;
         4'h6449 	:	val_out <= 4'hd084;
         4'h644a 	:	val_out <= 4'hd084;
         4'h644b 	:	val_out <= 4'hd084;
         4'h6450 	:	val_out <= 4'hd070;
         4'h6451 	:	val_out <= 4'hd070;
         4'h6452 	:	val_out <= 4'hd070;
         4'h6453 	:	val_out <= 4'hd070;
         4'h6458 	:	val_out <= 4'hd05d;
         4'h6459 	:	val_out <= 4'hd05d;
         4'h645a 	:	val_out <= 4'hd05d;
         4'h645b 	:	val_out <= 4'hd05d;
         4'h6460 	:	val_out <= 4'hd049;
         4'h6461 	:	val_out <= 4'hd049;
         4'h6462 	:	val_out <= 4'hd049;
         4'h6463 	:	val_out <= 4'hd049;
         4'h6468 	:	val_out <= 4'hd036;
         4'h6469 	:	val_out <= 4'hd036;
         4'h646a 	:	val_out <= 4'hd036;
         4'h646b 	:	val_out <= 4'hd036;
         4'h6470 	:	val_out <= 4'hd022;
         4'h6471 	:	val_out <= 4'hd022;
         4'h6472 	:	val_out <= 4'hd022;
         4'h6473 	:	val_out <= 4'hd022;
         4'h6478 	:	val_out <= 4'hd00f;
         4'h6479 	:	val_out <= 4'hd00f;
         4'h647a 	:	val_out <= 4'hd00f;
         4'h647b 	:	val_out <= 4'hd00f;
         4'h6480 	:	val_out <= 4'hcffb;
         4'h6481 	:	val_out <= 4'hcffb;
         4'h6482 	:	val_out <= 4'hcffb;
         4'h6483 	:	val_out <= 4'hcffb;
         4'h6488 	:	val_out <= 4'hcfe7;
         4'h6489 	:	val_out <= 4'hcfe7;
         4'h648a 	:	val_out <= 4'hcfe7;
         4'h648b 	:	val_out <= 4'hcfe7;
         4'h6490 	:	val_out <= 4'hcfd4;
         4'h6491 	:	val_out <= 4'hcfd4;
         4'h6492 	:	val_out <= 4'hcfd4;
         4'h6493 	:	val_out <= 4'hcfd4;
         4'h6498 	:	val_out <= 4'hcfc0;
         4'h6499 	:	val_out <= 4'hcfc0;
         4'h649a 	:	val_out <= 4'hcfc0;
         4'h649b 	:	val_out <= 4'hcfc0;
         4'h64a0 	:	val_out <= 4'hcfac;
         4'h64a1 	:	val_out <= 4'hcfac;
         4'h64a2 	:	val_out <= 4'hcfac;
         4'h64a3 	:	val_out <= 4'hcfac;
         4'h64a8 	:	val_out <= 4'hcf99;
         4'h64a9 	:	val_out <= 4'hcf99;
         4'h64aa 	:	val_out <= 4'hcf99;
         4'h64ab 	:	val_out <= 4'hcf99;
         4'h64b0 	:	val_out <= 4'hcf85;
         4'h64b1 	:	val_out <= 4'hcf85;
         4'h64b2 	:	val_out <= 4'hcf85;
         4'h64b3 	:	val_out <= 4'hcf85;
         4'h64b8 	:	val_out <= 4'hcf71;
         4'h64b9 	:	val_out <= 4'hcf71;
         4'h64ba 	:	val_out <= 4'hcf71;
         4'h64bb 	:	val_out <= 4'hcf71;
         4'h64c0 	:	val_out <= 4'hcf5e;
         4'h64c1 	:	val_out <= 4'hcf5e;
         4'h64c2 	:	val_out <= 4'hcf5e;
         4'h64c3 	:	val_out <= 4'hcf5e;
         4'h64c8 	:	val_out <= 4'hcf4a;
         4'h64c9 	:	val_out <= 4'hcf4a;
         4'h64ca 	:	val_out <= 4'hcf4a;
         4'h64cb 	:	val_out <= 4'hcf4a;
         4'h64d0 	:	val_out <= 4'hcf36;
         4'h64d1 	:	val_out <= 4'hcf36;
         4'h64d2 	:	val_out <= 4'hcf36;
         4'h64d3 	:	val_out <= 4'hcf36;
         4'h64d8 	:	val_out <= 4'hcf22;
         4'h64d9 	:	val_out <= 4'hcf22;
         4'h64da 	:	val_out <= 4'hcf22;
         4'h64db 	:	val_out <= 4'hcf22;
         4'h64e0 	:	val_out <= 4'hcf0f;
         4'h64e1 	:	val_out <= 4'hcf0f;
         4'h64e2 	:	val_out <= 4'hcf0f;
         4'h64e3 	:	val_out <= 4'hcf0f;
         4'h64e8 	:	val_out <= 4'hcefb;
         4'h64e9 	:	val_out <= 4'hcefb;
         4'h64ea 	:	val_out <= 4'hcefb;
         4'h64eb 	:	val_out <= 4'hcefb;
         4'h64f0 	:	val_out <= 4'hcee7;
         4'h64f1 	:	val_out <= 4'hcee7;
         4'h64f2 	:	val_out <= 4'hcee7;
         4'h64f3 	:	val_out <= 4'hcee7;
         4'h64f8 	:	val_out <= 4'hced3;
         4'h64f9 	:	val_out <= 4'hced3;
         4'h64fa 	:	val_out <= 4'hced3;
         4'h64fb 	:	val_out <= 4'hced3;
         4'h6500 	:	val_out <= 4'hcebf;
         4'h6501 	:	val_out <= 4'hcebf;
         4'h6502 	:	val_out <= 4'hcebf;
         4'h6503 	:	val_out <= 4'hcebf;
         4'h6508 	:	val_out <= 4'hceac;
         4'h6509 	:	val_out <= 4'hceac;
         4'h650a 	:	val_out <= 4'hceac;
         4'h650b 	:	val_out <= 4'hceac;
         4'h6510 	:	val_out <= 4'hce98;
         4'h6511 	:	val_out <= 4'hce98;
         4'h6512 	:	val_out <= 4'hce98;
         4'h6513 	:	val_out <= 4'hce98;
         4'h6518 	:	val_out <= 4'hce84;
         4'h6519 	:	val_out <= 4'hce84;
         4'h651a 	:	val_out <= 4'hce84;
         4'h651b 	:	val_out <= 4'hce84;
         4'h6520 	:	val_out <= 4'hce70;
         4'h6521 	:	val_out <= 4'hce70;
         4'h6522 	:	val_out <= 4'hce70;
         4'h6523 	:	val_out <= 4'hce70;
         4'h6528 	:	val_out <= 4'hce5c;
         4'h6529 	:	val_out <= 4'hce5c;
         4'h652a 	:	val_out <= 4'hce5c;
         4'h652b 	:	val_out <= 4'hce5c;
         4'h6530 	:	val_out <= 4'hce48;
         4'h6531 	:	val_out <= 4'hce48;
         4'h6532 	:	val_out <= 4'hce48;
         4'h6533 	:	val_out <= 4'hce48;
         4'h6538 	:	val_out <= 4'hce34;
         4'h6539 	:	val_out <= 4'hce34;
         4'h653a 	:	val_out <= 4'hce34;
         4'h653b 	:	val_out <= 4'hce34;
         4'h6540 	:	val_out <= 4'hce21;
         4'h6541 	:	val_out <= 4'hce21;
         4'h6542 	:	val_out <= 4'hce21;
         4'h6543 	:	val_out <= 4'hce21;
         4'h6548 	:	val_out <= 4'hce0d;
         4'h6549 	:	val_out <= 4'hce0d;
         4'h654a 	:	val_out <= 4'hce0d;
         4'h654b 	:	val_out <= 4'hce0d;
         4'h6550 	:	val_out <= 4'hcdf9;
         4'h6551 	:	val_out <= 4'hcdf9;
         4'h6552 	:	val_out <= 4'hcdf9;
         4'h6553 	:	val_out <= 4'hcdf9;
         4'h6558 	:	val_out <= 4'hcde5;
         4'h6559 	:	val_out <= 4'hcde5;
         4'h655a 	:	val_out <= 4'hcde5;
         4'h655b 	:	val_out <= 4'hcde5;
         4'h6560 	:	val_out <= 4'hcdd1;
         4'h6561 	:	val_out <= 4'hcdd1;
         4'h6562 	:	val_out <= 4'hcdd1;
         4'h6563 	:	val_out <= 4'hcdd1;
         4'h6568 	:	val_out <= 4'hcdbd;
         4'h6569 	:	val_out <= 4'hcdbd;
         4'h656a 	:	val_out <= 4'hcdbd;
         4'h656b 	:	val_out <= 4'hcdbd;
         4'h6570 	:	val_out <= 4'hcda9;
         4'h6571 	:	val_out <= 4'hcda9;
         4'h6572 	:	val_out <= 4'hcda9;
         4'h6573 	:	val_out <= 4'hcda9;
         4'h6578 	:	val_out <= 4'hcd95;
         4'h6579 	:	val_out <= 4'hcd95;
         4'h657a 	:	val_out <= 4'hcd95;
         4'h657b 	:	val_out <= 4'hcd95;
         4'h6580 	:	val_out <= 4'hcd81;
         4'h6581 	:	val_out <= 4'hcd81;
         4'h6582 	:	val_out <= 4'hcd81;
         4'h6583 	:	val_out <= 4'hcd81;
         4'h6588 	:	val_out <= 4'hcd6d;
         4'h6589 	:	val_out <= 4'hcd6d;
         4'h658a 	:	val_out <= 4'hcd6d;
         4'h658b 	:	val_out <= 4'hcd6d;
         4'h6590 	:	val_out <= 4'hcd59;
         4'h6591 	:	val_out <= 4'hcd59;
         4'h6592 	:	val_out <= 4'hcd59;
         4'h6593 	:	val_out <= 4'hcd59;
         4'h6598 	:	val_out <= 4'hcd45;
         4'h6599 	:	val_out <= 4'hcd45;
         4'h659a 	:	val_out <= 4'hcd45;
         4'h659b 	:	val_out <= 4'hcd45;
         4'h65a0 	:	val_out <= 4'hcd31;
         4'h65a1 	:	val_out <= 4'hcd31;
         4'h65a2 	:	val_out <= 4'hcd31;
         4'h65a3 	:	val_out <= 4'hcd31;
         4'h65a8 	:	val_out <= 4'hcd1d;
         4'h65a9 	:	val_out <= 4'hcd1d;
         4'h65aa 	:	val_out <= 4'hcd1d;
         4'h65ab 	:	val_out <= 4'hcd1d;
         4'h65b0 	:	val_out <= 4'hcd09;
         4'h65b1 	:	val_out <= 4'hcd09;
         4'h65b2 	:	val_out <= 4'hcd09;
         4'h65b3 	:	val_out <= 4'hcd09;
         4'h65b8 	:	val_out <= 4'hccf5;
         4'h65b9 	:	val_out <= 4'hccf5;
         4'h65ba 	:	val_out <= 4'hccf5;
         4'h65bb 	:	val_out <= 4'hccf5;
         4'h65c0 	:	val_out <= 4'hcce1;
         4'h65c1 	:	val_out <= 4'hcce1;
         4'h65c2 	:	val_out <= 4'hcce1;
         4'h65c3 	:	val_out <= 4'hcce1;
         4'h65c8 	:	val_out <= 4'hcccc;
         4'h65c9 	:	val_out <= 4'hcccc;
         4'h65ca 	:	val_out <= 4'hcccc;
         4'h65cb 	:	val_out <= 4'hcccc;
         4'h65d0 	:	val_out <= 4'hccb8;
         4'h65d1 	:	val_out <= 4'hccb8;
         4'h65d2 	:	val_out <= 4'hccb8;
         4'h65d3 	:	val_out <= 4'hccb8;
         4'h65d8 	:	val_out <= 4'hcca4;
         4'h65d9 	:	val_out <= 4'hcca4;
         4'h65da 	:	val_out <= 4'hcca4;
         4'h65db 	:	val_out <= 4'hcca4;
         4'h65e0 	:	val_out <= 4'hcc90;
         4'h65e1 	:	val_out <= 4'hcc90;
         4'h65e2 	:	val_out <= 4'hcc90;
         4'h65e3 	:	val_out <= 4'hcc90;
         4'h65e8 	:	val_out <= 4'hcc7c;
         4'h65e9 	:	val_out <= 4'hcc7c;
         4'h65ea 	:	val_out <= 4'hcc7c;
         4'h65eb 	:	val_out <= 4'hcc7c;
         4'h65f0 	:	val_out <= 4'hcc68;
         4'h65f1 	:	val_out <= 4'hcc68;
         4'h65f2 	:	val_out <= 4'hcc68;
         4'h65f3 	:	val_out <= 4'hcc68;
         4'h65f8 	:	val_out <= 4'hcc54;
         4'h65f9 	:	val_out <= 4'hcc54;
         4'h65fa 	:	val_out <= 4'hcc54;
         4'h65fb 	:	val_out <= 4'hcc54;
         4'h6600 	:	val_out <= 4'hcc3f;
         4'h6601 	:	val_out <= 4'hcc3f;
         4'h6602 	:	val_out <= 4'hcc3f;
         4'h6603 	:	val_out <= 4'hcc3f;
         4'h6608 	:	val_out <= 4'hcc2b;
         4'h6609 	:	val_out <= 4'hcc2b;
         4'h660a 	:	val_out <= 4'hcc2b;
         4'h660b 	:	val_out <= 4'hcc2b;
         4'h6610 	:	val_out <= 4'hcc17;
         4'h6611 	:	val_out <= 4'hcc17;
         4'h6612 	:	val_out <= 4'hcc17;
         4'h6613 	:	val_out <= 4'hcc17;
         4'h6618 	:	val_out <= 4'hcc03;
         4'h6619 	:	val_out <= 4'hcc03;
         4'h661a 	:	val_out <= 4'hcc03;
         4'h661b 	:	val_out <= 4'hcc03;
         4'h6620 	:	val_out <= 4'hcbef;
         4'h6621 	:	val_out <= 4'hcbef;
         4'h6622 	:	val_out <= 4'hcbef;
         4'h6623 	:	val_out <= 4'hcbef;
         4'h6628 	:	val_out <= 4'hcbda;
         4'h6629 	:	val_out <= 4'hcbda;
         4'h662a 	:	val_out <= 4'hcbda;
         4'h662b 	:	val_out <= 4'hcbda;
         4'h6630 	:	val_out <= 4'hcbc6;
         4'h6631 	:	val_out <= 4'hcbc6;
         4'h6632 	:	val_out <= 4'hcbc6;
         4'h6633 	:	val_out <= 4'hcbc6;
         4'h6638 	:	val_out <= 4'hcbb2;
         4'h6639 	:	val_out <= 4'hcbb2;
         4'h663a 	:	val_out <= 4'hcbb2;
         4'h663b 	:	val_out <= 4'hcbb2;
         4'h6640 	:	val_out <= 4'hcb9e;
         4'h6641 	:	val_out <= 4'hcb9e;
         4'h6642 	:	val_out <= 4'hcb9e;
         4'h6643 	:	val_out <= 4'hcb9e;
         4'h6648 	:	val_out <= 4'hcb89;
         4'h6649 	:	val_out <= 4'hcb89;
         4'h664a 	:	val_out <= 4'hcb89;
         4'h664b 	:	val_out <= 4'hcb89;
         4'h6650 	:	val_out <= 4'hcb75;
         4'h6651 	:	val_out <= 4'hcb75;
         4'h6652 	:	val_out <= 4'hcb75;
         4'h6653 	:	val_out <= 4'hcb75;
         4'h6658 	:	val_out <= 4'hcb61;
         4'h6659 	:	val_out <= 4'hcb61;
         4'h665a 	:	val_out <= 4'hcb61;
         4'h665b 	:	val_out <= 4'hcb61;
         4'h6660 	:	val_out <= 4'hcb4c;
         4'h6661 	:	val_out <= 4'hcb4c;
         4'h6662 	:	val_out <= 4'hcb4c;
         4'h6663 	:	val_out <= 4'hcb4c;
         4'h6668 	:	val_out <= 4'hcb38;
         4'h6669 	:	val_out <= 4'hcb38;
         4'h666a 	:	val_out <= 4'hcb38;
         4'h666b 	:	val_out <= 4'hcb38;
         4'h6670 	:	val_out <= 4'hcb24;
         4'h6671 	:	val_out <= 4'hcb24;
         4'h6672 	:	val_out <= 4'hcb24;
         4'h6673 	:	val_out <= 4'hcb24;
         4'h6678 	:	val_out <= 4'hcb0f;
         4'h6679 	:	val_out <= 4'hcb0f;
         4'h667a 	:	val_out <= 4'hcb0f;
         4'h667b 	:	val_out <= 4'hcb0f;
         4'h6680 	:	val_out <= 4'hcafb;
         4'h6681 	:	val_out <= 4'hcafb;
         4'h6682 	:	val_out <= 4'hcafb;
         4'h6683 	:	val_out <= 4'hcafb;
         4'h6688 	:	val_out <= 4'hcae7;
         4'h6689 	:	val_out <= 4'hcae7;
         4'h668a 	:	val_out <= 4'hcae7;
         4'h668b 	:	val_out <= 4'hcae7;
         4'h6690 	:	val_out <= 4'hcad2;
         4'h6691 	:	val_out <= 4'hcad2;
         4'h6692 	:	val_out <= 4'hcad2;
         4'h6693 	:	val_out <= 4'hcad2;
         4'h6698 	:	val_out <= 4'hcabe;
         4'h6699 	:	val_out <= 4'hcabe;
         4'h669a 	:	val_out <= 4'hcabe;
         4'h669b 	:	val_out <= 4'hcabe;
         4'h66a0 	:	val_out <= 4'hcaa9;
         4'h66a1 	:	val_out <= 4'hcaa9;
         4'h66a2 	:	val_out <= 4'hcaa9;
         4'h66a3 	:	val_out <= 4'hcaa9;
         4'h66a8 	:	val_out <= 4'hca95;
         4'h66a9 	:	val_out <= 4'hca95;
         4'h66aa 	:	val_out <= 4'hca95;
         4'h66ab 	:	val_out <= 4'hca95;
         4'h66b0 	:	val_out <= 4'hca81;
         4'h66b1 	:	val_out <= 4'hca81;
         4'h66b2 	:	val_out <= 4'hca81;
         4'h66b3 	:	val_out <= 4'hca81;
         4'h66b8 	:	val_out <= 4'hca6c;
         4'h66b9 	:	val_out <= 4'hca6c;
         4'h66ba 	:	val_out <= 4'hca6c;
         4'h66bb 	:	val_out <= 4'hca6c;
         4'h66c0 	:	val_out <= 4'hca58;
         4'h66c1 	:	val_out <= 4'hca58;
         4'h66c2 	:	val_out <= 4'hca58;
         4'h66c3 	:	val_out <= 4'hca58;
         4'h66c8 	:	val_out <= 4'hca43;
         4'h66c9 	:	val_out <= 4'hca43;
         4'h66ca 	:	val_out <= 4'hca43;
         4'h66cb 	:	val_out <= 4'hca43;
         4'h66d0 	:	val_out <= 4'hca2f;
         4'h66d1 	:	val_out <= 4'hca2f;
         4'h66d2 	:	val_out <= 4'hca2f;
         4'h66d3 	:	val_out <= 4'hca2f;
         4'h66d8 	:	val_out <= 4'hca1a;
         4'h66d9 	:	val_out <= 4'hca1a;
         4'h66da 	:	val_out <= 4'hca1a;
         4'h66db 	:	val_out <= 4'hca1a;
         4'h66e0 	:	val_out <= 4'hca06;
         4'h66e1 	:	val_out <= 4'hca06;
         4'h66e2 	:	val_out <= 4'hca06;
         4'h66e3 	:	val_out <= 4'hca06;
         4'h66e8 	:	val_out <= 4'hc9f1;
         4'h66e9 	:	val_out <= 4'hc9f1;
         4'h66ea 	:	val_out <= 4'hc9f1;
         4'h66eb 	:	val_out <= 4'hc9f1;
         4'h66f0 	:	val_out <= 4'hc9dd;
         4'h66f1 	:	val_out <= 4'hc9dd;
         4'h66f2 	:	val_out <= 4'hc9dd;
         4'h66f3 	:	val_out <= 4'hc9dd;
         4'h66f8 	:	val_out <= 4'hc9c8;
         4'h66f9 	:	val_out <= 4'hc9c8;
         4'h66fa 	:	val_out <= 4'hc9c8;
         4'h66fb 	:	val_out <= 4'hc9c8;
         4'h6700 	:	val_out <= 4'hc9b4;
         4'h6701 	:	val_out <= 4'hc9b4;
         4'h6702 	:	val_out <= 4'hc9b4;
         4'h6703 	:	val_out <= 4'hc9b4;
         4'h6708 	:	val_out <= 4'hc99f;
         4'h6709 	:	val_out <= 4'hc99f;
         4'h670a 	:	val_out <= 4'hc99f;
         4'h670b 	:	val_out <= 4'hc99f;
         4'h6710 	:	val_out <= 4'hc98a;
         4'h6711 	:	val_out <= 4'hc98a;
         4'h6712 	:	val_out <= 4'hc98a;
         4'h6713 	:	val_out <= 4'hc98a;
         4'h6718 	:	val_out <= 4'hc976;
         4'h6719 	:	val_out <= 4'hc976;
         4'h671a 	:	val_out <= 4'hc976;
         4'h671b 	:	val_out <= 4'hc976;
         4'h6720 	:	val_out <= 4'hc961;
         4'h6721 	:	val_out <= 4'hc961;
         4'h6722 	:	val_out <= 4'hc961;
         4'h6723 	:	val_out <= 4'hc961;
         4'h6728 	:	val_out <= 4'hc94d;
         4'h6729 	:	val_out <= 4'hc94d;
         4'h672a 	:	val_out <= 4'hc94d;
         4'h672b 	:	val_out <= 4'hc94d;
         4'h6730 	:	val_out <= 4'hc938;
         4'h6731 	:	val_out <= 4'hc938;
         4'h6732 	:	val_out <= 4'hc938;
         4'h6733 	:	val_out <= 4'hc938;
         4'h6738 	:	val_out <= 4'hc923;
         4'h6739 	:	val_out <= 4'hc923;
         4'h673a 	:	val_out <= 4'hc923;
         4'h673b 	:	val_out <= 4'hc923;
         4'h6740 	:	val_out <= 4'hc90f;
         4'h6741 	:	val_out <= 4'hc90f;
         4'h6742 	:	val_out <= 4'hc90f;
         4'h6743 	:	val_out <= 4'hc90f;
         4'h6748 	:	val_out <= 4'hc8fa;
         4'h6749 	:	val_out <= 4'hc8fa;
         4'h674a 	:	val_out <= 4'hc8fa;
         4'h674b 	:	val_out <= 4'hc8fa;
         4'h6750 	:	val_out <= 4'hc8e6;
         4'h6751 	:	val_out <= 4'hc8e6;
         4'h6752 	:	val_out <= 4'hc8e6;
         4'h6753 	:	val_out <= 4'hc8e6;
         4'h6758 	:	val_out <= 4'hc8d1;
         4'h6759 	:	val_out <= 4'hc8d1;
         4'h675a 	:	val_out <= 4'hc8d1;
         4'h675b 	:	val_out <= 4'hc8d1;
         4'h6760 	:	val_out <= 4'hc8bc;
         4'h6761 	:	val_out <= 4'hc8bc;
         4'h6762 	:	val_out <= 4'hc8bc;
         4'h6763 	:	val_out <= 4'hc8bc;
         4'h6768 	:	val_out <= 4'hc8a8;
         4'h6769 	:	val_out <= 4'hc8a8;
         4'h676a 	:	val_out <= 4'hc8a8;
         4'h676b 	:	val_out <= 4'hc8a8;
         4'h6770 	:	val_out <= 4'hc893;
         4'h6771 	:	val_out <= 4'hc893;
         4'h6772 	:	val_out <= 4'hc893;
         4'h6773 	:	val_out <= 4'hc893;
         4'h6778 	:	val_out <= 4'hc87e;
         4'h6779 	:	val_out <= 4'hc87e;
         4'h677a 	:	val_out <= 4'hc87e;
         4'h677b 	:	val_out <= 4'hc87e;
         4'h6780 	:	val_out <= 4'hc869;
         4'h6781 	:	val_out <= 4'hc869;
         4'h6782 	:	val_out <= 4'hc869;
         4'h6783 	:	val_out <= 4'hc869;
         4'h6788 	:	val_out <= 4'hc855;
         4'h6789 	:	val_out <= 4'hc855;
         4'h678a 	:	val_out <= 4'hc855;
         4'h678b 	:	val_out <= 4'hc855;
         4'h6790 	:	val_out <= 4'hc840;
         4'h6791 	:	val_out <= 4'hc840;
         4'h6792 	:	val_out <= 4'hc840;
         4'h6793 	:	val_out <= 4'hc840;
         4'h6798 	:	val_out <= 4'hc82b;
         4'h6799 	:	val_out <= 4'hc82b;
         4'h679a 	:	val_out <= 4'hc82b;
         4'h679b 	:	val_out <= 4'hc82b;
         4'h67a0 	:	val_out <= 4'hc816;
         4'h67a1 	:	val_out <= 4'hc816;
         4'h67a2 	:	val_out <= 4'hc816;
         4'h67a3 	:	val_out <= 4'hc816;
         4'h67a8 	:	val_out <= 4'hc802;
         4'h67a9 	:	val_out <= 4'hc802;
         4'h67aa 	:	val_out <= 4'hc802;
         4'h67ab 	:	val_out <= 4'hc802;
         4'h67b0 	:	val_out <= 4'hc7ed;
         4'h67b1 	:	val_out <= 4'hc7ed;
         4'h67b2 	:	val_out <= 4'hc7ed;
         4'h67b3 	:	val_out <= 4'hc7ed;
         4'h67b8 	:	val_out <= 4'hc7d8;
         4'h67b9 	:	val_out <= 4'hc7d8;
         4'h67ba 	:	val_out <= 4'hc7d8;
         4'h67bb 	:	val_out <= 4'hc7d8;
         4'h67c0 	:	val_out <= 4'hc7c3;
         4'h67c1 	:	val_out <= 4'hc7c3;
         4'h67c2 	:	val_out <= 4'hc7c3;
         4'h67c3 	:	val_out <= 4'hc7c3;
         4'h67c8 	:	val_out <= 4'hc7ae;
         4'h67c9 	:	val_out <= 4'hc7ae;
         4'h67ca 	:	val_out <= 4'hc7ae;
         4'h67cb 	:	val_out <= 4'hc7ae;
         4'h67d0 	:	val_out <= 4'hc79a;
         4'h67d1 	:	val_out <= 4'hc79a;
         4'h67d2 	:	val_out <= 4'hc79a;
         4'h67d3 	:	val_out <= 4'hc79a;
         4'h67d8 	:	val_out <= 4'hc785;
         4'h67d9 	:	val_out <= 4'hc785;
         4'h67da 	:	val_out <= 4'hc785;
         4'h67db 	:	val_out <= 4'hc785;
         4'h67e0 	:	val_out <= 4'hc770;
         4'h67e1 	:	val_out <= 4'hc770;
         4'h67e2 	:	val_out <= 4'hc770;
         4'h67e3 	:	val_out <= 4'hc770;
         4'h67e8 	:	val_out <= 4'hc75b;
         4'h67e9 	:	val_out <= 4'hc75b;
         4'h67ea 	:	val_out <= 4'hc75b;
         4'h67eb 	:	val_out <= 4'hc75b;
         4'h67f0 	:	val_out <= 4'hc746;
         4'h67f1 	:	val_out <= 4'hc746;
         4'h67f2 	:	val_out <= 4'hc746;
         4'h67f3 	:	val_out <= 4'hc746;
         4'h67f8 	:	val_out <= 4'hc731;
         4'h67f9 	:	val_out <= 4'hc731;
         4'h67fa 	:	val_out <= 4'hc731;
         4'h67fb 	:	val_out <= 4'hc731;
         4'h6800 	:	val_out <= 4'hc71c;
         4'h6801 	:	val_out <= 4'hc71c;
         4'h6802 	:	val_out <= 4'hc71c;
         4'h6803 	:	val_out <= 4'hc71c;
         4'h6808 	:	val_out <= 4'hc708;
         4'h6809 	:	val_out <= 4'hc708;
         4'h680a 	:	val_out <= 4'hc708;
         4'h680b 	:	val_out <= 4'hc708;
         4'h6810 	:	val_out <= 4'hc6f3;
         4'h6811 	:	val_out <= 4'hc6f3;
         4'h6812 	:	val_out <= 4'hc6f3;
         4'h6813 	:	val_out <= 4'hc6f3;
         4'h6818 	:	val_out <= 4'hc6de;
         4'h6819 	:	val_out <= 4'hc6de;
         4'h681a 	:	val_out <= 4'hc6de;
         4'h681b 	:	val_out <= 4'hc6de;
         4'h6820 	:	val_out <= 4'hc6c9;
         4'h6821 	:	val_out <= 4'hc6c9;
         4'h6822 	:	val_out <= 4'hc6c9;
         4'h6823 	:	val_out <= 4'hc6c9;
         4'h6828 	:	val_out <= 4'hc6b4;
         4'h6829 	:	val_out <= 4'hc6b4;
         4'h682a 	:	val_out <= 4'hc6b4;
         4'h682b 	:	val_out <= 4'hc6b4;
         4'h6830 	:	val_out <= 4'hc69f;
         4'h6831 	:	val_out <= 4'hc69f;
         4'h6832 	:	val_out <= 4'hc69f;
         4'h6833 	:	val_out <= 4'hc69f;
         4'h6838 	:	val_out <= 4'hc68a;
         4'h6839 	:	val_out <= 4'hc68a;
         4'h683a 	:	val_out <= 4'hc68a;
         4'h683b 	:	val_out <= 4'hc68a;
         4'h6840 	:	val_out <= 4'hc675;
         4'h6841 	:	val_out <= 4'hc675;
         4'h6842 	:	val_out <= 4'hc675;
         4'h6843 	:	val_out <= 4'hc675;
         4'h6848 	:	val_out <= 4'hc660;
         4'h6849 	:	val_out <= 4'hc660;
         4'h684a 	:	val_out <= 4'hc660;
         4'h684b 	:	val_out <= 4'hc660;
         4'h6850 	:	val_out <= 4'hc64b;
         4'h6851 	:	val_out <= 4'hc64b;
         4'h6852 	:	val_out <= 4'hc64b;
         4'h6853 	:	val_out <= 4'hc64b;
         4'h6858 	:	val_out <= 4'hc636;
         4'h6859 	:	val_out <= 4'hc636;
         4'h685a 	:	val_out <= 4'hc636;
         4'h685b 	:	val_out <= 4'hc636;
         4'h6860 	:	val_out <= 4'hc621;
         4'h6861 	:	val_out <= 4'hc621;
         4'h6862 	:	val_out <= 4'hc621;
         4'h6863 	:	val_out <= 4'hc621;
         4'h6868 	:	val_out <= 4'hc60c;
         4'h6869 	:	val_out <= 4'hc60c;
         4'h686a 	:	val_out <= 4'hc60c;
         4'h686b 	:	val_out <= 4'hc60c;
         4'h6870 	:	val_out <= 4'hc5f7;
         4'h6871 	:	val_out <= 4'hc5f7;
         4'h6872 	:	val_out <= 4'hc5f7;
         4'h6873 	:	val_out <= 4'hc5f7;
         4'h6878 	:	val_out <= 4'hc5e2;
         4'h6879 	:	val_out <= 4'hc5e2;
         4'h687a 	:	val_out <= 4'hc5e2;
         4'h687b 	:	val_out <= 4'hc5e2;
         4'h6880 	:	val_out <= 4'hc5cd;
         4'h6881 	:	val_out <= 4'hc5cd;
         4'h6882 	:	val_out <= 4'hc5cd;
         4'h6883 	:	val_out <= 4'hc5cd;
         4'h6888 	:	val_out <= 4'hc5b8;
         4'h6889 	:	val_out <= 4'hc5b8;
         4'h688a 	:	val_out <= 4'hc5b8;
         4'h688b 	:	val_out <= 4'hc5b8;
         4'h6890 	:	val_out <= 4'hc5a3;
         4'h6891 	:	val_out <= 4'hc5a3;
         4'h6892 	:	val_out <= 4'hc5a3;
         4'h6893 	:	val_out <= 4'hc5a3;
         4'h6898 	:	val_out <= 4'hc58d;
         4'h6899 	:	val_out <= 4'hc58d;
         4'h689a 	:	val_out <= 4'hc58d;
         4'h689b 	:	val_out <= 4'hc58d;
         4'h68a0 	:	val_out <= 4'hc578;
         4'h68a1 	:	val_out <= 4'hc578;
         4'h68a2 	:	val_out <= 4'hc578;
         4'h68a3 	:	val_out <= 4'hc578;
         4'h68a8 	:	val_out <= 4'hc563;
         4'h68a9 	:	val_out <= 4'hc563;
         4'h68aa 	:	val_out <= 4'hc563;
         4'h68ab 	:	val_out <= 4'hc563;
         4'h68b0 	:	val_out <= 4'hc54e;
         4'h68b1 	:	val_out <= 4'hc54e;
         4'h68b2 	:	val_out <= 4'hc54e;
         4'h68b3 	:	val_out <= 4'hc54e;
         4'h68b8 	:	val_out <= 4'hc539;
         4'h68b9 	:	val_out <= 4'hc539;
         4'h68ba 	:	val_out <= 4'hc539;
         4'h68bb 	:	val_out <= 4'hc539;
         4'h68c0 	:	val_out <= 4'hc524;
         4'h68c1 	:	val_out <= 4'hc524;
         4'h68c2 	:	val_out <= 4'hc524;
         4'h68c3 	:	val_out <= 4'hc524;
         4'h68c8 	:	val_out <= 4'hc50f;
         4'h68c9 	:	val_out <= 4'hc50f;
         4'h68ca 	:	val_out <= 4'hc50f;
         4'h68cb 	:	val_out <= 4'hc50f;
         4'h68d0 	:	val_out <= 4'hc4fa;
         4'h68d1 	:	val_out <= 4'hc4fa;
         4'h68d2 	:	val_out <= 4'hc4fa;
         4'h68d3 	:	val_out <= 4'hc4fa;
         4'h68d8 	:	val_out <= 4'hc4e4;
         4'h68d9 	:	val_out <= 4'hc4e4;
         4'h68da 	:	val_out <= 4'hc4e4;
         4'h68db 	:	val_out <= 4'hc4e4;
         4'h68e0 	:	val_out <= 4'hc4cf;
         4'h68e1 	:	val_out <= 4'hc4cf;
         4'h68e2 	:	val_out <= 4'hc4cf;
         4'h68e3 	:	val_out <= 4'hc4cf;
         4'h68e8 	:	val_out <= 4'hc4ba;
         4'h68e9 	:	val_out <= 4'hc4ba;
         4'h68ea 	:	val_out <= 4'hc4ba;
         4'h68eb 	:	val_out <= 4'hc4ba;
         4'h68f0 	:	val_out <= 4'hc4a5;
         4'h68f1 	:	val_out <= 4'hc4a5;
         4'h68f2 	:	val_out <= 4'hc4a5;
         4'h68f3 	:	val_out <= 4'hc4a5;
         4'h68f8 	:	val_out <= 4'hc490;
         4'h68f9 	:	val_out <= 4'hc490;
         4'h68fa 	:	val_out <= 4'hc490;
         4'h68fb 	:	val_out <= 4'hc490;
         4'h6900 	:	val_out <= 4'hc47a;
         4'h6901 	:	val_out <= 4'hc47a;
         4'h6902 	:	val_out <= 4'hc47a;
         4'h6903 	:	val_out <= 4'hc47a;
         4'h6908 	:	val_out <= 4'hc465;
         4'h6909 	:	val_out <= 4'hc465;
         4'h690a 	:	val_out <= 4'hc465;
         4'h690b 	:	val_out <= 4'hc465;
         4'h6910 	:	val_out <= 4'hc450;
         4'h6911 	:	val_out <= 4'hc450;
         4'h6912 	:	val_out <= 4'hc450;
         4'h6913 	:	val_out <= 4'hc450;
         4'h6918 	:	val_out <= 4'hc43b;
         4'h6919 	:	val_out <= 4'hc43b;
         4'h691a 	:	val_out <= 4'hc43b;
         4'h691b 	:	val_out <= 4'hc43b;
         4'h6920 	:	val_out <= 4'hc425;
         4'h6921 	:	val_out <= 4'hc425;
         4'h6922 	:	val_out <= 4'hc425;
         4'h6923 	:	val_out <= 4'hc425;
         4'h6928 	:	val_out <= 4'hc410;
         4'h6929 	:	val_out <= 4'hc410;
         4'h692a 	:	val_out <= 4'hc410;
         4'h692b 	:	val_out <= 4'hc410;
         4'h6930 	:	val_out <= 4'hc3fb;
         4'h6931 	:	val_out <= 4'hc3fb;
         4'h6932 	:	val_out <= 4'hc3fb;
         4'h6933 	:	val_out <= 4'hc3fb;
         4'h6938 	:	val_out <= 4'hc3e5;
         4'h6939 	:	val_out <= 4'hc3e5;
         4'h693a 	:	val_out <= 4'hc3e5;
         4'h693b 	:	val_out <= 4'hc3e5;
         4'h6940 	:	val_out <= 4'hc3d0;
         4'h6941 	:	val_out <= 4'hc3d0;
         4'h6942 	:	val_out <= 4'hc3d0;
         4'h6943 	:	val_out <= 4'hc3d0;
         4'h6948 	:	val_out <= 4'hc3bb;
         4'h6949 	:	val_out <= 4'hc3bb;
         4'h694a 	:	val_out <= 4'hc3bb;
         4'h694b 	:	val_out <= 4'hc3bb;
         4'h6950 	:	val_out <= 4'hc3a5;
         4'h6951 	:	val_out <= 4'hc3a5;
         4'h6952 	:	val_out <= 4'hc3a5;
         4'h6953 	:	val_out <= 4'hc3a5;
         4'h6958 	:	val_out <= 4'hc390;
         4'h6959 	:	val_out <= 4'hc390;
         4'h695a 	:	val_out <= 4'hc390;
         4'h695b 	:	val_out <= 4'hc390;
         4'h6960 	:	val_out <= 4'hc37b;
         4'h6961 	:	val_out <= 4'hc37b;
         4'h6962 	:	val_out <= 4'hc37b;
         4'h6963 	:	val_out <= 4'hc37b;
         4'h6968 	:	val_out <= 4'hc365;
         4'h6969 	:	val_out <= 4'hc365;
         4'h696a 	:	val_out <= 4'hc365;
         4'h696b 	:	val_out <= 4'hc365;
         4'h6970 	:	val_out <= 4'hc350;
         4'h6971 	:	val_out <= 4'hc350;
         4'h6972 	:	val_out <= 4'hc350;
         4'h6973 	:	val_out <= 4'hc350;
         4'h6978 	:	val_out <= 4'hc33b;
         4'h6979 	:	val_out <= 4'hc33b;
         4'h697a 	:	val_out <= 4'hc33b;
         4'h697b 	:	val_out <= 4'hc33b;
         4'h6980 	:	val_out <= 4'hc325;
         4'h6981 	:	val_out <= 4'hc325;
         4'h6982 	:	val_out <= 4'hc325;
         4'h6983 	:	val_out <= 4'hc325;
         4'h6988 	:	val_out <= 4'hc310;
         4'h6989 	:	val_out <= 4'hc310;
         4'h698a 	:	val_out <= 4'hc310;
         4'h698b 	:	val_out <= 4'hc310;
         4'h6990 	:	val_out <= 4'hc2fa;
         4'h6991 	:	val_out <= 4'hc2fa;
         4'h6992 	:	val_out <= 4'hc2fa;
         4'h6993 	:	val_out <= 4'hc2fa;
         4'h6998 	:	val_out <= 4'hc2e5;
         4'h6999 	:	val_out <= 4'hc2e5;
         4'h699a 	:	val_out <= 4'hc2e5;
         4'h699b 	:	val_out <= 4'hc2e5;
         4'h69a0 	:	val_out <= 4'hc2d0;
         4'h69a1 	:	val_out <= 4'hc2d0;
         4'h69a2 	:	val_out <= 4'hc2d0;
         4'h69a3 	:	val_out <= 4'hc2d0;
         4'h69a8 	:	val_out <= 4'hc2ba;
         4'h69a9 	:	val_out <= 4'hc2ba;
         4'h69aa 	:	val_out <= 4'hc2ba;
         4'h69ab 	:	val_out <= 4'hc2ba;
         4'h69b0 	:	val_out <= 4'hc2a5;
         4'h69b1 	:	val_out <= 4'hc2a5;
         4'h69b2 	:	val_out <= 4'hc2a5;
         4'h69b3 	:	val_out <= 4'hc2a5;
         4'h69b8 	:	val_out <= 4'hc28f;
         4'h69b9 	:	val_out <= 4'hc28f;
         4'h69ba 	:	val_out <= 4'hc28f;
         4'h69bb 	:	val_out <= 4'hc28f;
         4'h69c0 	:	val_out <= 4'hc27a;
         4'h69c1 	:	val_out <= 4'hc27a;
         4'h69c2 	:	val_out <= 4'hc27a;
         4'h69c3 	:	val_out <= 4'hc27a;
         4'h69c8 	:	val_out <= 4'hc264;
         4'h69c9 	:	val_out <= 4'hc264;
         4'h69ca 	:	val_out <= 4'hc264;
         4'h69cb 	:	val_out <= 4'hc264;
         4'h69d0 	:	val_out <= 4'hc24f;
         4'h69d1 	:	val_out <= 4'hc24f;
         4'h69d2 	:	val_out <= 4'hc24f;
         4'h69d3 	:	val_out <= 4'hc24f;
         4'h69d8 	:	val_out <= 4'hc239;
         4'h69d9 	:	val_out <= 4'hc239;
         4'h69da 	:	val_out <= 4'hc239;
         4'h69db 	:	val_out <= 4'hc239;
         4'h69e0 	:	val_out <= 4'hc224;
         4'h69e1 	:	val_out <= 4'hc224;
         4'h69e2 	:	val_out <= 4'hc224;
         4'h69e3 	:	val_out <= 4'hc224;
         4'h69e8 	:	val_out <= 4'hc20e;
         4'h69e9 	:	val_out <= 4'hc20e;
         4'h69ea 	:	val_out <= 4'hc20e;
         4'h69eb 	:	val_out <= 4'hc20e;
         4'h69f0 	:	val_out <= 4'hc1f9;
         4'h69f1 	:	val_out <= 4'hc1f9;
         4'h69f2 	:	val_out <= 4'hc1f9;
         4'h69f3 	:	val_out <= 4'hc1f9;
         4'h69f8 	:	val_out <= 4'hc1e3;
         4'h69f9 	:	val_out <= 4'hc1e3;
         4'h69fa 	:	val_out <= 4'hc1e3;
         4'h69fb 	:	val_out <= 4'hc1e3;
         4'h6a00 	:	val_out <= 4'hc1ce;
         4'h6a01 	:	val_out <= 4'hc1ce;
         4'h6a02 	:	val_out <= 4'hc1ce;
         4'h6a03 	:	val_out <= 4'hc1ce;
         4'h6a08 	:	val_out <= 4'hc1b8;
         4'h6a09 	:	val_out <= 4'hc1b8;
         4'h6a0a 	:	val_out <= 4'hc1b8;
         4'h6a0b 	:	val_out <= 4'hc1b8;
         4'h6a10 	:	val_out <= 4'hc1a2;
         4'h6a11 	:	val_out <= 4'hc1a2;
         4'h6a12 	:	val_out <= 4'hc1a2;
         4'h6a13 	:	val_out <= 4'hc1a2;
         4'h6a18 	:	val_out <= 4'hc18d;
         4'h6a19 	:	val_out <= 4'hc18d;
         4'h6a1a 	:	val_out <= 4'hc18d;
         4'h6a1b 	:	val_out <= 4'hc18d;
         4'h6a20 	:	val_out <= 4'hc177;
         4'h6a21 	:	val_out <= 4'hc177;
         4'h6a22 	:	val_out <= 4'hc177;
         4'h6a23 	:	val_out <= 4'hc177;
         4'h6a28 	:	val_out <= 4'hc162;
         4'h6a29 	:	val_out <= 4'hc162;
         4'h6a2a 	:	val_out <= 4'hc162;
         4'h6a2b 	:	val_out <= 4'hc162;
         4'h6a30 	:	val_out <= 4'hc14c;
         4'h6a31 	:	val_out <= 4'hc14c;
         4'h6a32 	:	val_out <= 4'hc14c;
         4'h6a33 	:	val_out <= 4'hc14c;
         4'h6a38 	:	val_out <= 4'hc136;
         4'h6a39 	:	val_out <= 4'hc136;
         4'h6a3a 	:	val_out <= 4'hc136;
         4'h6a3b 	:	val_out <= 4'hc136;
         4'h6a40 	:	val_out <= 4'hc121;
         4'h6a41 	:	val_out <= 4'hc121;
         4'h6a42 	:	val_out <= 4'hc121;
         4'h6a43 	:	val_out <= 4'hc121;
         4'h6a48 	:	val_out <= 4'hc10b;
         4'h6a49 	:	val_out <= 4'hc10b;
         4'h6a4a 	:	val_out <= 4'hc10b;
         4'h6a4b 	:	val_out <= 4'hc10b;
         4'h6a50 	:	val_out <= 4'hc0f6;
         4'h6a51 	:	val_out <= 4'hc0f6;
         4'h6a52 	:	val_out <= 4'hc0f6;
         4'h6a53 	:	val_out <= 4'hc0f6;
         4'h6a58 	:	val_out <= 4'hc0e0;
         4'h6a59 	:	val_out <= 4'hc0e0;
         4'h6a5a 	:	val_out <= 4'hc0e0;
         4'h6a5b 	:	val_out <= 4'hc0e0;
         4'h6a60 	:	val_out <= 4'hc0ca;
         4'h6a61 	:	val_out <= 4'hc0ca;
         4'h6a62 	:	val_out <= 4'hc0ca;
         4'h6a63 	:	val_out <= 4'hc0ca;
         4'h6a68 	:	val_out <= 4'hc0b5;
         4'h6a69 	:	val_out <= 4'hc0b5;
         4'h6a6a 	:	val_out <= 4'hc0b5;
         4'h6a6b 	:	val_out <= 4'hc0b5;
         4'h6a70 	:	val_out <= 4'hc09f;
         4'h6a71 	:	val_out <= 4'hc09f;
         4'h6a72 	:	val_out <= 4'hc09f;
         4'h6a73 	:	val_out <= 4'hc09f;
         4'h6a78 	:	val_out <= 4'hc089;
         4'h6a79 	:	val_out <= 4'hc089;
         4'h6a7a 	:	val_out <= 4'hc089;
         4'h6a7b 	:	val_out <= 4'hc089;
         4'h6a80 	:	val_out <= 4'hc073;
         4'h6a81 	:	val_out <= 4'hc073;
         4'h6a82 	:	val_out <= 4'hc073;
         4'h6a83 	:	val_out <= 4'hc073;
         4'h6a88 	:	val_out <= 4'hc05e;
         4'h6a89 	:	val_out <= 4'hc05e;
         4'h6a8a 	:	val_out <= 4'hc05e;
         4'h6a8b 	:	val_out <= 4'hc05e;
         4'h6a90 	:	val_out <= 4'hc048;
         4'h6a91 	:	val_out <= 4'hc048;
         4'h6a92 	:	val_out <= 4'hc048;
         4'h6a93 	:	val_out <= 4'hc048;
         4'h6a98 	:	val_out <= 4'hc032;
         4'h6a99 	:	val_out <= 4'hc032;
         4'h6a9a 	:	val_out <= 4'hc032;
         4'h6a9b 	:	val_out <= 4'hc032;
         4'h6aa0 	:	val_out <= 4'hc01d;
         4'h6aa1 	:	val_out <= 4'hc01d;
         4'h6aa2 	:	val_out <= 4'hc01d;
         4'h6aa3 	:	val_out <= 4'hc01d;
         4'h6aa8 	:	val_out <= 4'hc007;
         4'h6aa9 	:	val_out <= 4'hc007;
         4'h6aaa 	:	val_out <= 4'hc007;
         4'h6aab 	:	val_out <= 4'hc007;
         4'h6ab0 	:	val_out <= 4'hbff1;
         4'h6ab1 	:	val_out <= 4'hbff1;
         4'h6ab2 	:	val_out <= 4'hbff1;
         4'h6ab3 	:	val_out <= 4'hbff1;
         4'h6ab8 	:	val_out <= 4'hbfdb;
         4'h6ab9 	:	val_out <= 4'hbfdb;
         4'h6aba 	:	val_out <= 4'hbfdb;
         4'h6abb 	:	val_out <= 4'hbfdb;
         4'h6ac0 	:	val_out <= 4'hbfc5;
         4'h6ac1 	:	val_out <= 4'hbfc5;
         4'h6ac2 	:	val_out <= 4'hbfc5;
         4'h6ac3 	:	val_out <= 4'hbfc5;
         4'h6ac8 	:	val_out <= 4'hbfb0;
         4'h6ac9 	:	val_out <= 4'hbfb0;
         4'h6aca 	:	val_out <= 4'hbfb0;
         4'h6acb 	:	val_out <= 4'hbfb0;
         4'h6ad0 	:	val_out <= 4'hbf9a;
         4'h6ad1 	:	val_out <= 4'hbf9a;
         4'h6ad2 	:	val_out <= 4'hbf9a;
         4'h6ad3 	:	val_out <= 4'hbf9a;
         4'h6ad8 	:	val_out <= 4'hbf84;
         4'h6ad9 	:	val_out <= 4'hbf84;
         4'h6ada 	:	val_out <= 4'hbf84;
         4'h6adb 	:	val_out <= 4'hbf84;
         4'h6ae0 	:	val_out <= 4'hbf6e;
         4'h6ae1 	:	val_out <= 4'hbf6e;
         4'h6ae2 	:	val_out <= 4'hbf6e;
         4'h6ae3 	:	val_out <= 4'hbf6e;
         4'h6ae8 	:	val_out <= 4'hbf58;
         4'h6ae9 	:	val_out <= 4'hbf58;
         4'h6aea 	:	val_out <= 4'hbf58;
         4'h6aeb 	:	val_out <= 4'hbf58;
         4'h6af0 	:	val_out <= 4'hbf43;
         4'h6af1 	:	val_out <= 4'hbf43;
         4'h6af2 	:	val_out <= 4'hbf43;
         4'h6af3 	:	val_out <= 4'hbf43;
         4'h6af8 	:	val_out <= 4'hbf2d;
         4'h6af9 	:	val_out <= 4'hbf2d;
         4'h6afa 	:	val_out <= 4'hbf2d;
         4'h6afb 	:	val_out <= 4'hbf2d;
         4'h6b00 	:	val_out <= 4'hbf17;
         4'h6b01 	:	val_out <= 4'hbf17;
         4'h6b02 	:	val_out <= 4'hbf17;
         4'h6b03 	:	val_out <= 4'hbf17;
         4'h6b08 	:	val_out <= 4'hbf01;
         4'h6b09 	:	val_out <= 4'hbf01;
         4'h6b0a 	:	val_out <= 4'hbf01;
         4'h6b0b 	:	val_out <= 4'hbf01;
         4'h6b10 	:	val_out <= 4'hbeeb;
         4'h6b11 	:	val_out <= 4'hbeeb;
         4'h6b12 	:	val_out <= 4'hbeeb;
         4'h6b13 	:	val_out <= 4'hbeeb;
         4'h6b18 	:	val_out <= 4'hbed5;
         4'h6b19 	:	val_out <= 4'hbed5;
         4'h6b1a 	:	val_out <= 4'hbed5;
         4'h6b1b 	:	val_out <= 4'hbed5;
         4'h6b20 	:	val_out <= 4'hbebf;
         4'h6b21 	:	val_out <= 4'hbebf;
         4'h6b22 	:	val_out <= 4'hbebf;
         4'h6b23 	:	val_out <= 4'hbebf;
         4'h6b28 	:	val_out <= 4'hbea9;
         4'h6b29 	:	val_out <= 4'hbea9;
         4'h6b2a 	:	val_out <= 4'hbea9;
         4'h6b2b 	:	val_out <= 4'hbea9;
         4'h6b30 	:	val_out <= 4'hbe93;
         4'h6b31 	:	val_out <= 4'hbe93;
         4'h6b32 	:	val_out <= 4'hbe93;
         4'h6b33 	:	val_out <= 4'hbe93;
         4'h6b38 	:	val_out <= 4'hbe7d;
         4'h6b39 	:	val_out <= 4'hbe7d;
         4'h6b3a 	:	val_out <= 4'hbe7d;
         4'h6b3b 	:	val_out <= 4'hbe7d;
         4'h6b40 	:	val_out <= 4'hbe68;
         4'h6b41 	:	val_out <= 4'hbe68;
         4'h6b42 	:	val_out <= 4'hbe68;
         4'h6b43 	:	val_out <= 4'hbe68;
         4'h6b48 	:	val_out <= 4'hbe52;
         4'h6b49 	:	val_out <= 4'hbe52;
         4'h6b4a 	:	val_out <= 4'hbe52;
         4'h6b4b 	:	val_out <= 4'hbe52;
         4'h6b50 	:	val_out <= 4'hbe3c;
         4'h6b51 	:	val_out <= 4'hbe3c;
         4'h6b52 	:	val_out <= 4'hbe3c;
         4'h6b53 	:	val_out <= 4'hbe3c;
         4'h6b58 	:	val_out <= 4'hbe26;
         4'h6b59 	:	val_out <= 4'hbe26;
         4'h6b5a 	:	val_out <= 4'hbe26;
         4'h6b5b 	:	val_out <= 4'hbe26;
         4'h6b60 	:	val_out <= 4'hbe10;
         4'h6b61 	:	val_out <= 4'hbe10;
         4'h6b62 	:	val_out <= 4'hbe10;
         4'h6b63 	:	val_out <= 4'hbe10;
         4'h6b68 	:	val_out <= 4'hbdfa;
         4'h6b69 	:	val_out <= 4'hbdfa;
         4'h6b6a 	:	val_out <= 4'hbdfa;
         4'h6b6b 	:	val_out <= 4'hbdfa;
         4'h6b70 	:	val_out <= 4'hbde4;
         4'h6b71 	:	val_out <= 4'hbde4;
         4'h6b72 	:	val_out <= 4'hbde4;
         4'h6b73 	:	val_out <= 4'hbde4;
         4'h6b78 	:	val_out <= 4'hbdce;
         4'h6b79 	:	val_out <= 4'hbdce;
         4'h6b7a 	:	val_out <= 4'hbdce;
         4'h6b7b 	:	val_out <= 4'hbdce;
         4'h6b80 	:	val_out <= 4'hbdb8;
         4'h6b81 	:	val_out <= 4'hbdb8;
         4'h6b82 	:	val_out <= 4'hbdb8;
         4'h6b83 	:	val_out <= 4'hbdb8;
         4'h6b88 	:	val_out <= 4'hbda2;
         4'h6b89 	:	val_out <= 4'hbda2;
         4'h6b8a 	:	val_out <= 4'hbda2;
         4'h6b8b 	:	val_out <= 4'hbda2;
         4'h6b90 	:	val_out <= 4'hbd8c;
         4'h6b91 	:	val_out <= 4'hbd8c;
         4'h6b92 	:	val_out <= 4'hbd8c;
         4'h6b93 	:	val_out <= 4'hbd8c;
         4'h6b98 	:	val_out <= 4'hbd76;
         4'h6b99 	:	val_out <= 4'hbd76;
         4'h6b9a 	:	val_out <= 4'hbd76;
         4'h6b9b 	:	val_out <= 4'hbd76;
         4'h6ba0 	:	val_out <= 4'hbd60;
         4'h6ba1 	:	val_out <= 4'hbd60;
         4'h6ba2 	:	val_out <= 4'hbd60;
         4'h6ba3 	:	val_out <= 4'hbd60;
         4'h6ba8 	:	val_out <= 4'hbd49;
         4'h6ba9 	:	val_out <= 4'hbd49;
         4'h6baa 	:	val_out <= 4'hbd49;
         4'h6bab 	:	val_out <= 4'hbd49;
         4'h6bb0 	:	val_out <= 4'hbd33;
         4'h6bb1 	:	val_out <= 4'hbd33;
         4'h6bb2 	:	val_out <= 4'hbd33;
         4'h6bb3 	:	val_out <= 4'hbd33;
         4'h6bb8 	:	val_out <= 4'hbd1d;
         4'h6bb9 	:	val_out <= 4'hbd1d;
         4'h6bba 	:	val_out <= 4'hbd1d;
         4'h6bbb 	:	val_out <= 4'hbd1d;
         4'h6bc0 	:	val_out <= 4'hbd07;
         4'h6bc1 	:	val_out <= 4'hbd07;
         4'h6bc2 	:	val_out <= 4'hbd07;
         4'h6bc3 	:	val_out <= 4'hbd07;
         4'h6bc8 	:	val_out <= 4'hbcf1;
         4'h6bc9 	:	val_out <= 4'hbcf1;
         4'h6bca 	:	val_out <= 4'hbcf1;
         4'h6bcb 	:	val_out <= 4'hbcf1;
         4'h6bd0 	:	val_out <= 4'hbcdb;
         4'h6bd1 	:	val_out <= 4'hbcdb;
         4'h6bd2 	:	val_out <= 4'hbcdb;
         4'h6bd3 	:	val_out <= 4'hbcdb;
         4'h6bd8 	:	val_out <= 4'hbcc5;
         4'h6bd9 	:	val_out <= 4'hbcc5;
         4'h6bda 	:	val_out <= 4'hbcc5;
         4'h6bdb 	:	val_out <= 4'hbcc5;
         4'h6be0 	:	val_out <= 4'hbcaf;
         4'h6be1 	:	val_out <= 4'hbcaf;
         4'h6be2 	:	val_out <= 4'hbcaf;
         4'h6be3 	:	val_out <= 4'hbcaf;
         4'h6be8 	:	val_out <= 4'hbc99;
         4'h6be9 	:	val_out <= 4'hbc99;
         4'h6bea 	:	val_out <= 4'hbc99;
         4'h6beb 	:	val_out <= 4'hbc99;
         4'h6bf0 	:	val_out <= 4'hbc83;
         4'h6bf1 	:	val_out <= 4'hbc83;
         4'h6bf2 	:	val_out <= 4'hbc83;
         4'h6bf3 	:	val_out <= 4'hbc83;
         4'h6bf8 	:	val_out <= 4'hbc6c;
         4'h6bf9 	:	val_out <= 4'hbc6c;
         4'h6bfa 	:	val_out <= 4'hbc6c;
         4'h6bfb 	:	val_out <= 4'hbc6c;
         4'h6c00 	:	val_out <= 4'hbc56;
         4'h6c01 	:	val_out <= 4'hbc56;
         4'h6c02 	:	val_out <= 4'hbc56;
         4'h6c03 	:	val_out <= 4'hbc56;
         4'h6c08 	:	val_out <= 4'hbc40;
         4'h6c09 	:	val_out <= 4'hbc40;
         4'h6c0a 	:	val_out <= 4'hbc40;
         4'h6c0b 	:	val_out <= 4'hbc40;
         4'h6c10 	:	val_out <= 4'hbc2a;
         4'h6c11 	:	val_out <= 4'hbc2a;
         4'h6c12 	:	val_out <= 4'hbc2a;
         4'h6c13 	:	val_out <= 4'hbc2a;
         4'h6c18 	:	val_out <= 4'hbc14;
         4'h6c19 	:	val_out <= 4'hbc14;
         4'h6c1a 	:	val_out <= 4'hbc14;
         4'h6c1b 	:	val_out <= 4'hbc14;
         4'h6c20 	:	val_out <= 4'hbbfd;
         4'h6c21 	:	val_out <= 4'hbbfd;
         4'h6c22 	:	val_out <= 4'hbbfd;
         4'h6c23 	:	val_out <= 4'hbbfd;
         4'h6c28 	:	val_out <= 4'hbbe7;
         4'h6c29 	:	val_out <= 4'hbbe7;
         4'h6c2a 	:	val_out <= 4'hbbe7;
         4'h6c2b 	:	val_out <= 4'hbbe7;
         4'h6c30 	:	val_out <= 4'hbbd1;
         4'h6c31 	:	val_out <= 4'hbbd1;
         4'h6c32 	:	val_out <= 4'hbbd1;
         4'h6c33 	:	val_out <= 4'hbbd1;
         4'h6c38 	:	val_out <= 4'hbbbb;
         4'h6c39 	:	val_out <= 4'hbbbb;
         4'h6c3a 	:	val_out <= 4'hbbbb;
         4'h6c3b 	:	val_out <= 4'hbbbb;
         4'h6c40 	:	val_out <= 4'hbba5;
         4'h6c41 	:	val_out <= 4'hbba5;
         4'h6c42 	:	val_out <= 4'hbba5;
         4'h6c43 	:	val_out <= 4'hbba5;
         4'h6c48 	:	val_out <= 4'hbb8e;
         4'h6c49 	:	val_out <= 4'hbb8e;
         4'h6c4a 	:	val_out <= 4'hbb8e;
         4'h6c4b 	:	val_out <= 4'hbb8e;
         4'h6c50 	:	val_out <= 4'hbb78;
         4'h6c51 	:	val_out <= 4'hbb78;
         4'h6c52 	:	val_out <= 4'hbb78;
         4'h6c53 	:	val_out <= 4'hbb78;
         4'h6c58 	:	val_out <= 4'hbb62;
         4'h6c59 	:	val_out <= 4'hbb62;
         4'h6c5a 	:	val_out <= 4'hbb62;
         4'h6c5b 	:	val_out <= 4'hbb62;
         4'h6c60 	:	val_out <= 4'hbb4c;
         4'h6c61 	:	val_out <= 4'hbb4c;
         4'h6c62 	:	val_out <= 4'hbb4c;
         4'h6c63 	:	val_out <= 4'hbb4c;
         4'h6c68 	:	val_out <= 4'hbb35;
         4'h6c69 	:	val_out <= 4'hbb35;
         4'h6c6a 	:	val_out <= 4'hbb35;
         4'h6c6b 	:	val_out <= 4'hbb35;
         4'h6c70 	:	val_out <= 4'hbb1f;
         4'h6c71 	:	val_out <= 4'hbb1f;
         4'h6c72 	:	val_out <= 4'hbb1f;
         4'h6c73 	:	val_out <= 4'hbb1f;
         4'h6c78 	:	val_out <= 4'hbb09;
         4'h6c79 	:	val_out <= 4'hbb09;
         4'h6c7a 	:	val_out <= 4'hbb09;
         4'h6c7b 	:	val_out <= 4'hbb09;
         4'h6c80 	:	val_out <= 4'hbaf2;
         4'h6c81 	:	val_out <= 4'hbaf2;
         4'h6c82 	:	val_out <= 4'hbaf2;
         4'h6c83 	:	val_out <= 4'hbaf2;
         4'h6c88 	:	val_out <= 4'hbadc;
         4'h6c89 	:	val_out <= 4'hbadc;
         4'h6c8a 	:	val_out <= 4'hbadc;
         4'h6c8b 	:	val_out <= 4'hbadc;
         4'h6c90 	:	val_out <= 4'hbac6;
         4'h6c91 	:	val_out <= 4'hbac6;
         4'h6c92 	:	val_out <= 4'hbac6;
         4'h6c93 	:	val_out <= 4'hbac6;
         4'h6c98 	:	val_out <= 4'hbaaf;
         4'h6c99 	:	val_out <= 4'hbaaf;
         4'h6c9a 	:	val_out <= 4'hbaaf;
         4'h6c9b 	:	val_out <= 4'hbaaf;
         4'h6ca0 	:	val_out <= 4'hba99;
         4'h6ca1 	:	val_out <= 4'hba99;
         4'h6ca2 	:	val_out <= 4'hba99;
         4'h6ca3 	:	val_out <= 4'hba99;
         4'h6ca8 	:	val_out <= 4'hba83;
         4'h6ca9 	:	val_out <= 4'hba83;
         4'h6caa 	:	val_out <= 4'hba83;
         4'h6cab 	:	val_out <= 4'hba83;
         4'h6cb0 	:	val_out <= 4'hba6c;
         4'h6cb1 	:	val_out <= 4'hba6c;
         4'h6cb2 	:	val_out <= 4'hba6c;
         4'h6cb3 	:	val_out <= 4'hba6c;
         4'h6cb8 	:	val_out <= 4'hba56;
         4'h6cb9 	:	val_out <= 4'hba56;
         4'h6cba 	:	val_out <= 4'hba56;
         4'h6cbb 	:	val_out <= 4'hba56;
         4'h6cc0 	:	val_out <= 4'hba40;
         4'h6cc1 	:	val_out <= 4'hba40;
         4'h6cc2 	:	val_out <= 4'hba40;
         4'h6cc3 	:	val_out <= 4'hba40;
         4'h6cc8 	:	val_out <= 4'hba29;
         4'h6cc9 	:	val_out <= 4'hba29;
         4'h6cca 	:	val_out <= 4'hba29;
         4'h6ccb 	:	val_out <= 4'hba29;
         4'h6cd0 	:	val_out <= 4'hba13;
         4'h6cd1 	:	val_out <= 4'hba13;
         4'h6cd2 	:	val_out <= 4'hba13;
         4'h6cd3 	:	val_out <= 4'hba13;
         4'h6cd8 	:	val_out <= 4'hb9fd;
         4'h6cd9 	:	val_out <= 4'hb9fd;
         4'h6cda 	:	val_out <= 4'hb9fd;
         4'h6cdb 	:	val_out <= 4'hb9fd;
         4'h6ce0 	:	val_out <= 4'hb9e6;
         4'h6ce1 	:	val_out <= 4'hb9e6;
         4'h6ce2 	:	val_out <= 4'hb9e6;
         4'h6ce3 	:	val_out <= 4'hb9e6;
         4'h6ce8 	:	val_out <= 4'hb9d0;
         4'h6ce9 	:	val_out <= 4'hb9d0;
         4'h6cea 	:	val_out <= 4'hb9d0;
         4'h6ceb 	:	val_out <= 4'hb9d0;
         4'h6cf0 	:	val_out <= 4'hb9b9;
         4'h6cf1 	:	val_out <= 4'hb9b9;
         4'h6cf2 	:	val_out <= 4'hb9b9;
         4'h6cf3 	:	val_out <= 4'hb9b9;
         4'h6cf8 	:	val_out <= 4'hb9a3;
         4'h6cf9 	:	val_out <= 4'hb9a3;
         4'h6cfa 	:	val_out <= 4'hb9a3;
         4'h6cfb 	:	val_out <= 4'hb9a3;
         4'h6d00 	:	val_out <= 4'hb98c;
         4'h6d01 	:	val_out <= 4'hb98c;
         4'h6d02 	:	val_out <= 4'hb98c;
         4'h6d03 	:	val_out <= 4'hb98c;
         4'h6d08 	:	val_out <= 4'hb976;
         4'h6d09 	:	val_out <= 4'hb976;
         4'h6d0a 	:	val_out <= 4'hb976;
         4'h6d0b 	:	val_out <= 4'hb976;
         4'h6d10 	:	val_out <= 4'hb95f;
         4'h6d11 	:	val_out <= 4'hb95f;
         4'h6d12 	:	val_out <= 4'hb95f;
         4'h6d13 	:	val_out <= 4'hb95f;
         4'h6d18 	:	val_out <= 4'hb949;
         4'h6d19 	:	val_out <= 4'hb949;
         4'h6d1a 	:	val_out <= 4'hb949;
         4'h6d1b 	:	val_out <= 4'hb949;
         4'h6d20 	:	val_out <= 4'hb932;
         4'h6d21 	:	val_out <= 4'hb932;
         4'h6d22 	:	val_out <= 4'hb932;
         4'h6d23 	:	val_out <= 4'hb932;
         4'h6d28 	:	val_out <= 4'hb91c;
         4'h6d29 	:	val_out <= 4'hb91c;
         4'h6d2a 	:	val_out <= 4'hb91c;
         4'h6d2b 	:	val_out <= 4'hb91c;
         4'h6d30 	:	val_out <= 4'hb906;
         4'h6d31 	:	val_out <= 4'hb906;
         4'h6d32 	:	val_out <= 4'hb906;
         4'h6d33 	:	val_out <= 4'hb906;
         4'h6d38 	:	val_out <= 4'hb8ef;
         4'h6d39 	:	val_out <= 4'hb8ef;
         4'h6d3a 	:	val_out <= 4'hb8ef;
         4'h6d3b 	:	val_out <= 4'hb8ef;
         4'h6d40 	:	val_out <= 4'hb8d8;
         4'h6d41 	:	val_out <= 4'hb8d8;
         4'h6d42 	:	val_out <= 4'hb8d8;
         4'h6d43 	:	val_out <= 4'hb8d8;
         4'h6d48 	:	val_out <= 4'hb8c2;
         4'h6d49 	:	val_out <= 4'hb8c2;
         4'h6d4a 	:	val_out <= 4'hb8c2;
         4'h6d4b 	:	val_out <= 4'hb8c2;
         4'h6d50 	:	val_out <= 4'hb8ab;
         4'h6d51 	:	val_out <= 4'hb8ab;
         4'h6d52 	:	val_out <= 4'hb8ab;
         4'h6d53 	:	val_out <= 4'hb8ab;
         4'h6d58 	:	val_out <= 4'hb895;
         4'h6d59 	:	val_out <= 4'hb895;
         4'h6d5a 	:	val_out <= 4'hb895;
         4'h6d5b 	:	val_out <= 4'hb895;
         4'h6d60 	:	val_out <= 4'hb87e;
         4'h6d61 	:	val_out <= 4'hb87e;
         4'h6d62 	:	val_out <= 4'hb87e;
         4'h6d63 	:	val_out <= 4'hb87e;
         4'h6d68 	:	val_out <= 4'hb868;
         4'h6d69 	:	val_out <= 4'hb868;
         4'h6d6a 	:	val_out <= 4'hb868;
         4'h6d6b 	:	val_out <= 4'hb868;
         4'h6d70 	:	val_out <= 4'hb851;
         4'h6d71 	:	val_out <= 4'hb851;
         4'h6d72 	:	val_out <= 4'hb851;
         4'h6d73 	:	val_out <= 4'hb851;
         4'h6d78 	:	val_out <= 4'hb83b;
         4'h6d79 	:	val_out <= 4'hb83b;
         4'h6d7a 	:	val_out <= 4'hb83b;
         4'h6d7b 	:	val_out <= 4'hb83b;
         4'h6d80 	:	val_out <= 4'hb824;
         4'h6d81 	:	val_out <= 4'hb824;
         4'h6d82 	:	val_out <= 4'hb824;
         4'h6d83 	:	val_out <= 4'hb824;
         4'h6d88 	:	val_out <= 4'hb80d;
         4'h6d89 	:	val_out <= 4'hb80d;
         4'h6d8a 	:	val_out <= 4'hb80d;
         4'h6d8b 	:	val_out <= 4'hb80d;
         4'h6d90 	:	val_out <= 4'hb7f7;
         4'h6d91 	:	val_out <= 4'hb7f7;
         4'h6d92 	:	val_out <= 4'hb7f7;
         4'h6d93 	:	val_out <= 4'hb7f7;
         4'h6d98 	:	val_out <= 4'hb7e0;
         4'h6d99 	:	val_out <= 4'hb7e0;
         4'h6d9a 	:	val_out <= 4'hb7e0;
         4'h6d9b 	:	val_out <= 4'hb7e0;
         4'h6da0 	:	val_out <= 4'hb7ca;
         4'h6da1 	:	val_out <= 4'hb7ca;
         4'h6da2 	:	val_out <= 4'hb7ca;
         4'h6da3 	:	val_out <= 4'hb7ca;
         4'h6da8 	:	val_out <= 4'hb7b3;
         4'h6da9 	:	val_out <= 4'hb7b3;
         4'h6daa 	:	val_out <= 4'hb7b3;
         4'h6dab 	:	val_out <= 4'hb7b3;
         4'h6db0 	:	val_out <= 4'hb79c;
         4'h6db1 	:	val_out <= 4'hb79c;
         4'h6db2 	:	val_out <= 4'hb79c;
         4'h6db3 	:	val_out <= 4'hb79c;
         4'h6db8 	:	val_out <= 4'hb786;
         4'h6db9 	:	val_out <= 4'hb786;
         4'h6dba 	:	val_out <= 4'hb786;
         4'h6dbb 	:	val_out <= 4'hb786;
         4'h6dc0 	:	val_out <= 4'hb76f;
         4'h6dc1 	:	val_out <= 4'hb76f;
         4'h6dc2 	:	val_out <= 4'hb76f;
         4'h6dc3 	:	val_out <= 4'hb76f;
         4'h6dc8 	:	val_out <= 4'hb758;
         4'h6dc9 	:	val_out <= 4'hb758;
         4'h6dca 	:	val_out <= 4'hb758;
         4'h6dcb 	:	val_out <= 4'hb758;
         4'h6dd0 	:	val_out <= 4'hb742;
         4'h6dd1 	:	val_out <= 4'hb742;
         4'h6dd2 	:	val_out <= 4'hb742;
         4'h6dd3 	:	val_out <= 4'hb742;
         4'h6dd8 	:	val_out <= 4'hb72b;
         4'h6dd9 	:	val_out <= 4'hb72b;
         4'h6dda 	:	val_out <= 4'hb72b;
         4'h6ddb 	:	val_out <= 4'hb72b;
         4'h6de0 	:	val_out <= 4'hb714;
         4'h6de1 	:	val_out <= 4'hb714;
         4'h6de2 	:	val_out <= 4'hb714;
         4'h6de3 	:	val_out <= 4'hb714;
         4'h6de8 	:	val_out <= 4'hb6fe;
         4'h6de9 	:	val_out <= 4'hb6fe;
         4'h6dea 	:	val_out <= 4'hb6fe;
         4'h6deb 	:	val_out <= 4'hb6fe;
         4'h6df0 	:	val_out <= 4'hb6e7;
         4'h6df1 	:	val_out <= 4'hb6e7;
         4'h6df2 	:	val_out <= 4'hb6e7;
         4'h6df3 	:	val_out <= 4'hb6e7;
         4'h6df8 	:	val_out <= 4'hb6d0;
         4'h6df9 	:	val_out <= 4'hb6d0;
         4'h6dfa 	:	val_out <= 4'hb6d0;
         4'h6dfb 	:	val_out <= 4'hb6d0;
         4'h6e00 	:	val_out <= 4'hb6ba;
         4'h6e01 	:	val_out <= 4'hb6ba;
         4'h6e02 	:	val_out <= 4'hb6ba;
         4'h6e03 	:	val_out <= 4'hb6ba;
         4'h6e08 	:	val_out <= 4'hb6a3;
         4'h6e09 	:	val_out <= 4'hb6a3;
         4'h6e0a 	:	val_out <= 4'hb6a3;
         4'h6e0b 	:	val_out <= 4'hb6a3;
         4'h6e10 	:	val_out <= 4'hb68c;
         4'h6e11 	:	val_out <= 4'hb68c;
         4'h6e12 	:	val_out <= 4'hb68c;
         4'h6e13 	:	val_out <= 4'hb68c;
         4'h6e18 	:	val_out <= 4'hb675;
         4'h6e19 	:	val_out <= 4'hb675;
         4'h6e1a 	:	val_out <= 4'hb675;
         4'h6e1b 	:	val_out <= 4'hb675;
         4'h6e20 	:	val_out <= 4'hb65f;
         4'h6e21 	:	val_out <= 4'hb65f;
         4'h6e22 	:	val_out <= 4'hb65f;
         4'h6e23 	:	val_out <= 4'hb65f;
         4'h6e28 	:	val_out <= 4'hb648;
         4'h6e29 	:	val_out <= 4'hb648;
         4'h6e2a 	:	val_out <= 4'hb648;
         4'h6e2b 	:	val_out <= 4'hb648;
         4'h6e30 	:	val_out <= 4'hb631;
         4'h6e31 	:	val_out <= 4'hb631;
         4'h6e32 	:	val_out <= 4'hb631;
         4'h6e33 	:	val_out <= 4'hb631;
         4'h6e38 	:	val_out <= 4'hb61a;
         4'h6e39 	:	val_out <= 4'hb61a;
         4'h6e3a 	:	val_out <= 4'hb61a;
         4'h6e3b 	:	val_out <= 4'hb61a;
         4'h6e40 	:	val_out <= 4'hb604;
         4'h6e41 	:	val_out <= 4'hb604;
         4'h6e42 	:	val_out <= 4'hb604;
         4'h6e43 	:	val_out <= 4'hb604;
         4'h6e48 	:	val_out <= 4'hb5ed;
         4'h6e49 	:	val_out <= 4'hb5ed;
         4'h6e4a 	:	val_out <= 4'hb5ed;
         4'h6e4b 	:	val_out <= 4'hb5ed;
         4'h6e50 	:	val_out <= 4'hb5d6;
         4'h6e51 	:	val_out <= 4'hb5d6;
         4'h6e52 	:	val_out <= 4'hb5d6;
         4'h6e53 	:	val_out <= 4'hb5d6;
         4'h6e58 	:	val_out <= 4'hb5bf;
         4'h6e59 	:	val_out <= 4'hb5bf;
         4'h6e5a 	:	val_out <= 4'hb5bf;
         4'h6e5b 	:	val_out <= 4'hb5bf;
         4'h6e60 	:	val_out <= 4'hb5a8;
         4'h6e61 	:	val_out <= 4'hb5a8;
         4'h6e62 	:	val_out <= 4'hb5a8;
         4'h6e63 	:	val_out <= 4'hb5a8;
         4'h6e68 	:	val_out <= 4'hb592;
         4'h6e69 	:	val_out <= 4'hb592;
         4'h6e6a 	:	val_out <= 4'hb592;
         4'h6e6b 	:	val_out <= 4'hb592;
         4'h6e70 	:	val_out <= 4'hb57b;
         4'h6e71 	:	val_out <= 4'hb57b;
         4'h6e72 	:	val_out <= 4'hb57b;
         4'h6e73 	:	val_out <= 4'hb57b;
         4'h6e78 	:	val_out <= 4'hb564;
         4'h6e79 	:	val_out <= 4'hb564;
         4'h6e7a 	:	val_out <= 4'hb564;
         4'h6e7b 	:	val_out <= 4'hb564;
         4'h6e80 	:	val_out <= 4'hb54d;
         4'h6e81 	:	val_out <= 4'hb54d;
         4'h6e82 	:	val_out <= 4'hb54d;
         4'h6e83 	:	val_out <= 4'hb54d;
         4'h6e88 	:	val_out <= 4'hb536;
         4'h6e89 	:	val_out <= 4'hb536;
         4'h6e8a 	:	val_out <= 4'hb536;
         4'h6e8b 	:	val_out <= 4'hb536;
         4'h6e90 	:	val_out <= 4'hb51f;
         4'h6e91 	:	val_out <= 4'hb51f;
         4'h6e92 	:	val_out <= 4'hb51f;
         4'h6e93 	:	val_out <= 4'hb51f;
         4'h6e98 	:	val_out <= 4'hb508;
         4'h6e99 	:	val_out <= 4'hb508;
         4'h6e9a 	:	val_out <= 4'hb508;
         4'h6e9b 	:	val_out <= 4'hb508;
         4'h6ea0 	:	val_out <= 4'hb4f2;
         4'h6ea1 	:	val_out <= 4'hb4f2;
         4'h6ea2 	:	val_out <= 4'hb4f2;
         4'h6ea3 	:	val_out <= 4'hb4f2;
         4'h6ea8 	:	val_out <= 4'hb4db;
         4'h6ea9 	:	val_out <= 4'hb4db;
         4'h6eaa 	:	val_out <= 4'hb4db;
         4'h6eab 	:	val_out <= 4'hb4db;
         4'h6eb0 	:	val_out <= 4'hb4c4;
         4'h6eb1 	:	val_out <= 4'hb4c4;
         4'h6eb2 	:	val_out <= 4'hb4c4;
         4'h6eb3 	:	val_out <= 4'hb4c4;
         4'h6eb8 	:	val_out <= 4'hb4ad;
         4'h6eb9 	:	val_out <= 4'hb4ad;
         4'h6eba 	:	val_out <= 4'hb4ad;
         4'h6ebb 	:	val_out <= 4'hb4ad;
         4'h6ec0 	:	val_out <= 4'hb496;
         4'h6ec1 	:	val_out <= 4'hb496;
         4'h6ec2 	:	val_out <= 4'hb496;
         4'h6ec3 	:	val_out <= 4'hb496;
         4'h6ec8 	:	val_out <= 4'hb47f;
         4'h6ec9 	:	val_out <= 4'hb47f;
         4'h6eca 	:	val_out <= 4'hb47f;
         4'h6ecb 	:	val_out <= 4'hb47f;
         4'h6ed0 	:	val_out <= 4'hb468;
         4'h6ed1 	:	val_out <= 4'hb468;
         4'h6ed2 	:	val_out <= 4'hb468;
         4'h6ed3 	:	val_out <= 4'hb468;
         4'h6ed8 	:	val_out <= 4'hb451;
         4'h6ed9 	:	val_out <= 4'hb451;
         4'h6eda 	:	val_out <= 4'hb451;
         4'h6edb 	:	val_out <= 4'hb451;
         4'h6ee0 	:	val_out <= 4'hb43a;
         4'h6ee1 	:	val_out <= 4'hb43a;
         4'h6ee2 	:	val_out <= 4'hb43a;
         4'h6ee3 	:	val_out <= 4'hb43a;
         4'h6ee8 	:	val_out <= 4'hb423;
         4'h6ee9 	:	val_out <= 4'hb423;
         4'h6eea 	:	val_out <= 4'hb423;
         4'h6eeb 	:	val_out <= 4'hb423;
         4'h6ef0 	:	val_out <= 4'hb40c;
         4'h6ef1 	:	val_out <= 4'hb40c;
         4'h6ef2 	:	val_out <= 4'hb40c;
         4'h6ef3 	:	val_out <= 4'hb40c;
         4'h6ef8 	:	val_out <= 4'hb3f5;
         4'h6ef9 	:	val_out <= 4'hb3f5;
         4'h6efa 	:	val_out <= 4'hb3f5;
         4'h6efb 	:	val_out <= 4'hb3f5;
         4'h6f00 	:	val_out <= 4'hb3de;
         4'h6f01 	:	val_out <= 4'hb3de;
         4'h6f02 	:	val_out <= 4'hb3de;
         4'h6f03 	:	val_out <= 4'hb3de;
         4'h6f08 	:	val_out <= 4'hb3c7;
         4'h6f09 	:	val_out <= 4'hb3c7;
         4'h6f0a 	:	val_out <= 4'hb3c7;
         4'h6f0b 	:	val_out <= 4'hb3c7;
         4'h6f10 	:	val_out <= 4'hb3b0;
         4'h6f11 	:	val_out <= 4'hb3b0;
         4'h6f12 	:	val_out <= 4'hb3b0;
         4'h6f13 	:	val_out <= 4'hb3b0;
         4'h6f18 	:	val_out <= 4'hb399;
         4'h6f19 	:	val_out <= 4'hb399;
         4'h6f1a 	:	val_out <= 4'hb399;
         4'h6f1b 	:	val_out <= 4'hb399;
         4'h6f20 	:	val_out <= 4'hb382;
         4'h6f21 	:	val_out <= 4'hb382;
         4'h6f22 	:	val_out <= 4'hb382;
         4'h6f23 	:	val_out <= 4'hb382;
         4'h6f28 	:	val_out <= 4'hb36b;
         4'h6f29 	:	val_out <= 4'hb36b;
         4'h6f2a 	:	val_out <= 4'hb36b;
         4'h6f2b 	:	val_out <= 4'hb36b;
         4'h6f30 	:	val_out <= 4'hb354;
         4'h6f31 	:	val_out <= 4'hb354;
         4'h6f32 	:	val_out <= 4'hb354;
         4'h6f33 	:	val_out <= 4'hb354;
         4'h6f38 	:	val_out <= 4'hb33d;
         4'h6f39 	:	val_out <= 4'hb33d;
         4'h6f3a 	:	val_out <= 4'hb33d;
         4'h6f3b 	:	val_out <= 4'hb33d;
         4'h6f40 	:	val_out <= 4'hb326;
         4'h6f41 	:	val_out <= 4'hb326;
         4'h6f42 	:	val_out <= 4'hb326;
         4'h6f43 	:	val_out <= 4'hb326;
         4'h6f48 	:	val_out <= 4'hb30f;
         4'h6f49 	:	val_out <= 4'hb30f;
         4'h6f4a 	:	val_out <= 4'hb30f;
         4'h6f4b 	:	val_out <= 4'hb30f;
         4'h6f50 	:	val_out <= 4'hb2f8;
         4'h6f51 	:	val_out <= 4'hb2f8;
         4'h6f52 	:	val_out <= 4'hb2f8;
         4'h6f53 	:	val_out <= 4'hb2f8;
         4'h6f58 	:	val_out <= 4'hb2e1;
         4'h6f59 	:	val_out <= 4'hb2e1;
         4'h6f5a 	:	val_out <= 4'hb2e1;
         4'h6f5b 	:	val_out <= 4'hb2e1;
         4'h6f60 	:	val_out <= 4'hb2ca;
         4'h6f61 	:	val_out <= 4'hb2ca;
         4'h6f62 	:	val_out <= 4'hb2ca;
         4'h6f63 	:	val_out <= 4'hb2ca;
         4'h6f68 	:	val_out <= 4'hb2b3;
         4'h6f69 	:	val_out <= 4'hb2b3;
         4'h6f6a 	:	val_out <= 4'hb2b3;
         4'h6f6b 	:	val_out <= 4'hb2b3;
         4'h6f70 	:	val_out <= 4'hb29c;
         4'h6f71 	:	val_out <= 4'hb29c;
         4'h6f72 	:	val_out <= 4'hb29c;
         4'h6f73 	:	val_out <= 4'hb29c;
         4'h6f78 	:	val_out <= 4'hb285;
         4'h6f79 	:	val_out <= 4'hb285;
         4'h6f7a 	:	val_out <= 4'hb285;
         4'h6f7b 	:	val_out <= 4'hb285;
         4'h6f80 	:	val_out <= 4'hb26e;
         4'h6f81 	:	val_out <= 4'hb26e;
         4'h6f82 	:	val_out <= 4'hb26e;
         4'h6f83 	:	val_out <= 4'hb26e;
         4'h6f88 	:	val_out <= 4'hb257;
         4'h6f89 	:	val_out <= 4'hb257;
         4'h6f8a 	:	val_out <= 4'hb257;
         4'h6f8b 	:	val_out <= 4'hb257;
         4'h6f90 	:	val_out <= 4'hb240;
         4'h6f91 	:	val_out <= 4'hb240;
         4'h6f92 	:	val_out <= 4'hb240;
         4'h6f93 	:	val_out <= 4'hb240;
         4'h6f98 	:	val_out <= 4'hb228;
         4'h6f99 	:	val_out <= 4'hb228;
         4'h6f9a 	:	val_out <= 4'hb228;
         4'h6f9b 	:	val_out <= 4'hb228;
         4'h6fa0 	:	val_out <= 4'hb211;
         4'h6fa1 	:	val_out <= 4'hb211;
         4'h6fa2 	:	val_out <= 4'hb211;
         4'h6fa3 	:	val_out <= 4'hb211;
         4'h6fa8 	:	val_out <= 4'hb1fa;
         4'h6fa9 	:	val_out <= 4'hb1fa;
         4'h6faa 	:	val_out <= 4'hb1fa;
         4'h6fab 	:	val_out <= 4'hb1fa;
         4'h6fb0 	:	val_out <= 4'hb1e3;
         4'h6fb1 	:	val_out <= 4'hb1e3;
         4'h6fb2 	:	val_out <= 4'hb1e3;
         4'h6fb3 	:	val_out <= 4'hb1e3;
         4'h6fb8 	:	val_out <= 4'hb1cc;
         4'h6fb9 	:	val_out <= 4'hb1cc;
         4'h6fba 	:	val_out <= 4'hb1cc;
         4'h6fbb 	:	val_out <= 4'hb1cc;
         4'h6fc0 	:	val_out <= 4'hb1b5;
         4'h6fc1 	:	val_out <= 4'hb1b5;
         4'h6fc2 	:	val_out <= 4'hb1b5;
         4'h6fc3 	:	val_out <= 4'hb1b5;
         4'h6fc8 	:	val_out <= 4'hb19e;
         4'h6fc9 	:	val_out <= 4'hb19e;
         4'h6fca 	:	val_out <= 4'hb19e;
         4'h6fcb 	:	val_out <= 4'hb19e;
         4'h6fd0 	:	val_out <= 4'hb186;
         4'h6fd1 	:	val_out <= 4'hb186;
         4'h6fd2 	:	val_out <= 4'hb186;
         4'h6fd3 	:	val_out <= 4'hb186;
         4'h6fd8 	:	val_out <= 4'hb16f;
         4'h6fd9 	:	val_out <= 4'hb16f;
         4'h6fda 	:	val_out <= 4'hb16f;
         4'h6fdb 	:	val_out <= 4'hb16f;
         4'h6fe0 	:	val_out <= 4'hb158;
         4'h6fe1 	:	val_out <= 4'hb158;
         4'h6fe2 	:	val_out <= 4'hb158;
         4'h6fe3 	:	val_out <= 4'hb158;
         4'h6fe8 	:	val_out <= 4'hb141;
         4'h6fe9 	:	val_out <= 4'hb141;
         4'h6fea 	:	val_out <= 4'hb141;
         4'h6feb 	:	val_out <= 4'hb141;
         4'h6ff0 	:	val_out <= 4'hb12a;
         4'h6ff1 	:	val_out <= 4'hb12a;
         4'h6ff2 	:	val_out <= 4'hb12a;
         4'h6ff3 	:	val_out <= 4'hb12a;
         4'h6ff8 	:	val_out <= 4'hb112;
         4'h6ff9 	:	val_out <= 4'hb112;
         4'h6ffa 	:	val_out <= 4'hb112;
         4'h6ffb 	:	val_out <= 4'hb112;
         4'h7000 	:	val_out <= 4'hb0fb;
         4'h7001 	:	val_out <= 4'hb0fb;
         4'h7002 	:	val_out <= 4'hb0fb;
         4'h7003 	:	val_out <= 4'hb0fb;
         4'h7008 	:	val_out <= 4'hb0e4;
         4'h7009 	:	val_out <= 4'hb0e4;
         4'h700a 	:	val_out <= 4'hb0e4;
         4'h700b 	:	val_out <= 4'hb0e4;
         4'h7010 	:	val_out <= 4'hb0cd;
         4'h7011 	:	val_out <= 4'hb0cd;
         4'h7012 	:	val_out <= 4'hb0cd;
         4'h7013 	:	val_out <= 4'hb0cd;
         4'h7018 	:	val_out <= 4'hb0b6;
         4'h7019 	:	val_out <= 4'hb0b6;
         4'h701a 	:	val_out <= 4'hb0b6;
         4'h701b 	:	val_out <= 4'hb0b6;
         4'h7020 	:	val_out <= 4'hb09e;
         4'h7021 	:	val_out <= 4'hb09e;
         4'h7022 	:	val_out <= 4'hb09e;
         4'h7023 	:	val_out <= 4'hb09e;
         4'h7028 	:	val_out <= 4'hb087;
         4'h7029 	:	val_out <= 4'hb087;
         4'h702a 	:	val_out <= 4'hb087;
         4'h702b 	:	val_out <= 4'hb087;
         4'h7030 	:	val_out <= 4'hb070;
         4'h7031 	:	val_out <= 4'hb070;
         4'h7032 	:	val_out <= 4'hb070;
         4'h7033 	:	val_out <= 4'hb070;
         4'h7038 	:	val_out <= 4'hb059;
         4'h7039 	:	val_out <= 4'hb059;
         4'h703a 	:	val_out <= 4'hb059;
         4'h703b 	:	val_out <= 4'hb059;
         4'h7040 	:	val_out <= 4'hb041;
         4'h7041 	:	val_out <= 4'hb041;
         4'h7042 	:	val_out <= 4'hb041;
         4'h7043 	:	val_out <= 4'hb041;
         4'h7048 	:	val_out <= 4'hb02a;
         4'h7049 	:	val_out <= 4'hb02a;
         4'h704a 	:	val_out <= 4'hb02a;
         4'h704b 	:	val_out <= 4'hb02a;
         4'h7050 	:	val_out <= 4'hb013;
         4'h7051 	:	val_out <= 4'hb013;
         4'h7052 	:	val_out <= 4'hb013;
         4'h7053 	:	val_out <= 4'hb013;
         4'h7058 	:	val_out <= 4'haffb;
         4'h7059 	:	val_out <= 4'haffb;
         4'h705a 	:	val_out <= 4'haffb;
         4'h705b 	:	val_out <= 4'haffb;
         4'h7060 	:	val_out <= 4'hafe4;
         4'h7061 	:	val_out <= 4'hafe4;
         4'h7062 	:	val_out <= 4'hafe4;
         4'h7063 	:	val_out <= 4'hafe4;
         4'h7068 	:	val_out <= 4'hafcd;
         4'h7069 	:	val_out <= 4'hafcd;
         4'h706a 	:	val_out <= 4'hafcd;
         4'h706b 	:	val_out <= 4'hafcd;
         4'h7070 	:	val_out <= 4'hafb5;
         4'h7071 	:	val_out <= 4'hafb5;
         4'h7072 	:	val_out <= 4'hafb5;
         4'h7073 	:	val_out <= 4'hafb5;
         4'h7078 	:	val_out <= 4'haf9e;
         4'h7079 	:	val_out <= 4'haf9e;
         4'h707a 	:	val_out <= 4'haf9e;
         4'h707b 	:	val_out <= 4'haf9e;
         4'h7080 	:	val_out <= 4'haf87;
         4'h7081 	:	val_out <= 4'haf87;
         4'h7082 	:	val_out <= 4'haf87;
         4'h7083 	:	val_out <= 4'haf87;
         4'h7088 	:	val_out <= 4'haf6f;
         4'h7089 	:	val_out <= 4'haf6f;
         4'h708a 	:	val_out <= 4'haf6f;
         4'h708b 	:	val_out <= 4'haf6f;
         4'h7090 	:	val_out <= 4'haf58;
         4'h7091 	:	val_out <= 4'haf58;
         4'h7092 	:	val_out <= 4'haf58;
         4'h7093 	:	val_out <= 4'haf58;
         4'h7098 	:	val_out <= 4'haf41;
         4'h7099 	:	val_out <= 4'haf41;
         4'h709a 	:	val_out <= 4'haf41;
         4'h709b 	:	val_out <= 4'haf41;
         4'h70a0 	:	val_out <= 4'haf29;
         4'h70a1 	:	val_out <= 4'haf29;
         4'h70a2 	:	val_out <= 4'haf29;
         4'h70a3 	:	val_out <= 4'haf29;
         4'h70a8 	:	val_out <= 4'haf12;
         4'h70a9 	:	val_out <= 4'haf12;
         4'h70aa 	:	val_out <= 4'haf12;
         4'h70ab 	:	val_out <= 4'haf12;
         4'h70b0 	:	val_out <= 4'haefb;
         4'h70b1 	:	val_out <= 4'haefb;
         4'h70b2 	:	val_out <= 4'haefb;
         4'h70b3 	:	val_out <= 4'haefb;
         4'h70b8 	:	val_out <= 4'haee3;
         4'h70b9 	:	val_out <= 4'haee3;
         4'h70ba 	:	val_out <= 4'haee3;
         4'h70bb 	:	val_out <= 4'haee3;
         4'h70c0 	:	val_out <= 4'haecc;
         4'h70c1 	:	val_out <= 4'haecc;
         4'h70c2 	:	val_out <= 4'haecc;
         4'h70c3 	:	val_out <= 4'haecc;
         4'h70c8 	:	val_out <= 4'haeb5;
         4'h70c9 	:	val_out <= 4'haeb5;
         4'h70ca 	:	val_out <= 4'haeb5;
         4'h70cb 	:	val_out <= 4'haeb5;
         4'h70d0 	:	val_out <= 4'hae9d;
         4'h70d1 	:	val_out <= 4'hae9d;
         4'h70d2 	:	val_out <= 4'hae9d;
         4'h70d3 	:	val_out <= 4'hae9d;
         4'h70d8 	:	val_out <= 4'hae86;
         4'h70d9 	:	val_out <= 4'hae86;
         4'h70da 	:	val_out <= 4'hae86;
         4'h70db 	:	val_out <= 4'hae86;
         4'h70e0 	:	val_out <= 4'hae6e;
         4'h70e1 	:	val_out <= 4'hae6e;
         4'h70e2 	:	val_out <= 4'hae6e;
         4'h70e3 	:	val_out <= 4'hae6e;
         4'h70e8 	:	val_out <= 4'hae57;
         4'h70e9 	:	val_out <= 4'hae57;
         4'h70ea 	:	val_out <= 4'hae57;
         4'h70eb 	:	val_out <= 4'hae57;
         4'h70f0 	:	val_out <= 4'hae3f;
         4'h70f1 	:	val_out <= 4'hae3f;
         4'h70f2 	:	val_out <= 4'hae3f;
         4'h70f3 	:	val_out <= 4'hae3f;
         4'h70f8 	:	val_out <= 4'hae28;
         4'h70f9 	:	val_out <= 4'hae28;
         4'h70fa 	:	val_out <= 4'hae28;
         4'h70fb 	:	val_out <= 4'hae28;
         4'h7100 	:	val_out <= 4'hae11;
         4'h7101 	:	val_out <= 4'hae11;
         4'h7102 	:	val_out <= 4'hae11;
         4'h7103 	:	val_out <= 4'hae11;
         4'h7108 	:	val_out <= 4'hadf9;
         4'h7109 	:	val_out <= 4'hadf9;
         4'h710a 	:	val_out <= 4'hadf9;
         4'h710b 	:	val_out <= 4'hadf9;
         4'h7110 	:	val_out <= 4'hade2;
         4'h7111 	:	val_out <= 4'hade2;
         4'h7112 	:	val_out <= 4'hade2;
         4'h7113 	:	val_out <= 4'hade2;
         4'h7118 	:	val_out <= 4'hadca;
         4'h7119 	:	val_out <= 4'hadca;
         4'h711a 	:	val_out <= 4'hadca;
         4'h711b 	:	val_out <= 4'hadca;
         4'h7120 	:	val_out <= 4'hadb3;
         4'h7121 	:	val_out <= 4'hadb3;
         4'h7122 	:	val_out <= 4'hadb3;
         4'h7123 	:	val_out <= 4'hadb3;
         4'h7128 	:	val_out <= 4'had9b;
         4'h7129 	:	val_out <= 4'had9b;
         4'h712a 	:	val_out <= 4'had9b;
         4'h712b 	:	val_out <= 4'had9b;
         4'h7130 	:	val_out <= 4'had84;
         4'h7131 	:	val_out <= 4'had84;
         4'h7132 	:	val_out <= 4'had84;
         4'h7133 	:	val_out <= 4'had84;
         4'h7138 	:	val_out <= 4'had6c;
         4'h7139 	:	val_out <= 4'had6c;
         4'h713a 	:	val_out <= 4'had6c;
         4'h713b 	:	val_out <= 4'had6c;
         4'h7140 	:	val_out <= 4'had55;
         4'h7141 	:	val_out <= 4'had55;
         4'h7142 	:	val_out <= 4'had55;
         4'h7143 	:	val_out <= 4'had55;
         4'h7148 	:	val_out <= 4'had3d;
         4'h7149 	:	val_out <= 4'had3d;
         4'h714a 	:	val_out <= 4'had3d;
         4'h714b 	:	val_out <= 4'had3d;
         4'h7150 	:	val_out <= 4'had26;
         4'h7151 	:	val_out <= 4'had26;
         4'h7152 	:	val_out <= 4'had26;
         4'h7153 	:	val_out <= 4'had26;
         4'h7158 	:	val_out <= 4'had0e;
         4'h7159 	:	val_out <= 4'had0e;
         4'h715a 	:	val_out <= 4'had0e;
         4'h715b 	:	val_out <= 4'had0e;
         4'h7160 	:	val_out <= 4'hacf7;
         4'h7161 	:	val_out <= 4'hacf7;
         4'h7162 	:	val_out <= 4'hacf7;
         4'h7163 	:	val_out <= 4'hacf7;
         4'h7168 	:	val_out <= 4'hacdf;
         4'h7169 	:	val_out <= 4'hacdf;
         4'h716a 	:	val_out <= 4'hacdf;
         4'h716b 	:	val_out <= 4'hacdf;
         4'h7170 	:	val_out <= 4'hacc8;
         4'h7171 	:	val_out <= 4'hacc8;
         4'h7172 	:	val_out <= 4'hacc8;
         4'h7173 	:	val_out <= 4'hacc8;
         4'h7178 	:	val_out <= 4'hacb0;
         4'h7179 	:	val_out <= 4'hacb0;
         4'h717a 	:	val_out <= 4'hacb0;
         4'h717b 	:	val_out <= 4'hacb0;
         4'h7180 	:	val_out <= 4'hac98;
         4'h7181 	:	val_out <= 4'hac98;
         4'h7182 	:	val_out <= 4'hac98;
         4'h7183 	:	val_out <= 4'hac98;
         4'h7188 	:	val_out <= 4'hac81;
         4'h7189 	:	val_out <= 4'hac81;
         4'h718a 	:	val_out <= 4'hac81;
         4'h718b 	:	val_out <= 4'hac81;
         4'h7190 	:	val_out <= 4'hac69;
         4'h7191 	:	val_out <= 4'hac69;
         4'h7192 	:	val_out <= 4'hac69;
         4'h7193 	:	val_out <= 4'hac69;
         4'h7198 	:	val_out <= 4'hac52;
         4'h7199 	:	val_out <= 4'hac52;
         4'h719a 	:	val_out <= 4'hac52;
         4'h719b 	:	val_out <= 4'hac52;
         4'h71a0 	:	val_out <= 4'hac3a;
         4'h71a1 	:	val_out <= 4'hac3a;
         4'h71a2 	:	val_out <= 4'hac3a;
         4'h71a3 	:	val_out <= 4'hac3a;
         4'h71a8 	:	val_out <= 4'hac23;
         4'h71a9 	:	val_out <= 4'hac23;
         4'h71aa 	:	val_out <= 4'hac23;
         4'h71ab 	:	val_out <= 4'hac23;
         4'h71b0 	:	val_out <= 4'hac0b;
         4'h71b1 	:	val_out <= 4'hac0b;
         4'h71b2 	:	val_out <= 4'hac0b;
         4'h71b3 	:	val_out <= 4'hac0b;
         4'h71b8 	:	val_out <= 4'habf3;
         4'h71b9 	:	val_out <= 4'habf3;
         4'h71ba 	:	val_out <= 4'habf3;
         4'h71bb 	:	val_out <= 4'habf3;
         4'h71c0 	:	val_out <= 4'habdc;
         4'h71c1 	:	val_out <= 4'habdc;
         4'h71c2 	:	val_out <= 4'habdc;
         4'h71c3 	:	val_out <= 4'habdc;
         4'h71c8 	:	val_out <= 4'habc4;
         4'h71c9 	:	val_out <= 4'habc4;
         4'h71ca 	:	val_out <= 4'habc4;
         4'h71cb 	:	val_out <= 4'habc4;
         4'h71d0 	:	val_out <= 4'habad;
         4'h71d1 	:	val_out <= 4'habad;
         4'h71d2 	:	val_out <= 4'habad;
         4'h71d3 	:	val_out <= 4'habad;
         4'h71d8 	:	val_out <= 4'hab95;
         4'h71d9 	:	val_out <= 4'hab95;
         4'h71da 	:	val_out <= 4'hab95;
         4'h71db 	:	val_out <= 4'hab95;
         4'h71e0 	:	val_out <= 4'hab7d;
         4'h71e1 	:	val_out <= 4'hab7d;
         4'h71e2 	:	val_out <= 4'hab7d;
         4'h71e3 	:	val_out <= 4'hab7d;
         4'h71e8 	:	val_out <= 4'hab66;
         4'h71e9 	:	val_out <= 4'hab66;
         4'h71ea 	:	val_out <= 4'hab66;
         4'h71eb 	:	val_out <= 4'hab66;
         4'h71f0 	:	val_out <= 4'hab4e;
         4'h71f1 	:	val_out <= 4'hab4e;
         4'h71f2 	:	val_out <= 4'hab4e;
         4'h71f3 	:	val_out <= 4'hab4e;
         4'h71f8 	:	val_out <= 4'hab36;
         4'h71f9 	:	val_out <= 4'hab36;
         4'h71fa 	:	val_out <= 4'hab36;
         4'h71fb 	:	val_out <= 4'hab36;
         4'h7200 	:	val_out <= 4'hab1f;
         4'h7201 	:	val_out <= 4'hab1f;
         4'h7202 	:	val_out <= 4'hab1f;
         4'h7203 	:	val_out <= 4'hab1f;
         4'h7208 	:	val_out <= 4'hab07;
         4'h7209 	:	val_out <= 4'hab07;
         4'h720a 	:	val_out <= 4'hab07;
         4'h720b 	:	val_out <= 4'hab07;
         4'h7210 	:	val_out <= 4'haaef;
         4'h7211 	:	val_out <= 4'haaef;
         4'h7212 	:	val_out <= 4'haaef;
         4'h7213 	:	val_out <= 4'haaef;
         4'h7218 	:	val_out <= 4'haad8;
         4'h7219 	:	val_out <= 4'haad8;
         4'h721a 	:	val_out <= 4'haad8;
         4'h721b 	:	val_out <= 4'haad8;
         4'h7220 	:	val_out <= 4'haac0;
         4'h7221 	:	val_out <= 4'haac0;
         4'h7222 	:	val_out <= 4'haac0;
         4'h7223 	:	val_out <= 4'haac0;
         4'h7228 	:	val_out <= 4'haaa8;
         4'h7229 	:	val_out <= 4'haaa8;
         4'h722a 	:	val_out <= 4'haaa8;
         4'h722b 	:	val_out <= 4'haaa8;
         4'h7230 	:	val_out <= 4'haa91;
         4'h7231 	:	val_out <= 4'haa91;
         4'h7232 	:	val_out <= 4'haa91;
         4'h7233 	:	val_out <= 4'haa91;
         4'h7238 	:	val_out <= 4'haa79;
         4'h7239 	:	val_out <= 4'haa79;
         4'h723a 	:	val_out <= 4'haa79;
         4'h723b 	:	val_out <= 4'haa79;
         4'h7240 	:	val_out <= 4'haa61;
         4'h7241 	:	val_out <= 4'haa61;
         4'h7242 	:	val_out <= 4'haa61;
         4'h7243 	:	val_out <= 4'haa61;
         4'h7248 	:	val_out <= 4'haa49;
         4'h7249 	:	val_out <= 4'haa49;
         4'h724a 	:	val_out <= 4'haa49;
         4'h724b 	:	val_out <= 4'haa49;
         4'h7250 	:	val_out <= 4'haa32;
         4'h7251 	:	val_out <= 4'haa32;
         4'h7252 	:	val_out <= 4'haa32;
         4'h7253 	:	val_out <= 4'haa32;
         4'h7258 	:	val_out <= 4'haa1a;
         4'h7259 	:	val_out <= 4'haa1a;
         4'h725a 	:	val_out <= 4'haa1a;
         4'h725b 	:	val_out <= 4'haa1a;
         4'h7260 	:	val_out <= 4'haa02;
         4'h7261 	:	val_out <= 4'haa02;
         4'h7262 	:	val_out <= 4'haa02;
         4'h7263 	:	val_out <= 4'haa02;
         4'h7268 	:	val_out <= 4'ha9eb;
         4'h7269 	:	val_out <= 4'ha9eb;
         4'h726a 	:	val_out <= 4'ha9eb;
         4'h726b 	:	val_out <= 4'ha9eb;
         4'h7270 	:	val_out <= 4'ha9d3;
         4'h7271 	:	val_out <= 4'ha9d3;
         4'h7272 	:	val_out <= 4'ha9d3;
         4'h7273 	:	val_out <= 4'ha9d3;
         4'h7278 	:	val_out <= 4'ha9bb;
         4'h7279 	:	val_out <= 4'ha9bb;
         4'h727a 	:	val_out <= 4'ha9bb;
         4'h727b 	:	val_out <= 4'ha9bb;
         4'h7280 	:	val_out <= 4'ha9a3;
         4'h7281 	:	val_out <= 4'ha9a3;
         4'h7282 	:	val_out <= 4'ha9a3;
         4'h7283 	:	val_out <= 4'ha9a3;
         4'h7288 	:	val_out <= 4'ha98b;
         4'h7289 	:	val_out <= 4'ha98b;
         4'h728a 	:	val_out <= 4'ha98b;
         4'h728b 	:	val_out <= 4'ha98b;
         4'h7290 	:	val_out <= 4'ha974;
         4'h7291 	:	val_out <= 4'ha974;
         4'h7292 	:	val_out <= 4'ha974;
         4'h7293 	:	val_out <= 4'ha974;
         4'h7298 	:	val_out <= 4'ha95c;
         4'h7299 	:	val_out <= 4'ha95c;
         4'h729a 	:	val_out <= 4'ha95c;
         4'h729b 	:	val_out <= 4'ha95c;
         4'h72a0 	:	val_out <= 4'ha944;
         4'h72a1 	:	val_out <= 4'ha944;
         4'h72a2 	:	val_out <= 4'ha944;
         4'h72a3 	:	val_out <= 4'ha944;
         4'h72a8 	:	val_out <= 4'ha92c;
         4'h72a9 	:	val_out <= 4'ha92c;
         4'h72aa 	:	val_out <= 4'ha92c;
         4'h72ab 	:	val_out <= 4'ha92c;
         4'h72b0 	:	val_out <= 4'ha915;
         4'h72b1 	:	val_out <= 4'ha915;
         4'h72b2 	:	val_out <= 4'ha915;
         4'h72b3 	:	val_out <= 4'ha915;
         4'h72b8 	:	val_out <= 4'ha8fd;
         4'h72b9 	:	val_out <= 4'ha8fd;
         4'h72ba 	:	val_out <= 4'ha8fd;
         4'h72bb 	:	val_out <= 4'ha8fd;
         4'h72c0 	:	val_out <= 4'ha8e5;
         4'h72c1 	:	val_out <= 4'ha8e5;
         4'h72c2 	:	val_out <= 4'ha8e5;
         4'h72c3 	:	val_out <= 4'ha8e5;
         4'h72c8 	:	val_out <= 4'ha8cd;
         4'h72c9 	:	val_out <= 4'ha8cd;
         4'h72ca 	:	val_out <= 4'ha8cd;
         4'h72cb 	:	val_out <= 4'ha8cd;
         4'h72d0 	:	val_out <= 4'ha8b5;
         4'h72d1 	:	val_out <= 4'ha8b5;
         4'h72d2 	:	val_out <= 4'ha8b5;
         4'h72d3 	:	val_out <= 4'ha8b5;
         4'h72d8 	:	val_out <= 4'ha89d;
         4'h72d9 	:	val_out <= 4'ha89d;
         4'h72da 	:	val_out <= 4'ha89d;
         4'h72db 	:	val_out <= 4'ha89d;
         4'h72e0 	:	val_out <= 4'ha886;
         4'h72e1 	:	val_out <= 4'ha886;
         4'h72e2 	:	val_out <= 4'ha886;
         4'h72e3 	:	val_out <= 4'ha886;
         4'h72e8 	:	val_out <= 4'ha86e;
         4'h72e9 	:	val_out <= 4'ha86e;
         4'h72ea 	:	val_out <= 4'ha86e;
         4'h72eb 	:	val_out <= 4'ha86e;
         4'h72f0 	:	val_out <= 4'ha856;
         4'h72f1 	:	val_out <= 4'ha856;
         4'h72f2 	:	val_out <= 4'ha856;
         4'h72f3 	:	val_out <= 4'ha856;
         4'h72f8 	:	val_out <= 4'ha83e;
         4'h72f9 	:	val_out <= 4'ha83e;
         4'h72fa 	:	val_out <= 4'ha83e;
         4'h72fb 	:	val_out <= 4'ha83e;
         4'h7300 	:	val_out <= 4'ha826;
         4'h7301 	:	val_out <= 4'ha826;
         4'h7302 	:	val_out <= 4'ha826;
         4'h7303 	:	val_out <= 4'ha826;
         4'h7308 	:	val_out <= 4'ha80e;
         4'h7309 	:	val_out <= 4'ha80e;
         4'h730a 	:	val_out <= 4'ha80e;
         4'h730b 	:	val_out <= 4'ha80e;
         4'h7310 	:	val_out <= 4'ha7f6;
         4'h7311 	:	val_out <= 4'ha7f6;
         4'h7312 	:	val_out <= 4'ha7f6;
         4'h7313 	:	val_out <= 4'ha7f6;
         4'h7318 	:	val_out <= 4'ha7df;
         4'h7319 	:	val_out <= 4'ha7df;
         4'h731a 	:	val_out <= 4'ha7df;
         4'h731b 	:	val_out <= 4'ha7df;
         4'h7320 	:	val_out <= 4'ha7c7;
         4'h7321 	:	val_out <= 4'ha7c7;
         4'h7322 	:	val_out <= 4'ha7c7;
         4'h7323 	:	val_out <= 4'ha7c7;
         4'h7328 	:	val_out <= 4'ha7af;
         4'h7329 	:	val_out <= 4'ha7af;
         4'h732a 	:	val_out <= 4'ha7af;
         4'h732b 	:	val_out <= 4'ha7af;
         4'h7330 	:	val_out <= 4'ha797;
         4'h7331 	:	val_out <= 4'ha797;
         4'h7332 	:	val_out <= 4'ha797;
         4'h7333 	:	val_out <= 4'ha797;
         4'h7338 	:	val_out <= 4'ha77f;
         4'h7339 	:	val_out <= 4'ha77f;
         4'h733a 	:	val_out <= 4'ha77f;
         4'h733b 	:	val_out <= 4'ha77f;
         4'h7340 	:	val_out <= 4'ha767;
         4'h7341 	:	val_out <= 4'ha767;
         4'h7342 	:	val_out <= 4'ha767;
         4'h7343 	:	val_out <= 4'ha767;
         4'h7348 	:	val_out <= 4'ha74f;
         4'h7349 	:	val_out <= 4'ha74f;
         4'h734a 	:	val_out <= 4'ha74f;
         4'h734b 	:	val_out <= 4'ha74f;
         4'h7350 	:	val_out <= 4'ha737;
         4'h7351 	:	val_out <= 4'ha737;
         4'h7352 	:	val_out <= 4'ha737;
         4'h7353 	:	val_out <= 4'ha737;
         4'h7358 	:	val_out <= 4'ha71f;
         4'h7359 	:	val_out <= 4'ha71f;
         4'h735a 	:	val_out <= 4'ha71f;
         4'h735b 	:	val_out <= 4'ha71f;
         4'h7360 	:	val_out <= 4'ha707;
         4'h7361 	:	val_out <= 4'ha707;
         4'h7362 	:	val_out <= 4'ha707;
         4'h7363 	:	val_out <= 4'ha707;
         4'h7368 	:	val_out <= 4'ha6ef;
         4'h7369 	:	val_out <= 4'ha6ef;
         4'h736a 	:	val_out <= 4'ha6ef;
         4'h736b 	:	val_out <= 4'ha6ef;
         4'h7370 	:	val_out <= 4'ha6d8;
         4'h7371 	:	val_out <= 4'ha6d8;
         4'h7372 	:	val_out <= 4'ha6d8;
         4'h7373 	:	val_out <= 4'ha6d8;
         4'h7378 	:	val_out <= 4'ha6c0;
         4'h7379 	:	val_out <= 4'ha6c0;
         4'h737a 	:	val_out <= 4'ha6c0;
         4'h737b 	:	val_out <= 4'ha6c0;
         4'h7380 	:	val_out <= 4'ha6a8;
         4'h7381 	:	val_out <= 4'ha6a8;
         4'h7382 	:	val_out <= 4'ha6a8;
         4'h7383 	:	val_out <= 4'ha6a8;
         4'h7388 	:	val_out <= 4'ha690;
         4'h7389 	:	val_out <= 4'ha690;
         4'h738a 	:	val_out <= 4'ha690;
         4'h738b 	:	val_out <= 4'ha690;
         4'h7390 	:	val_out <= 4'ha678;
         4'h7391 	:	val_out <= 4'ha678;
         4'h7392 	:	val_out <= 4'ha678;
         4'h7393 	:	val_out <= 4'ha678;
         4'h7398 	:	val_out <= 4'ha660;
         4'h7399 	:	val_out <= 4'ha660;
         4'h739a 	:	val_out <= 4'ha660;
         4'h739b 	:	val_out <= 4'ha660;
         4'h73a0 	:	val_out <= 4'ha648;
         4'h73a1 	:	val_out <= 4'ha648;
         4'h73a2 	:	val_out <= 4'ha648;
         4'h73a3 	:	val_out <= 4'ha648;
         4'h73a8 	:	val_out <= 4'ha630;
         4'h73a9 	:	val_out <= 4'ha630;
         4'h73aa 	:	val_out <= 4'ha630;
         4'h73ab 	:	val_out <= 4'ha630;
         4'h73b0 	:	val_out <= 4'ha618;
         4'h73b1 	:	val_out <= 4'ha618;
         4'h73b2 	:	val_out <= 4'ha618;
         4'h73b3 	:	val_out <= 4'ha618;
         4'h73b8 	:	val_out <= 4'ha600;
         4'h73b9 	:	val_out <= 4'ha600;
         4'h73ba 	:	val_out <= 4'ha600;
         4'h73bb 	:	val_out <= 4'ha600;
         4'h73c0 	:	val_out <= 4'ha5e8;
         4'h73c1 	:	val_out <= 4'ha5e8;
         4'h73c2 	:	val_out <= 4'ha5e8;
         4'h73c3 	:	val_out <= 4'ha5e8;
         4'h73c8 	:	val_out <= 4'ha5d0;
         4'h73c9 	:	val_out <= 4'ha5d0;
         4'h73ca 	:	val_out <= 4'ha5d0;
         4'h73cb 	:	val_out <= 4'ha5d0;
         4'h73d0 	:	val_out <= 4'ha5b8;
         4'h73d1 	:	val_out <= 4'ha5b8;
         4'h73d2 	:	val_out <= 4'ha5b8;
         4'h73d3 	:	val_out <= 4'ha5b8;
         4'h73d8 	:	val_out <= 4'ha5a0;
         4'h73d9 	:	val_out <= 4'ha5a0;
         4'h73da 	:	val_out <= 4'ha5a0;
         4'h73db 	:	val_out <= 4'ha5a0;
         4'h73e0 	:	val_out <= 4'ha588;
         4'h73e1 	:	val_out <= 4'ha588;
         4'h73e2 	:	val_out <= 4'ha588;
         4'h73e3 	:	val_out <= 4'ha588;
         4'h73e8 	:	val_out <= 4'ha570;
         4'h73e9 	:	val_out <= 4'ha570;
         4'h73ea 	:	val_out <= 4'ha570;
         4'h73eb 	:	val_out <= 4'ha570;
         4'h73f0 	:	val_out <= 4'ha558;
         4'h73f1 	:	val_out <= 4'ha558;
         4'h73f2 	:	val_out <= 4'ha558;
         4'h73f3 	:	val_out <= 4'ha558;
         4'h73f8 	:	val_out <= 4'ha540;
         4'h73f9 	:	val_out <= 4'ha540;
         4'h73fa 	:	val_out <= 4'ha540;
         4'h73fb 	:	val_out <= 4'ha540;
         4'h7400 	:	val_out <= 4'ha528;
         4'h7401 	:	val_out <= 4'ha528;
         4'h7402 	:	val_out <= 4'ha528;
         4'h7403 	:	val_out <= 4'ha528;
         4'h7408 	:	val_out <= 4'ha50f;
         4'h7409 	:	val_out <= 4'ha50f;
         4'h740a 	:	val_out <= 4'ha50f;
         4'h740b 	:	val_out <= 4'ha50f;
         4'h7410 	:	val_out <= 4'ha4f7;
         4'h7411 	:	val_out <= 4'ha4f7;
         4'h7412 	:	val_out <= 4'ha4f7;
         4'h7413 	:	val_out <= 4'ha4f7;
         4'h7418 	:	val_out <= 4'ha4df;
         4'h7419 	:	val_out <= 4'ha4df;
         4'h741a 	:	val_out <= 4'ha4df;
         4'h741b 	:	val_out <= 4'ha4df;
         4'h7420 	:	val_out <= 4'ha4c7;
         4'h7421 	:	val_out <= 4'ha4c7;
         4'h7422 	:	val_out <= 4'ha4c7;
         4'h7423 	:	val_out <= 4'ha4c7;
         4'h7428 	:	val_out <= 4'ha4af;
         4'h7429 	:	val_out <= 4'ha4af;
         4'h742a 	:	val_out <= 4'ha4af;
         4'h742b 	:	val_out <= 4'ha4af;
         4'h7430 	:	val_out <= 4'ha497;
         4'h7431 	:	val_out <= 4'ha497;
         4'h7432 	:	val_out <= 4'ha497;
         4'h7433 	:	val_out <= 4'ha497;
         4'h7438 	:	val_out <= 4'ha47f;
         4'h7439 	:	val_out <= 4'ha47f;
         4'h743a 	:	val_out <= 4'ha47f;
         4'h743b 	:	val_out <= 4'ha47f;
         4'h7440 	:	val_out <= 4'ha467;
         4'h7441 	:	val_out <= 4'ha467;
         4'h7442 	:	val_out <= 4'ha467;
         4'h7443 	:	val_out <= 4'ha467;
         4'h7448 	:	val_out <= 4'ha44f;
         4'h7449 	:	val_out <= 4'ha44f;
         4'h744a 	:	val_out <= 4'ha44f;
         4'h744b 	:	val_out <= 4'ha44f;
         4'h7450 	:	val_out <= 4'ha437;
         4'h7451 	:	val_out <= 4'ha437;
         4'h7452 	:	val_out <= 4'ha437;
         4'h7453 	:	val_out <= 4'ha437;
         4'h7458 	:	val_out <= 4'ha41f;
         4'h7459 	:	val_out <= 4'ha41f;
         4'h745a 	:	val_out <= 4'ha41f;
         4'h745b 	:	val_out <= 4'ha41f;
         4'h7460 	:	val_out <= 4'ha407;
         4'h7461 	:	val_out <= 4'ha407;
         4'h7462 	:	val_out <= 4'ha407;
         4'h7463 	:	val_out <= 4'ha407;
         4'h7468 	:	val_out <= 4'ha3ee;
         4'h7469 	:	val_out <= 4'ha3ee;
         4'h746a 	:	val_out <= 4'ha3ee;
         4'h746b 	:	val_out <= 4'ha3ee;
         4'h7470 	:	val_out <= 4'ha3d6;
         4'h7471 	:	val_out <= 4'ha3d6;
         4'h7472 	:	val_out <= 4'ha3d6;
         4'h7473 	:	val_out <= 4'ha3d6;
         4'h7478 	:	val_out <= 4'ha3be;
         4'h7479 	:	val_out <= 4'ha3be;
         4'h747a 	:	val_out <= 4'ha3be;
         4'h747b 	:	val_out <= 4'ha3be;
         4'h7480 	:	val_out <= 4'ha3a6;
         4'h7481 	:	val_out <= 4'ha3a6;
         4'h7482 	:	val_out <= 4'ha3a6;
         4'h7483 	:	val_out <= 4'ha3a6;
         4'h7488 	:	val_out <= 4'ha38e;
         4'h7489 	:	val_out <= 4'ha38e;
         4'h748a 	:	val_out <= 4'ha38e;
         4'h748b 	:	val_out <= 4'ha38e;
         4'h7490 	:	val_out <= 4'ha376;
         4'h7491 	:	val_out <= 4'ha376;
         4'h7492 	:	val_out <= 4'ha376;
         4'h7493 	:	val_out <= 4'ha376;
         4'h7498 	:	val_out <= 4'ha35e;
         4'h7499 	:	val_out <= 4'ha35e;
         4'h749a 	:	val_out <= 4'ha35e;
         4'h749b 	:	val_out <= 4'ha35e;
         4'h74a0 	:	val_out <= 4'ha345;
         4'h74a1 	:	val_out <= 4'ha345;
         4'h74a2 	:	val_out <= 4'ha345;
         4'h74a3 	:	val_out <= 4'ha345;
         4'h74a8 	:	val_out <= 4'ha32d;
         4'h74a9 	:	val_out <= 4'ha32d;
         4'h74aa 	:	val_out <= 4'ha32d;
         4'h74ab 	:	val_out <= 4'ha32d;
         4'h74b0 	:	val_out <= 4'ha315;
         4'h74b1 	:	val_out <= 4'ha315;
         4'h74b2 	:	val_out <= 4'ha315;
         4'h74b3 	:	val_out <= 4'ha315;
         4'h74b8 	:	val_out <= 4'ha2fd;
         4'h74b9 	:	val_out <= 4'ha2fd;
         4'h74ba 	:	val_out <= 4'ha2fd;
         4'h74bb 	:	val_out <= 4'ha2fd;
         4'h74c0 	:	val_out <= 4'ha2e5;
         4'h74c1 	:	val_out <= 4'ha2e5;
         4'h74c2 	:	val_out <= 4'ha2e5;
         4'h74c3 	:	val_out <= 4'ha2e5;
         4'h74c8 	:	val_out <= 4'ha2cd;
         4'h74c9 	:	val_out <= 4'ha2cd;
         4'h74ca 	:	val_out <= 4'ha2cd;
         4'h74cb 	:	val_out <= 4'ha2cd;
         4'h74d0 	:	val_out <= 4'ha2b4;
         4'h74d1 	:	val_out <= 4'ha2b4;
         4'h74d2 	:	val_out <= 4'ha2b4;
         4'h74d3 	:	val_out <= 4'ha2b4;
         4'h74d8 	:	val_out <= 4'ha29c;
         4'h74d9 	:	val_out <= 4'ha29c;
         4'h74da 	:	val_out <= 4'ha29c;
         4'h74db 	:	val_out <= 4'ha29c;
         4'h74e0 	:	val_out <= 4'ha284;
         4'h74e1 	:	val_out <= 4'ha284;
         4'h74e2 	:	val_out <= 4'ha284;
         4'h74e3 	:	val_out <= 4'ha284;
         4'h74e8 	:	val_out <= 4'ha26c;
         4'h74e9 	:	val_out <= 4'ha26c;
         4'h74ea 	:	val_out <= 4'ha26c;
         4'h74eb 	:	val_out <= 4'ha26c;
         4'h74f0 	:	val_out <= 4'ha254;
         4'h74f1 	:	val_out <= 4'ha254;
         4'h74f2 	:	val_out <= 4'ha254;
         4'h74f3 	:	val_out <= 4'ha254;
         4'h74f8 	:	val_out <= 4'ha23b;
         4'h74f9 	:	val_out <= 4'ha23b;
         4'h74fa 	:	val_out <= 4'ha23b;
         4'h74fb 	:	val_out <= 4'ha23b;
         4'h7500 	:	val_out <= 4'ha223;
         4'h7501 	:	val_out <= 4'ha223;
         4'h7502 	:	val_out <= 4'ha223;
         4'h7503 	:	val_out <= 4'ha223;
         4'h7508 	:	val_out <= 4'ha20b;
         4'h7509 	:	val_out <= 4'ha20b;
         4'h750a 	:	val_out <= 4'ha20b;
         4'h750b 	:	val_out <= 4'ha20b;
         4'h7510 	:	val_out <= 4'ha1f3;
         4'h7511 	:	val_out <= 4'ha1f3;
         4'h7512 	:	val_out <= 4'ha1f3;
         4'h7513 	:	val_out <= 4'ha1f3;
         4'h7518 	:	val_out <= 4'ha1da;
         4'h7519 	:	val_out <= 4'ha1da;
         4'h751a 	:	val_out <= 4'ha1da;
         4'h751b 	:	val_out <= 4'ha1da;
         4'h7520 	:	val_out <= 4'ha1c2;
         4'h7521 	:	val_out <= 4'ha1c2;
         4'h7522 	:	val_out <= 4'ha1c2;
         4'h7523 	:	val_out <= 4'ha1c2;
         4'h7528 	:	val_out <= 4'ha1aa;
         4'h7529 	:	val_out <= 4'ha1aa;
         4'h752a 	:	val_out <= 4'ha1aa;
         4'h752b 	:	val_out <= 4'ha1aa;
         4'h7530 	:	val_out <= 4'ha192;
         4'h7531 	:	val_out <= 4'ha192;
         4'h7532 	:	val_out <= 4'ha192;
         4'h7533 	:	val_out <= 4'ha192;
         4'h7538 	:	val_out <= 4'ha179;
         4'h7539 	:	val_out <= 4'ha179;
         4'h753a 	:	val_out <= 4'ha179;
         4'h753b 	:	val_out <= 4'ha179;
         4'h7540 	:	val_out <= 4'ha161;
         4'h7541 	:	val_out <= 4'ha161;
         4'h7542 	:	val_out <= 4'ha161;
         4'h7543 	:	val_out <= 4'ha161;
         4'h7548 	:	val_out <= 4'ha149;
         4'h7549 	:	val_out <= 4'ha149;
         4'h754a 	:	val_out <= 4'ha149;
         4'h754b 	:	val_out <= 4'ha149;
         4'h7550 	:	val_out <= 4'ha131;
         4'h7551 	:	val_out <= 4'ha131;
         4'h7552 	:	val_out <= 4'ha131;
         4'h7553 	:	val_out <= 4'ha131;
         4'h7558 	:	val_out <= 4'ha118;
         4'h7559 	:	val_out <= 4'ha118;
         4'h755a 	:	val_out <= 4'ha118;
         4'h755b 	:	val_out <= 4'ha118;
         4'h7560 	:	val_out <= 4'ha100;
         4'h7561 	:	val_out <= 4'ha100;
         4'h7562 	:	val_out <= 4'ha100;
         4'h7563 	:	val_out <= 4'ha100;
         4'h7568 	:	val_out <= 4'ha0e8;
         4'h7569 	:	val_out <= 4'ha0e8;
         4'h756a 	:	val_out <= 4'ha0e8;
         4'h756b 	:	val_out <= 4'ha0e8;
         4'h7570 	:	val_out <= 4'ha0d0;
         4'h7571 	:	val_out <= 4'ha0d0;
         4'h7572 	:	val_out <= 4'ha0d0;
         4'h7573 	:	val_out <= 4'ha0d0;
         4'h7578 	:	val_out <= 4'ha0b7;
         4'h7579 	:	val_out <= 4'ha0b7;
         4'h757a 	:	val_out <= 4'ha0b7;
         4'h757b 	:	val_out <= 4'ha0b7;
         4'h7580 	:	val_out <= 4'ha09f;
         4'h7581 	:	val_out <= 4'ha09f;
         4'h7582 	:	val_out <= 4'ha09f;
         4'h7583 	:	val_out <= 4'ha09f;
         4'h7588 	:	val_out <= 4'ha087;
         4'h7589 	:	val_out <= 4'ha087;
         4'h758a 	:	val_out <= 4'ha087;
         4'h758b 	:	val_out <= 4'ha087;
         4'h7590 	:	val_out <= 4'ha06e;
         4'h7591 	:	val_out <= 4'ha06e;
         4'h7592 	:	val_out <= 4'ha06e;
         4'h7593 	:	val_out <= 4'ha06e;
         4'h7598 	:	val_out <= 4'ha056;
         4'h7599 	:	val_out <= 4'ha056;
         4'h759a 	:	val_out <= 4'ha056;
         4'h759b 	:	val_out <= 4'ha056;
         4'h75a0 	:	val_out <= 4'ha03e;
         4'h75a1 	:	val_out <= 4'ha03e;
         4'h75a2 	:	val_out <= 4'ha03e;
         4'h75a3 	:	val_out <= 4'ha03e;
         4'h75a8 	:	val_out <= 4'ha025;
         4'h75a9 	:	val_out <= 4'ha025;
         4'h75aa 	:	val_out <= 4'ha025;
         4'h75ab 	:	val_out <= 4'ha025;
         4'h75b0 	:	val_out <= 4'ha00d;
         4'h75b1 	:	val_out <= 4'ha00d;
         4'h75b2 	:	val_out <= 4'ha00d;
         4'h75b3 	:	val_out <= 4'ha00d;
         4'h75b8 	:	val_out <= 4'h9ff5;
         4'h75b9 	:	val_out <= 4'h9ff5;
         4'h75ba 	:	val_out <= 4'h9ff5;
         4'h75bb 	:	val_out <= 4'h9ff5;
         4'h75c0 	:	val_out <= 4'h9fdc;
         4'h75c1 	:	val_out <= 4'h9fdc;
         4'h75c2 	:	val_out <= 4'h9fdc;
         4'h75c3 	:	val_out <= 4'h9fdc;
         4'h75c8 	:	val_out <= 4'h9fc4;
         4'h75c9 	:	val_out <= 4'h9fc4;
         4'h75ca 	:	val_out <= 4'h9fc4;
         4'h75cb 	:	val_out <= 4'h9fc4;
         4'h75d0 	:	val_out <= 4'h9fac;
         4'h75d1 	:	val_out <= 4'h9fac;
         4'h75d2 	:	val_out <= 4'h9fac;
         4'h75d3 	:	val_out <= 4'h9fac;
         4'h75d8 	:	val_out <= 4'h9f93;
         4'h75d9 	:	val_out <= 4'h9f93;
         4'h75da 	:	val_out <= 4'h9f93;
         4'h75db 	:	val_out <= 4'h9f93;
         4'h75e0 	:	val_out <= 4'h9f7b;
         4'h75e1 	:	val_out <= 4'h9f7b;
         4'h75e2 	:	val_out <= 4'h9f7b;
         4'h75e3 	:	val_out <= 4'h9f7b;
         4'h75e8 	:	val_out <= 4'h9f63;
         4'h75e9 	:	val_out <= 4'h9f63;
         4'h75ea 	:	val_out <= 4'h9f63;
         4'h75eb 	:	val_out <= 4'h9f63;
         4'h75f0 	:	val_out <= 4'h9f4a;
         4'h75f1 	:	val_out <= 4'h9f4a;
         4'h75f2 	:	val_out <= 4'h9f4a;
         4'h75f3 	:	val_out <= 4'h9f4a;
         4'h75f8 	:	val_out <= 4'h9f32;
         4'h75f9 	:	val_out <= 4'h9f32;
         4'h75fa 	:	val_out <= 4'h9f32;
         4'h75fb 	:	val_out <= 4'h9f32;
         4'h7600 	:	val_out <= 4'h9f19;
         4'h7601 	:	val_out <= 4'h9f19;
         4'h7602 	:	val_out <= 4'h9f19;
         4'h7603 	:	val_out <= 4'h9f19;
         4'h7608 	:	val_out <= 4'h9f01;
         4'h7609 	:	val_out <= 4'h9f01;
         4'h760a 	:	val_out <= 4'h9f01;
         4'h760b 	:	val_out <= 4'h9f01;
         4'h7610 	:	val_out <= 4'h9ee9;
         4'h7611 	:	val_out <= 4'h9ee9;
         4'h7612 	:	val_out <= 4'h9ee9;
         4'h7613 	:	val_out <= 4'h9ee9;
         4'h7618 	:	val_out <= 4'h9ed0;
         4'h7619 	:	val_out <= 4'h9ed0;
         4'h761a 	:	val_out <= 4'h9ed0;
         4'h761b 	:	val_out <= 4'h9ed0;
         4'h7620 	:	val_out <= 4'h9eb8;
         4'h7621 	:	val_out <= 4'h9eb8;
         4'h7622 	:	val_out <= 4'h9eb8;
         4'h7623 	:	val_out <= 4'h9eb8;
         4'h7628 	:	val_out <= 4'h9ea0;
         4'h7629 	:	val_out <= 4'h9ea0;
         4'h762a 	:	val_out <= 4'h9ea0;
         4'h762b 	:	val_out <= 4'h9ea0;
         4'h7630 	:	val_out <= 4'h9e87;
         4'h7631 	:	val_out <= 4'h9e87;
         4'h7632 	:	val_out <= 4'h9e87;
         4'h7633 	:	val_out <= 4'h9e87;
         4'h7638 	:	val_out <= 4'h9e6f;
         4'h7639 	:	val_out <= 4'h9e6f;
         4'h763a 	:	val_out <= 4'h9e6f;
         4'h763b 	:	val_out <= 4'h9e6f;
         4'h7640 	:	val_out <= 4'h9e56;
         4'h7641 	:	val_out <= 4'h9e56;
         4'h7642 	:	val_out <= 4'h9e56;
         4'h7643 	:	val_out <= 4'h9e56;
         4'h7648 	:	val_out <= 4'h9e3e;
         4'h7649 	:	val_out <= 4'h9e3e;
         4'h764a 	:	val_out <= 4'h9e3e;
         4'h764b 	:	val_out <= 4'h9e3e;
         4'h7650 	:	val_out <= 4'h9e25;
         4'h7651 	:	val_out <= 4'h9e25;
         4'h7652 	:	val_out <= 4'h9e25;
         4'h7653 	:	val_out <= 4'h9e25;
         4'h7658 	:	val_out <= 4'h9e0d;
         4'h7659 	:	val_out <= 4'h9e0d;
         4'h765a 	:	val_out <= 4'h9e0d;
         4'h765b 	:	val_out <= 4'h9e0d;
         4'h7660 	:	val_out <= 4'h9df5;
         4'h7661 	:	val_out <= 4'h9df5;
         4'h7662 	:	val_out <= 4'h9df5;
         4'h7663 	:	val_out <= 4'h9df5;
         4'h7668 	:	val_out <= 4'h9ddc;
         4'h7669 	:	val_out <= 4'h9ddc;
         4'h766a 	:	val_out <= 4'h9ddc;
         4'h766b 	:	val_out <= 4'h9ddc;
         4'h7670 	:	val_out <= 4'h9dc4;
         4'h7671 	:	val_out <= 4'h9dc4;
         4'h7672 	:	val_out <= 4'h9dc4;
         4'h7673 	:	val_out <= 4'h9dc4;
         4'h7678 	:	val_out <= 4'h9dab;
         4'h7679 	:	val_out <= 4'h9dab;
         4'h767a 	:	val_out <= 4'h9dab;
         4'h767b 	:	val_out <= 4'h9dab;
         4'h7680 	:	val_out <= 4'h9d93;
         4'h7681 	:	val_out <= 4'h9d93;
         4'h7682 	:	val_out <= 4'h9d93;
         4'h7683 	:	val_out <= 4'h9d93;
         4'h7688 	:	val_out <= 4'h9d7a;
         4'h7689 	:	val_out <= 4'h9d7a;
         4'h768a 	:	val_out <= 4'h9d7a;
         4'h768b 	:	val_out <= 4'h9d7a;
         4'h7690 	:	val_out <= 4'h9d62;
         4'h7691 	:	val_out <= 4'h9d62;
         4'h7692 	:	val_out <= 4'h9d62;
         4'h7693 	:	val_out <= 4'h9d62;
         4'h7698 	:	val_out <= 4'h9d49;
         4'h7699 	:	val_out <= 4'h9d49;
         4'h769a 	:	val_out <= 4'h9d49;
         4'h769b 	:	val_out <= 4'h9d49;
         4'h76a0 	:	val_out <= 4'h9d31;
         4'h76a1 	:	val_out <= 4'h9d31;
         4'h76a2 	:	val_out <= 4'h9d31;
         4'h76a3 	:	val_out <= 4'h9d31;
         4'h76a8 	:	val_out <= 4'h9d18;
         4'h76a9 	:	val_out <= 4'h9d18;
         4'h76aa 	:	val_out <= 4'h9d18;
         4'h76ab 	:	val_out <= 4'h9d18;
         4'h76b0 	:	val_out <= 4'h9d00;
         4'h76b1 	:	val_out <= 4'h9d00;
         4'h76b2 	:	val_out <= 4'h9d00;
         4'h76b3 	:	val_out <= 4'h9d00;
         4'h76b8 	:	val_out <= 4'h9ce8;
         4'h76b9 	:	val_out <= 4'h9ce8;
         4'h76ba 	:	val_out <= 4'h9ce8;
         4'h76bb 	:	val_out <= 4'h9ce8;
         4'h76c0 	:	val_out <= 4'h9ccf;
         4'h76c1 	:	val_out <= 4'h9ccf;
         4'h76c2 	:	val_out <= 4'h9ccf;
         4'h76c3 	:	val_out <= 4'h9ccf;
         4'h76c8 	:	val_out <= 4'h9cb7;
         4'h76c9 	:	val_out <= 4'h9cb7;
         4'h76ca 	:	val_out <= 4'h9cb7;
         4'h76cb 	:	val_out <= 4'h9cb7;
         4'h76d0 	:	val_out <= 4'h9c9e;
         4'h76d1 	:	val_out <= 4'h9c9e;
         4'h76d2 	:	val_out <= 4'h9c9e;
         4'h76d3 	:	val_out <= 4'h9c9e;
         4'h76d8 	:	val_out <= 4'h9c86;
         4'h76d9 	:	val_out <= 4'h9c86;
         4'h76da 	:	val_out <= 4'h9c86;
         4'h76db 	:	val_out <= 4'h9c86;
         4'h76e0 	:	val_out <= 4'h9c6d;
         4'h76e1 	:	val_out <= 4'h9c6d;
         4'h76e2 	:	val_out <= 4'h9c6d;
         4'h76e3 	:	val_out <= 4'h9c6d;
         4'h76e8 	:	val_out <= 4'h9c55;
         4'h76e9 	:	val_out <= 4'h9c55;
         4'h76ea 	:	val_out <= 4'h9c55;
         4'h76eb 	:	val_out <= 4'h9c55;
         4'h76f0 	:	val_out <= 4'h9c3c;
         4'h76f1 	:	val_out <= 4'h9c3c;
         4'h76f2 	:	val_out <= 4'h9c3c;
         4'h76f3 	:	val_out <= 4'h9c3c;
         4'h76f8 	:	val_out <= 4'h9c24;
         4'h76f9 	:	val_out <= 4'h9c24;
         4'h76fa 	:	val_out <= 4'h9c24;
         4'h76fb 	:	val_out <= 4'h9c24;
         4'h7700 	:	val_out <= 4'h9c0b;
         4'h7701 	:	val_out <= 4'h9c0b;
         4'h7702 	:	val_out <= 4'h9c0b;
         4'h7703 	:	val_out <= 4'h9c0b;
         4'h7708 	:	val_out <= 4'h9bf2;
         4'h7709 	:	val_out <= 4'h9bf2;
         4'h770a 	:	val_out <= 4'h9bf2;
         4'h770b 	:	val_out <= 4'h9bf2;
         4'h7710 	:	val_out <= 4'h9bda;
         4'h7711 	:	val_out <= 4'h9bda;
         4'h7712 	:	val_out <= 4'h9bda;
         4'h7713 	:	val_out <= 4'h9bda;
         4'h7718 	:	val_out <= 4'h9bc1;
         4'h7719 	:	val_out <= 4'h9bc1;
         4'h771a 	:	val_out <= 4'h9bc1;
         4'h771b 	:	val_out <= 4'h9bc1;
         4'h7720 	:	val_out <= 4'h9ba9;
         4'h7721 	:	val_out <= 4'h9ba9;
         4'h7722 	:	val_out <= 4'h9ba9;
         4'h7723 	:	val_out <= 4'h9ba9;
         4'h7728 	:	val_out <= 4'h9b90;
         4'h7729 	:	val_out <= 4'h9b90;
         4'h772a 	:	val_out <= 4'h9b90;
         4'h772b 	:	val_out <= 4'h9b90;
         4'h7730 	:	val_out <= 4'h9b78;
         4'h7731 	:	val_out <= 4'h9b78;
         4'h7732 	:	val_out <= 4'h9b78;
         4'h7733 	:	val_out <= 4'h9b78;
         4'h7738 	:	val_out <= 4'h9b5f;
         4'h7739 	:	val_out <= 4'h9b5f;
         4'h773a 	:	val_out <= 4'h9b5f;
         4'h773b 	:	val_out <= 4'h9b5f;
         4'h7740 	:	val_out <= 4'h9b47;
         4'h7741 	:	val_out <= 4'h9b47;
         4'h7742 	:	val_out <= 4'h9b47;
         4'h7743 	:	val_out <= 4'h9b47;
         4'h7748 	:	val_out <= 4'h9b2e;
         4'h7749 	:	val_out <= 4'h9b2e;
         4'h774a 	:	val_out <= 4'h9b2e;
         4'h774b 	:	val_out <= 4'h9b2e;
         4'h7750 	:	val_out <= 4'h9b16;
         4'h7751 	:	val_out <= 4'h9b16;
         4'h7752 	:	val_out <= 4'h9b16;
         4'h7753 	:	val_out <= 4'h9b16;
         4'h7758 	:	val_out <= 4'h9afd;
         4'h7759 	:	val_out <= 4'h9afd;
         4'h775a 	:	val_out <= 4'h9afd;
         4'h775b 	:	val_out <= 4'h9afd;
         4'h7760 	:	val_out <= 4'h9ae4;
         4'h7761 	:	val_out <= 4'h9ae4;
         4'h7762 	:	val_out <= 4'h9ae4;
         4'h7763 	:	val_out <= 4'h9ae4;
         4'h7768 	:	val_out <= 4'h9acc;
         4'h7769 	:	val_out <= 4'h9acc;
         4'h776a 	:	val_out <= 4'h9acc;
         4'h776b 	:	val_out <= 4'h9acc;
         4'h7770 	:	val_out <= 4'h9ab3;
         4'h7771 	:	val_out <= 4'h9ab3;
         4'h7772 	:	val_out <= 4'h9ab3;
         4'h7773 	:	val_out <= 4'h9ab3;
         4'h7778 	:	val_out <= 4'h9a9b;
         4'h7779 	:	val_out <= 4'h9a9b;
         4'h777a 	:	val_out <= 4'h9a9b;
         4'h777b 	:	val_out <= 4'h9a9b;
         4'h7780 	:	val_out <= 4'h9a82;
         4'h7781 	:	val_out <= 4'h9a82;
         4'h7782 	:	val_out <= 4'h9a82;
         4'h7783 	:	val_out <= 4'h9a82;
         4'h7788 	:	val_out <= 4'h9a6a;
         4'h7789 	:	val_out <= 4'h9a6a;
         4'h778a 	:	val_out <= 4'h9a6a;
         4'h778b 	:	val_out <= 4'h9a6a;
         4'h7790 	:	val_out <= 4'h9a51;
         4'h7791 	:	val_out <= 4'h9a51;
         4'h7792 	:	val_out <= 4'h9a51;
         4'h7793 	:	val_out <= 4'h9a51;
         4'h7798 	:	val_out <= 4'h9a38;
         4'h7799 	:	val_out <= 4'h9a38;
         4'h779a 	:	val_out <= 4'h9a38;
         4'h779b 	:	val_out <= 4'h9a38;
         4'h77a0 	:	val_out <= 4'h9a20;
         4'h77a1 	:	val_out <= 4'h9a20;
         4'h77a2 	:	val_out <= 4'h9a20;
         4'h77a3 	:	val_out <= 4'h9a20;
         4'h77a8 	:	val_out <= 4'h9a07;
         4'h77a9 	:	val_out <= 4'h9a07;
         4'h77aa 	:	val_out <= 4'h9a07;
         4'h77ab 	:	val_out <= 4'h9a07;
         4'h77b0 	:	val_out <= 4'h99ef;
         4'h77b1 	:	val_out <= 4'h99ef;
         4'h77b2 	:	val_out <= 4'h99ef;
         4'h77b3 	:	val_out <= 4'h99ef;
         4'h77b8 	:	val_out <= 4'h99d6;
         4'h77b9 	:	val_out <= 4'h99d6;
         4'h77ba 	:	val_out <= 4'h99d6;
         4'h77bb 	:	val_out <= 4'h99d6;
         4'h77c0 	:	val_out <= 4'h99bd;
         4'h77c1 	:	val_out <= 4'h99bd;
         4'h77c2 	:	val_out <= 4'h99bd;
         4'h77c3 	:	val_out <= 4'h99bd;
         4'h77c8 	:	val_out <= 4'h99a5;
         4'h77c9 	:	val_out <= 4'h99a5;
         4'h77ca 	:	val_out <= 4'h99a5;
         4'h77cb 	:	val_out <= 4'h99a5;
         4'h77d0 	:	val_out <= 4'h998c;
         4'h77d1 	:	val_out <= 4'h998c;
         4'h77d2 	:	val_out <= 4'h998c;
         4'h77d3 	:	val_out <= 4'h998c;
         4'h77d8 	:	val_out <= 4'h9973;
         4'h77d9 	:	val_out <= 4'h9973;
         4'h77da 	:	val_out <= 4'h9973;
         4'h77db 	:	val_out <= 4'h9973;
         4'h77e0 	:	val_out <= 4'h995b;
         4'h77e1 	:	val_out <= 4'h995b;
         4'h77e2 	:	val_out <= 4'h995b;
         4'h77e3 	:	val_out <= 4'h995b;
         4'h77e8 	:	val_out <= 4'h9942;
         4'h77e9 	:	val_out <= 4'h9942;
         4'h77ea 	:	val_out <= 4'h9942;
         4'h77eb 	:	val_out <= 4'h9942;
         4'h77f0 	:	val_out <= 4'h992a;
         4'h77f1 	:	val_out <= 4'h992a;
         4'h77f2 	:	val_out <= 4'h992a;
         4'h77f3 	:	val_out <= 4'h992a;
         4'h77f8 	:	val_out <= 4'h9911;
         4'h77f9 	:	val_out <= 4'h9911;
         4'h77fa 	:	val_out <= 4'h9911;
         4'h77fb 	:	val_out <= 4'h9911;
         4'h7800 	:	val_out <= 4'h98f8;
         4'h7801 	:	val_out <= 4'h98f8;
         4'h7802 	:	val_out <= 4'h98f8;
         4'h7803 	:	val_out <= 4'h98f8;
         4'h7808 	:	val_out <= 4'h98e0;
         4'h7809 	:	val_out <= 4'h98e0;
         4'h780a 	:	val_out <= 4'h98e0;
         4'h780b 	:	val_out <= 4'h98e0;
         4'h7810 	:	val_out <= 4'h98c7;
         4'h7811 	:	val_out <= 4'h98c7;
         4'h7812 	:	val_out <= 4'h98c7;
         4'h7813 	:	val_out <= 4'h98c7;
         4'h7818 	:	val_out <= 4'h98ae;
         4'h7819 	:	val_out <= 4'h98ae;
         4'h781a 	:	val_out <= 4'h98ae;
         4'h781b 	:	val_out <= 4'h98ae;
         4'h7820 	:	val_out <= 4'h9896;
         4'h7821 	:	val_out <= 4'h9896;
         4'h7822 	:	val_out <= 4'h9896;
         4'h7823 	:	val_out <= 4'h9896;
         4'h7828 	:	val_out <= 4'h987d;
         4'h7829 	:	val_out <= 4'h987d;
         4'h782a 	:	val_out <= 4'h987d;
         4'h782b 	:	val_out <= 4'h987d;
         4'h7830 	:	val_out <= 4'h9864;
         4'h7831 	:	val_out <= 4'h9864;
         4'h7832 	:	val_out <= 4'h9864;
         4'h7833 	:	val_out <= 4'h9864;
         4'h7838 	:	val_out <= 4'h984c;
         4'h7839 	:	val_out <= 4'h984c;
         4'h783a 	:	val_out <= 4'h984c;
         4'h783b 	:	val_out <= 4'h984c;
         4'h7840 	:	val_out <= 4'h9833;
         4'h7841 	:	val_out <= 4'h9833;
         4'h7842 	:	val_out <= 4'h9833;
         4'h7843 	:	val_out <= 4'h9833;
         4'h7848 	:	val_out <= 4'h981a;
         4'h7849 	:	val_out <= 4'h981a;
         4'h784a 	:	val_out <= 4'h981a;
         4'h784b 	:	val_out <= 4'h981a;
         4'h7850 	:	val_out <= 4'h9802;
         4'h7851 	:	val_out <= 4'h9802;
         4'h7852 	:	val_out <= 4'h9802;
         4'h7853 	:	val_out <= 4'h9802;
         4'h7858 	:	val_out <= 4'h97e9;
         4'h7859 	:	val_out <= 4'h97e9;
         4'h785a 	:	val_out <= 4'h97e9;
         4'h785b 	:	val_out <= 4'h97e9;
         4'h7860 	:	val_out <= 4'h97d0;
         4'h7861 	:	val_out <= 4'h97d0;
         4'h7862 	:	val_out <= 4'h97d0;
         4'h7863 	:	val_out <= 4'h97d0;
         4'h7868 	:	val_out <= 4'h97b7;
         4'h7869 	:	val_out <= 4'h97b7;
         4'h786a 	:	val_out <= 4'h97b7;
         4'h786b 	:	val_out <= 4'h97b7;
         4'h7870 	:	val_out <= 4'h979f;
         4'h7871 	:	val_out <= 4'h979f;
         4'h7872 	:	val_out <= 4'h979f;
         4'h7873 	:	val_out <= 4'h979f;
         4'h7878 	:	val_out <= 4'h9786;
         4'h7879 	:	val_out <= 4'h9786;
         4'h787a 	:	val_out <= 4'h9786;
         4'h787b 	:	val_out <= 4'h9786;
         4'h7880 	:	val_out <= 4'h976d;
         4'h7881 	:	val_out <= 4'h976d;
         4'h7882 	:	val_out <= 4'h976d;
         4'h7883 	:	val_out <= 4'h976d;
         4'h7888 	:	val_out <= 4'h9755;
         4'h7889 	:	val_out <= 4'h9755;
         4'h788a 	:	val_out <= 4'h9755;
         4'h788b 	:	val_out <= 4'h9755;
         4'h7890 	:	val_out <= 4'h973c;
         4'h7891 	:	val_out <= 4'h973c;
         4'h7892 	:	val_out <= 4'h973c;
         4'h7893 	:	val_out <= 4'h973c;
         4'h7898 	:	val_out <= 4'h9723;
         4'h7899 	:	val_out <= 4'h9723;
         4'h789a 	:	val_out <= 4'h9723;
         4'h789b 	:	val_out <= 4'h9723;
         4'h78a0 	:	val_out <= 4'h970a;
         4'h78a1 	:	val_out <= 4'h970a;
         4'h78a2 	:	val_out <= 4'h970a;
         4'h78a3 	:	val_out <= 4'h970a;
         4'h78a8 	:	val_out <= 4'h96f2;
         4'h78a9 	:	val_out <= 4'h96f2;
         4'h78aa 	:	val_out <= 4'h96f2;
         4'h78ab 	:	val_out <= 4'h96f2;
         4'h78b0 	:	val_out <= 4'h96d9;
         4'h78b1 	:	val_out <= 4'h96d9;
         4'h78b2 	:	val_out <= 4'h96d9;
         4'h78b3 	:	val_out <= 4'h96d9;
         4'h78b8 	:	val_out <= 4'h96c0;
         4'h78b9 	:	val_out <= 4'h96c0;
         4'h78ba 	:	val_out <= 4'h96c0;
         4'h78bb 	:	val_out <= 4'h96c0;
         4'h78c0 	:	val_out <= 4'h96a8;
         4'h78c1 	:	val_out <= 4'h96a8;
         4'h78c2 	:	val_out <= 4'h96a8;
         4'h78c3 	:	val_out <= 4'h96a8;
         4'h78c8 	:	val_out <= 4'h968f;
         4'h78c9 	:	val_out <= 4'h968f;
         4'h78ca 	:	val_out <= 4'h968f;
         4'h78cb 	:	val_out <= 4'h968f;
         4'h78d0 	:	val_out <= 4'h9676;
         4'h78d1 	:	val_out <= 4'h9676;
         4'h78d2 	:	val_out <= 4'h9676;
         4'h78d3 	:	val_out <= 4'h9676;
         4'h78d8 	:	val_out <= 4'h965d;
         4'h78d9 	:	val_out <= 4'h965d;
         4'h78da 	:	val_out <= 4'h965d;
         4'h78db 	:	val_out <= 4'h965d;
         4'h78e0 	:	val_out <= 4'h9645;
         4'h78e1 	:	val_out <= 4'h9645;
         4'h78e2 	:	val_out <= 4'h9645;
         4'h78e3 	:	val_out <= 4'h9645;
         4'h78e8 	:	val_out <= 4'h962c;
         4'h78e9 	:	val_out <= 4'h962c;
         4'h78ea 	:	val_out <= 4'h962c;
         4'h78eb 	:	val_out <= 4'h962c;
         4'h78f0 	:	val_out <= 4'h9613;
         4'h78f1 	:	val_out <= 4'h9613;
         4'h78f2 	:	val_out <= 4'h9613;
         4'h78f3 	:	val_out <= 4'h9613;
         4'h78f8 	:	val_out <= 4'h95fa;
         4'h78f9 	:	val_out <= 4'h95fa;
         4'h78fa 	:	val_out <= 4'h95fa;
         4'h78fb 	:	val_out <= 4'h95fa;
         4'h7900 	:	val_out <= 4'h95e2;
         4'h7901 	:	val_out <= 4'h95e2;
         4'h7902 	:	val_out <= 4'h95e2;
         4'h7903 	:	val_out <= 4'h95e2;
         4'h7908 	:	val_out <= 4'h95c9;
         4'h7909 	:	val_out <= 4'h95c9;
         4'h790a 	:	val_out <= 4'h95c9;
         4'h790b 	:	val_out <= 4'h95c9;
         4'h7910 	:	val_out <= 4'h95b0;
         4'h7911 	:	val_out <= 4'h95b0;
         4'h7912 	:	val_out <= 4'h95b0;
         4'h7913 	:	val_out <= 4'h95b0;
         4'h7918 	:	val_out <= 4'h9597;
         4'h7919 	:	val_out <= 4'h9597;
         4'h791a 	:	val_out <= 4'h9597;
         4'h791b 	:	val_out <= 4'h9597;
         4'h7920 	:	val_out <= 4'h957f;
         4'h7921 	:	val_out <= 4'h957f;
         4'h7922 	:	val_out <= 4'h957f;
         4'h7923 	:	val_out <= 4'h957f;
         4'h7928 	:	val_out <= 4'h9566;
         4'h7929 	:	val_out <= 4'h9566;
         4'h792a 	:	val_out <= 4'h9566;
         4'h792b 	:	val_out <= 4'h9566;
         4'h7930 	:	val_out <= 4'h954d;
         4'h7931 	:	val_out <= 4'h954d;
         4'h7932 	:	val_out <= 4'h954d;
         4'h7933 	:	val_out <= 4'h954d;
         4'h7938 	:	val_out <= 4'h9534;
         4'h7939 	:	val_out <= 4'h9534;
         4'h793a 	:	val_out <= 4'h9534;
         4'h793b 	:	val_out <= 4'h9534;
         4'h7940 	:	val_out <= 4'h951b;
         4'h7941 	:	val_out <= 4'h951b;
         4'h7942 	:	val_out <= 4'h951b;
         4'h7943 	:	val_out <= 4'h951b;
         4'h7948 	:	val_out <= 4'h9503;
         4'h7949 	:	val_out <= 4'h9503;
         4'h794a 	:	val_out <= 4'h9503;
         4'h794b 	:	val_out <= 4'h9503;
         4'h7950 	:	val_out <= 4'h94ea;
         4'h7951 	:	val_out <= 4'h94ea;
         4'h7952 	:	val_out <= 4'h94ea;
         4'h7953 	:	val_out <= 4'h94ea;
         4'h7958 	:	val_out <= 4'h94d1;
         4'h7959 	:	val_out <= 4'h94d1;
         4'h795a 	:	val_out <= 4'h94d1;
         4'h795b 	:	val_out <= 4'h94d1;
         4'h7960 	:	val_out <= 4'h94b8;
         4'h7961 	:	val_out <= 4'h94b8;
         4'h7962 	:	val_out <= 4'h94b8;
         4'h7963 	:	val_out <= 4'h94b8;
         4'h7968 	:	val_out <= 4'h949f;
         4'h7969 	:	val_out <= 4'h949f;
         4'h796a 	:	val_out <= 4'h949f;
         4'h796b 	:	val_out <= 4'h949f;
         4'h7970 	:	val_out <= 4'h9487;
         4'h7971 	:	val_out <= 4'h9487;
         4'h7972 	:	val_out <= 4'h9487;
         4'h7973 	:	val_out <= 4'h9487;
         4'h7978 	:	val_out <= 4'h946e;
         4'h7979 	:	val_out <= 4'h946e;
         4'h797a 	:	val_out <= 4'h946e;
         4'h797b 	:	val_out <= 4'h946e;
         4'h7980 	:	val_out <= 4'h9455;
         4'h7981 	:	val_out <= 4'h9455;
         4'h7982 	:	val_out <= 4'h9455;
         4'h7983 	:	val_out <= 4'h9455;
         4'h7988 	:	val_out <= 4'h943c;
         4'h7989 	:	val_out <= 4'h943c;
         4'h798a 	:	val_out <= 4'h943c;
         4'h798b 	:	val_out <= 4'h943c;
         4'h7990 	:	val_out <= 4'h9423;
         4'h7991 	:	val_out <= 4'h9423;
         4'h7992 	:	val_out <= 4'h9423;
         4'h7993 	:	val_out <= 4'h9423;
         4'h7998 	:	val_out <= 4'h940b;
         4'h7999 	:	val_out <= 4'h940b;
         4'h799a 	:	val_out <= 4'h940b;
         4'h799b 	:	val_out <= 4'h940b;
         4'h79a0 	:	val_out <= 4'h93f2;
         4'h79a1 	:	val_out <= 4'h93f2;
         4'h79a2 	:	val_out <= 4'h93f2;
         4'h79a3 	:	val_out <= 4'h93f2;
         4'h79a8 	:	val_out <= 4'h93d9;
         4'h79a9 	:	val_out <= 4'h93d9;
         4'h79aa 	:	val_out <= 4'h93d9;
         4'h79ab 	:	val_out <= 4'h93d9;
         4'h79b0 	:	val_out <= 4'h93c0;
         4'h79b1 	:	val_out <= 4'h93c0;
         4'h79b2 	:	val_out <= 4'h93c0;
         4'h79b3 	:	val_out <= 4'h93c0;
         4'h79b8 	:	val_out <= 4'h93a7;
         4'h79b9 	:	val_out <= 4'h93a7;
         4'h79ba 	:	val_out <= 4'h93a7;
         4'h79bb 	:	val_out <= 4'h93a7;
         4'h79c0 	:	val_out <= 4'h938e;
         4'h79c1 	:	val_out <= 4'h938e;
         4'h79c2 	:	val_out <= 4'h938e;
         4'h79c3 	:	val_out <= 4'h938e;
         4'h79c8 	:	val_out <= 4'h9376;
         4'h79c9 	:	val_out <= 4'h9376;
         4'h79ca 	:	val_out <= 4'h9376;
         4'h79cb 	:	val_out <= 4'h9376;
         4'h79d0 	:	val_out <= 4'h935d;
         4'h79d1 	:	val_out <= 4'h935d;
         4'h79d2 	:	val_out <= 4'h935d;
         4'h79d3 	:	val_out <= 4'h935d;
         4'h79d8 	:	val_out <= 4'h9344;
         4'h79d9 	:	val_out <= 4'h9344;
         4'h79da 	:	val_out <= 4'h9344;
         4'h79db 	:	val_out <= 4'h9344;
         4'h79e0 	:	val_out <= 4'h932b;
         4'h79e1 	:	val_out <= 4'h932b;
         4'h79e2 	:	val_out <= 4'h932b;
         4'h79e3 	:	val_out <= 4'h932b;
         4'h79e8 	:	val_out <= 4'h9312;
         4'h79e9 	:	val_out <= 4'h9312;
         4'h79ea 	:	val_out <= 4'h9312;
         4'h79eb 	:	val_out <= 4'h9312;
         4'h79f0 	:	val_out <= 4'h92f9;
         4'h79f1 	:	val_out <= 4'h92f9;
         4'h79f2 	:	val_out <= 4'h92f9;
         4'h79f3 	:	val_out <= 4'h92f9;
         4'h79f8 	:	val_out <= 4'h92e0;
         4'h79f9 	:	val_out <= 4'h92e0;
         4'h79fa 	:	val_out <= 4'h92e0;
         4'h79fb 	:	val_out <= 4'h92e0;
         4'h7a00 	:	val_out <= 4'h92c8;
         4'h7a01 	:	val_out <= 4'h92c8;
         4'h7a02 	:	val_out <= 4'h92c8;
         4'h7a03 	:	val_out <= 4'h92c8;
         4'h7a08 	:	val_out <= 4'h92af;
         4'h7a09 	:	val_out <= 4'h92af;
         4'h7a0a 	:	val_out <= 4'h92af;
         4'h7a0b 	:	val_out <= 4'h92af;
         4'h7a10 	:	val_out <= 4'h9296;
         4'h7a11 	:	val_out <= 4'h9296;
         4'h7a12 	:	val_out <= 4'h9296;
         4'h7a13 	:	val_out <= 4'h9296;
         4'h7a18 	:	val_out <= 4'h927d;
         4'h7a19 	:	val_out <= 4'h927d;
         4'h7a1a 	:	val_out <= 4'h927d;
         4'h7a1b 	:	val_out <= 4'h927d;
         4'h7a20 	:	val_out <= 4'h9264;
         4'h7a21 	:	val_out <= 4'h9264;
         4'h7a22 	:	val_out <= 4'h9264;
         4'h7a23 	:	val_out <= 4'h9264;
         4'h7a28 	:	val_out <= 4'h924b;
         4'h7a29 	:	val_out <= 4'h924b;
         4'h7a2a 	:	val_out <= 4'h924b;
         4'h7a2b 	:	val_out <= 4'h924b;
         4'h7a30 	:	val_out <= 4'h9232;
         4'h7a31 	:	val_out <= 4'h9232;
         4'h7a32 	:	val_out <= 4'h9232;
         4'h7a33 	:	val_out <= 4'h9232;
         4'h7a38 	:	val_out <= 4'h9219;
         4'h7a39 	:	val_out <= 4'h9219;
         4'h7a3a 	:	val_out <= 4'h9219;
         4'h7a3b 	:	val_out <= 4'h9219;
         4'h7a40 	:	val_out <= 4'h9201;
         4'h7a41 	:	val_out <= 4'h9201;
         4'h7a42 	:	val_out <= 4'h9201;
         4'h7a43 	:	val_out <= 4'h9201;
         4'h7a48 	:	val_out <= 4'h91e8;
         4'h7a49 	:	val_out <= 4'h91e8;
         4'h7a4a 	:	val_out <= 4'h91e8;
         4'h7a4b 	:	val_out <= 4'h91e8;
         4'h7a50 	:	val_out <= 4'h91cf;
         4'h7a51 	:	val_out <= 4'h91cf;
         4'h7a52 	:	val_out <= 4'h91cf;
         4'h7a53 	:	val_out <= 4'h91cf;
         4'h7a58 	:	val_out <= 4'h91b6;
         4'h7a59 	:	val_out <= 4'h91b6;
         4'h7a5a 	:	val_out <= 4'h91b6;
         4'h7a5b 	:	val_out <= 4'h91b6;
         4'h7a60 	:	val_out <= 4'h919d;
         4'h7a61 	:	val_out <= 4'h919d;
         4'h7a62 	:	val_out <= 4'h919d;
         4'h7a63 	:	val_out <= 4'h919d;
         4'h7a68 	:	val_out <= 4'h9184;
         4'h7a69 	:	val_out <= 4'h9184;
         4'h7a6a 	:	val_out <= 4'h9184;
         4'h7a6b 	:	val_out <= 4'h9184;
         4'h7a70 	:	val_out <= 4'h916b;
         4'h7a71 	:	val_out <= 4'h916b;
         4'h7a72 	:	val_out <= 4'h916b;
         4'h7a73 	:	val_out <= 4'h916b;
         4'h7a78 	:	val_out <= 4'h9152;
         4'h7a79 	:	val_out <= 4'h9152;
         4'h7a7a 	:	val_out <= 4'h9152;
         4'h7a7b 	:	val_out <= 4'h9152;
         4'h7a80 	:	val_out <= 4'h9139;
         4'h7a81 	:	val_out <= 4'h9139;
         4'h7a82 	:	val_out <= 4'h9139;
         4'h7a83 	:	val_out <= 4'h9139;
         4'h7a88 	:	val_out <= 4'h9121;
         4'h7a89 	:	val_out <= 4'h9121;
         4'h7a8a 	:	val_out <= 4'h9121;
         4'h7a8b 	:	val_out <= 4'h9121;
         4'h7a90 	:	val_out <= 4'h9108;
         4'h7a91 	:	val_out <= 4'h9108;
         4'h7a92 	:	val_out <= 4'h9108;
         4'h7a93 	:	val_out <= 4'h9108;
         4'h7a98 	:	val_out <= 4'h90ef;
         4'h7a99 	:	val_out <= 4'h90ef;
         4'h7a9a 	:	val_out <= 4'h90ef;
         4'h7a9b 	:	val_out <= 4'h90ef;
         4'h7aa0 	:	val_out <= 4'h90d6;
         4'h7aa1 	:	val_out <= 4'h90d6;
         4'h7aa2 	:	val_out <= 4'h90d6;
         4'h7aa3 	:	val_out <= 4'h90d6;
         4'h7aa8 	:	val_out <= 4'h90bd;
         4'h7aa9 	:	val_out <= 4'h90bd;
         4'h7aaa 	:	val_out <= 4'h90bd;
         4'h7aab 	:	val_out <= 4'h90bd;
         4'h7ab0 	:	val_out <= 4'h90a4;
         4'h7ab1 	:	val_out <= 4'h90a4;
         4'h7ab2 	:	val_out <= 4'h90a4;
         4'h7ab3 	:	val_out <= 4'h90a4;
         4'h7ab8 	:	val_out <= 4'h908b;
         4'h7ab9 	:	val_out <= 4'h908b;
         4'h7aba 	:	val_out <= 4'h908b;
         4'h7abb 	:	val_out <= 4'h908b;
         4'h7ac0 	:	val_out <= 4'h9072;
         4'h7ac1 	:	val_out <= 4'h9072;
         4'h7ac2 	:	val_out <= 4'h9072;
         4'h7ac3 	:	val_out <= 4'h9072;
         4'h7ac8 	:	val_out <= 4'h9059;
         4'h7ac9 	:	val_out <= 4'h9059;
         4'h7aca 	:	val_out <= 4'h9059;
         4'h7acb 	:	val_out <= 4'h9059;
         4'h7ad0 	:	val_out <= 4'h9040;
         4'h7ad1 	:	val_out <= 4'h9040;
         4'h7ad2 	:	val_out <= 4'h9040;
         4'h7ad3 	:	val_out <= 4'h9040;
         4'h7ad8 	:	val_out <= 4'h9027;
         4'h7ad9 	:	val_out <= 4'h9027;
         4'h7ada 	:	val_out <= 4'h9027;
         4'h7adb 	:	val_out <= 4'h9027;
         4'h7ae0 	:	val_out <= 4'h900e;
         4'h7ae1 	:	val_out <= 4'h900e;
         4'h7ae2 	:	val_out <= 4'h900e;
         4'h7ae3 	:	val_out <= 4'h900e;
         4'h7ae8 	:	val_out <= 4'h8ff5;
         4'h7ae9 	:	val_out <= 4'h8ff5;
         4'h7aea 	:	val_out <= 4'h8ff5;
         4'h7aeb 	:	val_out <= 4'h8ff5;
         4'h7af0 	:	val_out <= 4'h8fdd;
         4'h7af1 	:	val_out <= 4'h8fdd;
         4'h7af2 	:	val_out <= 4'h8fdd;
         4'h7af3 	:	val_out <= 4'h8fdd;
         4'h7af8 	:	val_out <= 4'h8fc4;
         4'h7af9 	:	val_out <= 4'h8fc4;
         4'h7afa 	:	val_out <= 4'h8fc4;
         4'h7afb 	:	val_out <= 4'h8fc4;
         4'h7b00 	:	val_out <= 4'h8fab;
         4'h7b01 	:	val_out <= 4'h8fab;
         4'h7b02 	:	val_out <= 4'h8fab;
         4'h7b03 	:	val_out <= 4'h8fab;
         4'h7b08 	:	val_out <= 4'h8f92;
         4'h7b09 	:	val_out <= 4'h8f92;
         4'h7b0a 	:	val_out <= 4'h8f92;
         4'h7b0b 	:	val_out <= 4'h8f92;
         4'h7b10 	:	val_out <= 4'h8f79;
         4'h7b11 	:	val_out <= 4'h8f79;
         4'h7b12 	:	val_out <= 4'h8f79;
         4'h7b13 	:	val_out <= 4'h8f79;
         4'h7b18 	:	val_out <= 4'h8f60;
         4'h7b19 	:	val_out <= 4'h8f60;
         4'h7b1a 	:	val_out <= 4'h8f60;
         4'h7b1b 	:	val_out <= 4'h8f60;
         4'h7b20 	:	val_out <= 4'h8f47;
         4'h7b21 	:	val_out <= 4'h8f47;
         4'h7b22 	:	val_out <= 4'h8f47;
         4'h7b23 	:	val_out <= 4'h8f47;
         4'h7b28 	:	val_out <= 4'h8f2e;
         4'h7b29 	:	val_out <= 4'h8f2e;
         4'h7b2a 	:	val_out <= 4'h8f2e;
         4'h7b2b 	:	val_out <= 4'h8f2e;
         4'h7b30 	:	val_out <= 4'h8f15;
         4'h7b31 	:	val_out <= 4'h8f15;
         4'h7b32 	:	val_out <= 4'h8f15;
         4'h7b33 	:	val_out <= 4'h8f15;
         4'h7b38 	:	val_out <= 4'h8efc;
         4'h7b39 	:	val_out <= 4'h8efc;
         4'h7b3a 	:	val_out <= 4'h8efc;
         4'h7b3b 	:	val_out <= 4'h8efc;
         4'h7b40 	:	val_out <= 4'h8ee3;
         4'h7b41 	:	val_out <= 4'h8ee3;
         4'h7b42 	:	val_out <= 4'h8ee3;
         4'h7b43 	:	val_out <= 4'h8ee3;
         4'h7b48 	:	val_out <= 4'h8eca;
         4'h7b49 	:	val_out <= 4'h8eca;
         4'h7b4a 	:	val_out <= 4'h8eca;
         4'h7b4b 	:	val_out <= 4'h8eca;
         4'h7b50 	:	val_out <= 4'h8eb1;
         4'h7b51 	:	val_out <= 4'h8eb1;
         4'h7b52 	:	val_out <= 4'h8eb1;
         4'h7b53 	:	val_out <= 4'h8eb1;
         4'h7b58 	:	val_out <= 4'h8e98;
         4'h7b59 	:	val_out <= 4'h8e98;
         4'h7b5a 	:	val_out <= 4'h8e98;
         4'h7b5b 	:	val_out <= 4'h8e98;
         4'h7b60 	:	val_out <= 4'h8e7f;
         4'h7b61 	:	val_out <= 4'h8e7f;
         4'h7b62 	:	val_out <= 4'h8e7f;
         4'h7b63 	:	val_out <= 4'h8e7f;
         4'h7b68 	:	val_out <= 4'h8e66;
         4'h7b69 	:	val_out <= 4'h8e66;
         4'h7b6a 	:	val_out <= 4'h8e66;
         4'h7b6b 	:	val_out <= 4'h8e66;
         4'h7b70 	:	val_out <= 4'h8e4d;
         4'h7b71 	:	val_out <= 4'h8e4d;
         4'h7b72 	:	val_out <= 4'h8e4d;
         4'h7b73 	:	val_out <= 4'h8e4d;
         4'h7b78 	:	val_out <= 4'h8e34;
         4'h7b79 	:	val_out <= 4'h8e34;
         4'h7b7a 	:	val_out <= 4'h8e34;
         4'h7b7b 	:	val_out <= 4'h8e34;
         4'h7b80 	:	val_out <= 4'h8e1b;
         4'h7b81 	:	val_out <= 4'h8e1b;
         4'h7b82 	:	val_out <= 4'h8e1b;
         4'h7b83 	:	val_out <= 4'h8e1b;
         4'h7b88 	:	val_out <= 4'h8e02;
         4'h7b89 	:	val_out <= 4'h8e02;
         4'h7b8a 	:	val_out <= 4'h8e02;
         4'h7b8b 	:	val_out <= 4'h8e02;
         4'h7b90 	:	val_out <= 4'h8de9;
         4'h7b91 	:	val_out <= 4'h8de9;
         4'h7b92 	:	val_out <= 4'h8de9;
         4'h7b93 	:	val_out <= 4'h8de9;
         4'h7b98 	:	val_out <= 4'h8dd0;
         4'h7b99 	:	val_out <= 4'h8dd0;
         4'h7b9a 	:	val_out <= 4'h8dd0;
         4'h7b9b 	:	val_out <= 4'h8dd0;
         4'h7ba0 	:	val_out <= 4'h8db7;
         4'h7ba1 	:	val_out <= 4'h8db7;
         4'h7ba2 	:	val_out <= 4'h8db7;
         4'h7ba3 	:	val_out <= 4'h8db7;
         4'h7ba8 	:	val_out <= 4'h8d9e;
         4'h7ba9 	:	val_out <= 4'h8d9e;
         4'h7baa 	:	val_out <= 4'h8d9e;
         4'h7bab 	:	val_out <= 4'h8d9e;
         4'h7bb0 	:	val_out <= 4'h8d85;
         4'h7bb1 	:	val_out <= 4'h8d85;
         4'h7bb2 	:	val_out <= 4'h8d85;
         4'h7bb3 	:	val_out <= 4'h8d85;
         4'h7bb8 	:	val_out <= 4'h8d6c;
         4'h7bb9 	:	val_out <= 4'h8d6c;
         4'h7bba 	:	val_out <= 4'h8d6c;
         4'h7bbb 	:	val_out <= 4'h8d6c;
         4'h7bc0 	:	val_out <= 4'h8d53;
         4'h7bc1 	:	val_out <= 4'h8d53;
         4'h7bc2 	:	val_out <= 4'h8d53;
         4'h7bc3 	:	val_out <= 4'h8d53;
         4'h7bc8 	:	val_out <= 4'h8d3a;
         4'h7bc9 	:	val_out <= 4'h8d3a;
         4'h7bca 	:	val_out <= 4'h8d3a;
         4'h7bcb 	:	val_out <= 4'h8d3a;
         4'h7bd0 	:	val_out <= 4'h8d21;
         4'h7bd1 	:	val_out <= 4'h8d21;
         4'h7bd2 	:	val_out <= 4'h8d21;
         4'h7bd3 	:	val_out <= 4'h8d21;
         4'h7bd8 	:	val_out <= 4'h8d08;
         4'h7bd9 	:	val_out <= 4'h8d08;
         4'h7bda 	:	val_out <= 4'h8d08;
         4'h7bdb 	:	val_out <= 4'h8d08;
         4'h7be0 	:	val_out <= 4'h8cef;
         4'h7be1 	:	val_out <= 4'h8cef;
         4'h7be2 	:	val_out <= 4'h8cef;
         4'h7be3 	:	val_out <= 4'h8cef;
         4'h7be8 	:	val_out <= 4'h8cd6;
         4'h7be9 	:	val_out <= 4'h8cd6;
         4'h7bea 	:	val_out <= 4'h8cd6;
         4'h7beb 	:	val_out <= 4'h8cd6;
         4'h7bf0 	:	val_out <= 4'h8cbd;
         4'h7bf1 	:	val_out <= 4'h8cbd;
         4'h7bf2 	:	val_out <= 4'h8cbd;
         4'h7bf3 	:	val_out <= 4'h8cbd;
         4'h7bf8 	:	val_out <= 4'h8ca4;
         4'h7bf9 	:	val_out <= 4'h8ca4;
         4'h7bfa 	:	val_out <= 4'h8ca4;
         4'h7bfb 	:	val_out <= 4'h8ca4;
         4'h7c00 	:	val_out <= 4'h8c8b;
         4'h7c01 	:	val_out <= 4'h8c8b;
         4'h7c02 	:	val_out <= 4'h8c8b;
         4'h7c03 	:	val_out <= 4'h8c8b;
         4'h7c08 	:	val_out <= 4'h8c72;
         4'h7c09 	:	val_out <= 4'h8c72;
         4'h7c0a 	:	val_out <= 4'h8c72;
         4'h7c0b 	:	val_out <= 4'h8c72;
         4'h7c10 	:	val_out <= 4'h8c59;
         4'h7c11 	:	val_out <= 4'h8c59;
         4'h7c12 	:	val_out <= 4'h8c59;
         4'h7c13 	:	val_out <= 4'h8c59;
         4'h7c18 	:	val_out <= 4'h8c40;
         4'h7c19 	:	val_out <= 4'h8c40;
         4'h7c1a 	:	val_out <= 4'h8c40;
         4'h7c1b 	:	val_out <= 4'h8c40;
         4'h7c20 	:	val_out <= 4'h8c27;
         4'h7c21 	:	val_out <= 4'h8c27;
         4'h7c22 	:	val_out <= 4'h8c27;
         4'h7c23 	:	val_out <= 4'h8c27;
         4'h7c28 	:	val_out <= 4'h8c0e;
         4'h7c29 	:	val_out <= 4'h8c0e;
         4'h7c2a 	:	val_out <= 4'h8c0e;
         4'h7c2b 	:	val_out <= 4'h8c0e;
         4'h7c30 	:	val_out <= 4'h8bf5;
         4'h7c31 	:	val_out <= 4'h8bf5;
         4'h7c32 	:	val_out <= 4'h8bf5;
         4'h7c33 	:	val_out <= 4'h8bf5;
         4'h7c38 	:	val_out <= 4'h8bdc;
         4'h7c39 	:	val_out <= 4'h8bdc;
         4'h7c3a 	:	val_out <= 4'h8bdc;
         4'h7c3b 	:	val_out <= 4'h8bdc;
         4'h7c40 	:	val_out <= 4'h8bc3;
         4'h7c41 	:	val_out <= 4'h8bc3;
         4'h7c42 	:	val_out <= 4'h8bc3;
         4'h7c43 	:	val_out <= 4'h8bc3;
         4'h7c48 	:	val_out <= 4'h8baa;
         4'h7c49 	:	val_out <= 4'h8baa;
         4'h7c4a 	:	val_out <= 4'h8baa;
         4'h7c4b 	:	val_out <= 4'h8baa;
         4'h7c50 	:	val_out <= 4'h8b91;
         4'h7c51 	:	val_out <= 4'h8b91;
         4'h7c52 	:	val_out <= 4'h8b91;
         4'h7c53 	:	val_out <= 4'h8b91;
         4'h7c58 	:	val_out <= 4'h8b78;
         4'h7c59 	:	val_out <= 4'h8b78;
         4'h7c5a 	:	val_out <= 4'h8b78;
         4'h7c5b 	:	val_out <= 4'h8b78;
         4'h7c60 	:	val_out <= 4'h8b5f;
         4'h7c61 	:	val_out <= 4'h8b5f;
         4'h7c62 	:	val_out <= 4'h8b5f;
         4'h7c63 	:	val_out <= 4'h8b5f;
         4'h7c68 	:	val_out <= 4'h8b46;
         4'h7c69 	:	val_out <= 4'h8b46;
         4'h7c6a 	:	val_out <= 4'h8b46;
         4'h7c6b 	:	val_out <= 4'h8b46;
         4'h7c70 	:	val_out <= 4'h8b2d;
         4'h7c71 	:	val_out <= 4'h8b2d;
         4'h7c72 	:	val_out <= 4'h8b2d;
         4'h7c73 	:	val_out <= 4'h8b2d;
         4'h7c78 	:	val_out <= 4'h8b14;
         4'h7c79 	:	val_out <= 4'h8b14;
         4'h7c7a 	:	val_out <= 4'h8b14;
         4'h7c7b 	:	val_out <= 4'h8b14;
         4'h7c80 	:	val_out <= 4'h8afb;
         4'h7c81 	:	val_out <= 4'h8afb;
         4'h7c82 	:	val_out <= 4'h8afb;
         4'h7c83 	:	val_out <= 4'h8afb;
         4'h7c88 	:	val_out <= 4'h8ae2;
         4'h7c89 	:	val_out <= 4'h8ae2;
         4'h7c8a 	:	val_out <= 4'h8ae2;
         4'h7c8b 	:	val_out <= 4'h8ae2;
         4'h7c90 	:	val_out <= 4'h8ac9;
         4'h7c91 	:	val_out <= 4'h8ac9;
         4'h7c92 	:	val_out <= 4'h8ac9;
         4'h7c93 	:	val_out <= 4'h8ac9;
         4'h7c98 	:	val_out <= 4'h8ab0;
         4'h7c99 	:	val_out <= 4'h8ab0;
         4'h7c9a 	:	val_out <= 4'h8ab0;
         4'h7c9b 	:	val_out <= 4'h8ab0;
         4'h7ca0 	:	val_out <= 4'h8a97;
         4'h7ca1 	:	val_out <= 4'h8a97;
         4'h7ca2 	:	val_out <= 4'h8a97;
         4'h7ca3 	:	val_out <= 4'h8a97;
         4'h7ca8 	:	val_out <= 4'h8a7e;
         4'h7ca9 	:	val_out <= 4'h8a7e;
         4'h7caa 	:	val_out <= 4'h8a7e;
         4'h7cab 	:	val_out <= 4'h8a7e;
         4'h7cb0 	:	val_out <= 4'h8a65;
         4'h7cb1 	:	val_out <= 4'h8a65;
         4'h7cb2 	:	val_out <= 4'h8a65;
         4'h7cb3 	:	val_out <= 4'h8a65;
         4'h7cb8 	:	val_out <= 4'h8a4c;
         4'h7cb9 	:	val_out <= 4'h8a4c;
         4'h7cba 	:	val_out <= 4'h8a4c;
         4'h7cbb 	:	val_out <= 4'h8a4c;
         4'h7cc0 	:	val_out <= 4'h8a33;
         4'h7cc1 	:	val_out <= 4'h8a33;
         4'h7cc2 	:	val_out <= 4'h8a33;
         4'h7cc3 	:	val_out <= 4'h8a33;
         4'h7cc8 	:	val_out <= 4'h8a19;
         4'h7cc9 	:	val_out <= 4'h8a19;
         4'h7cca 	:	val_out <= 4'h8a19;
         4'h7ccb 	:	val_out <= 4'h8a19;
         4'h7cd0 	:	val_out <= 4'h8a00;
         4'h7cd1 	:	val_out <= 4'h8a00;
         4'h7cd2 	:	val_out <= 4'h8a00;
         4'h7cd3 	:	val_out <= 4'h8a00;
         4'h7cd8 	:	val_out <= 4'h89e7;
         4'h7cd9 	:	val_out <= 4'h89e7;
         4'h7cda 	:	val_out <= 4'h89e7;
         4'h7cdb 	:	val_out <= 4'h89e7;
         4'h7ce0 	:	val_out <= 4'h89ce;
         4'h7ce1 	:	val_out <= 4'h89ce;
         4'h7ce2 	:	val_out <= 4'h89ce;
         4'h7ce3 	:	val_out <= 4'h89ce;
         4'h7ce8 	:	val_out <= 4'h89b5;
         4'h7ce9 	:	val_out <= 4'h89b5;
         4'h7cea 	:	val_out <= 4'h89b5;
         4'h7ceb 	:	val_out <= 4'h89b5;
         4'h7cf0 	:	val_out <= 4'h899c;
         4'h7cf1 	:	val_out <= 4'h899c;
         4'h7cf2 	:	val_out <= 4'h899c;
         4'h7cf3 	:	val_out <= 4'h899c;
         4'h7cf8 	:	val_out <= 4'h8983;
         4'h7cf9 	:	val_out <= 4'h8983;
         4'h7cfa 	:	val_out <= 4'h8983;
         4'h7cfb 	:	val_out <= 4'h8983;
         4'h7d00 	:	val_out <= 4'h896a;
         4'h7d01 	:	val_out <= 4'h896a;
         4'h7d02 	:	val_out <= 4'h896a;
         4'h7d03 	:	val_out <= 4'h896a;
         4'h7d08 	:	val_out <= 4'h8951;
         4'h7d09 	:	val_out <= 4'h8951;
         4'h7d0a 	:	val_out <= 4'h8951;
         4'h7d0b 	:	val_out <= 4'h8951;
         4'h7d10 	:	val_out <= 4'h8938;
         4'h7d11 	:	val_out <= 4'h8938;
         4'h7d12 	:	val_out <= 4'h8938;
         4'h7d13 	:	val_out <= 4'h8938;
         4'h7d18 	:	val_out <= 4'h891f;
         4'h7d19 	:	val_out <= 4'h891f;
         4'h7d1a 	:	val_out <= 4'h891f;
         4'h7d1b 	:	val_out <= 4'h891f;
         4'h7d20 	:	val_out <= 4'h8906;
         4'h7d21 	:	val_out <= 4'h8906;
         4'h7d22 	:	val_out <= 4'h8906;
         4'h7d23 	:	val_out <= 4'h8906;
         4'h7d28 	:	val_out <= 4'h88ed;
         4'h7d29 	:	val_out <= 4'h88ed;
         4'h7d2a 	:	val_out <= 4'h88ed;
         4'h7d2b 	:	val_out <= 4'h88ed;
         4'h7d30 	:	val_out <= 4'h88d4;
         4'h7d31 	:	val_out <= 4'h88d4;
         4'h7d32 	:	val_out <= 4'h88d4;
         4'h7d33 	:	val_out <= 4'h88d4;
         4'h7d38 	:	val_out <= 4'h88bb;
         4'h7d39 	:	val_out <= 4'h88bb;
         4'h7d3a 	:	val_out <= 4'h88bb;
         4'h7d3b 	:	val_out <= 4'h88bb;
         4'h7d40 	:	val_out <= 4'h88a2;
         4'h7d41 	:	val_out <= 4'h88a2;
         4'h7d42 	:	val_out <= 4'h88a2;
         4'h7d43 	:	val_out <= 4'h88a2;
         4'h7d48 	:	val_out <= 4'h8888;
         4'h7d49 	:	val_out <= 4'h8888;
         4'h7d4a 	:	val_out <= 4'h8888;
         4'h7d4b 	:	val_out <= 4'h8888;
         4'h7d50 	:	val_out <= 4'h886f;
         4'h7d51 	:	val_out <= 4'h886f;
         4'h7d52 	:	val_out <= 4'h886f;
         4'h7d53 	:	val_out <= 4'h886f;
         4'h7d58 	:	val_out <= 4'h8856;
         4'h7d59 	:	val_out <= 4'h8856;
         4'h7d5a 	:	val_out <= 4'h8856;
         4'h7d5b 	:	val_out <= 4'h8856;
         4'h7d60 	:	val_out <= 4'h883d;
         4'h7d61 	:	val_out <= 4'h883d;
         4'h7d62 	:	val_out <= 4'h883d;
         4'h7d63 	:	val_out <= 4'h883d;
         4'h7d68 	:	val_out <= 4'h8824;
         4'h7d69 	:	val_out <= 4'h8824;
         4'h7d6a 	:	val_out <= 4'h8824;
         4'h7d6b 	:	val_out <= 4'h8824;
         4'h7d70 	:	val_out <= 4'h880b;
         4'h7d71 	:	val_out <= 4'h880b;
         4'h7d72 	:	val_out <= 4'h880b;
         4'h7d73 	:	val_out <= 4'h880b;
         4'h7d78 	:	val_out <= 4'h87f2;
         4'h7d79 	:	val_out <= 4'h87f2;
         4'h7d7a 	:	val_out <= 4'h87f2;
         4'h7d7b 	:	val_out <= 4'h87f2;
         4'h7d80 	:	val_out <= 4'h87d9;
         4'h7d81 	:	val_out <= 4'h87d9;
         4'h7d82 	:	val_out <= 4'h87d9;
         4'h7d83 	:	val_out <= 4'h87d9;
         4'h7d88 	:	val_out <= 4'h87c0;
         4'h7d89 	:	val_out <= 4'h87c0;
         4'h7d8a 	:	val_out <= 4'h87c0;
         4'h7d8b 	:	val_out <= 4'h87c0;
         4'h7d90 	:	val_out <= 4'h87a7;
         4'h7d91 	:	val_out <= 4'h87a7;
         4'h7d92 	:	val_out <= 4'h87a7;
         4'h7d93 	:	val_out <= 4'h87a7;
         4'h7d98 	:	val_out <= 4'h878e;
         4'h7d99 	:	val_out <= 4'h878e;
         4'h7d9a 	:	val_out <= 4'h878e;
         4'h7d9b 	:	val_out <= 4'h878e;
         4'h7da0 	:	val_out <= 4'h8775;
         4'h7da1 	:	val_out <= 4'h8775;
         4'h7da2 	:	val_out <= 4'h8775;
         4'h7da3 	:	val_out <= 4'h8775;
         4'h7da8 	:	val_out <= 4'h875b;
         4'h7da9 	:	val_out <= 4'h875b;
         4'h7daa 	:	val_out <= 4'h875b;
         4'h7dab 	:	val_out <= 4'h875b;
         4'h7db0 	:	val_out <= 4'h8742;
         4'h7db1 	:	val_out <= 4'h8742;
         4'h7db2 	:	val_out <= 4'h8742;
         4'h7db3 	:	val_out <= 4'h8742;
         4'h7db8 	:	val_out <= 4'h8729;
         4'h7db9 	:	val_out <= 4'h8729;
         4'h7dba 	:	val_out <= 4'h8729;
         4'h7dbb 	:	val_out <= 4'h8729;
         4'h7dc0 	:	val_out <= 4'h8710;
         4'h7dc1 	:	val_out <= 4'h8710;
         4'h7dc2 	:	val_out <= 4'h8710;
         4'h7dc3 	:	val_out <= 4'h8710;
         4'h7dc8 	:	val_out <= 4'h86f7;
         4'h7dc9 	:	val_out <= 4'h86f7;
         4'h7dca 	:	val_out <= 4'h86f7;
         4'h7dcb 	:	val_out <= 4'h86f7;
         4'h7dd0 	:	val_out <= 4'h86de;
         4'h7dd1 	:	val_out <= 4'h86de;
         4'h7dd2 	:	val_out <= 4'h86de;
         4'h7dd3 	:	val_out <= 4'h86de;
         4'h7dd8 	:	val_out <= 4'h86c5;
         4'h7dd9 	:	val_out <= 4'h86c5;
         4'h7dda 	:	val_out <= 4'h86c5;
         4'h7ddb 	:	val_out <= 4'h86c5;
         4'h7de0 	:	val_out <= 4'h86ac;
         4'h7de1 	:	val_out <= 4'h86ac;
         4'h7de2 	:	val_out <= 4'h86ac;
         4'h7de3 	:	val_out <= 4'h86ac;
         4'h7de8 	:	val_out <= 4'h8693;
         4'h7de9 	:	val_out <= 4'h8693;
         4'h7dea 	:	val_out <= 4'h8693;
         4'h7deb 	:	val_out <= 4'h8693;
         4'h7df0 	:	val_out <= 4'h867a;
         4'h7df1 	:	val_out <= 4'h867a;
         4'h7df2 	:	val_out <= 4'h867a;
         4'h7df3 	:	val_out <= 4'h867a;
         4'h7df8 	:	val_out <= 4'h8660;
         4'h7df9 	:	val_out <= 4'h8660;
         4'h7dfa 	:	val_out <= 4'h8660;
         4'h7dfb 	:	val_out <= 4'h8660;
         4'h7e00 	:	val_out <= 4'h8647;
         4'h7e01 	:	val_out <= 4'h8647;
         4'h7e02 	:	val_out <= 4'h8647;
         4'h7e03 	:	val_out <= 4'h8647;
         4'h7e08 	:	val_out <= 4'h862e;
         4'h7e09 	:	val_out <= 4'h862e;
         4'h7e0a 	:	val_out <= 4'h862e;
         4'h7e0b 	:	val_out <= 4'h862e;
         4'h7e10 	:	val_out <= 4'h8615;
         4'h7e11 	:	val_out <= 4'h8615;
         4'h7e12 	:	val_out <= 4'h8615;
         4'h7e13 	:	val_out <= 4'h8615;
         4'h7e18 	:	val_out <= 4'h85fc;
         4'h7e19 	:	val_out <= 4'h85fc;
         4'h7e1a 	:	val_out <= 4'h85fc;
         4'h7e1b 	:	val_out <= 4'h85fc;
         4'h7e20 	:	val_out <= 4'h85e3;
         4'h7e21 	:	val_out <= 4'h85e3;
         4'h7e22 	:	val_out <= 4'h85e3;
         4'h7e23 	:	val_out <= 4'h85e3;
         4'h7e28 	:	val_out <= 4'h85ca;
         4'h7e29 	:	val_out <= 4'h85ca;
         4'h7e2a 	:	val_out <= 4'h85ca;
         4'h7e2b 	:	val_out <= 4'h85ca;
         4'h7e30 	:	val_out <= 4'h85b1;
         4'h7e31 	:	val_out <= 4'h85b1;
         4'h7e32 	:	val_out <= 4'h85b1;
         4'h7e33 	:	val_out <= 4'h85b1;
         4'h7e38 	:	val_out <= 4'h8598;
         4'h7e39 	:	val_out <= 4'h8598;
         4'h7e3a 	:	val_out <= 4'h8598;
         4'h7e3b 	:	val_out <= 4'h8598;
         4'h7e40 	:	val_out <= 4'h857f;
         4'h7e41 	:	val_out <= 4'h857f;
         4'h7e42 	:	val_out <= 4'h857f;
         4'h7e43 	:	val_out <= 4'h857f;
         4'h7e48 	:	val_out <= 4'h8565;
         4'h7e49 	:	val_out <= 4'h8565;
         4'h7e4a 	:	val_out <= 4'h8565;
         4'h7e4b 	:	val_out <= 4'h8565;
         4'h7e50 	:	val_out <= 4'h854c;
         4'h7e51 	:	val_out <= 4'h854c;
         4'h7e52 	:	val_out <= 4'h854c;
         4'h7e53 	:	val_out <= 4'h854c;
         4'h7e58 	:	val_out <= 4'h8533;
         4'h7e59 	:	val_out <= 4'h8533;
         4'h7e5a 	:	val_out <= 4'h8533;
         4'h7e5b 	:	val_out <= 4'h8533;
         4'h7e60 	:	val_out <= 4'h851a;
         4'h7e61 	:	val_out <= 4'h851a;
         4'h7e62 	:	val_out <= 4'h851a;
         4'h7e63 	:	val_out <= 4'h851a;
         4'h7e68 	:	val_out <= 4'h8501;
         4'h7e69 	:	val_out <= 4'h8501;
         4'h7e6a 	:	val_out <= 4'h8501;
         4'h7e6b 	:	val_out <= 4'h8501;
         4'h7e70 	:	val_out <= 4'h84e8;
         4'h7e71 	:	val_out <= 4'h84e8;
         4'h7e72 	:	val_out <= 4'h84e8;
         4'h7e73 	:	val_out <= 4'h84e8;
         4'h7e78 	:	val_out <= 4'h84cf;
         4'h7e79 	:	val_out <= 4'h84cf;
         4'h7e7a 	:	val_out <= 4'h84cf;
         4'h7e7b 	:	val_out <= 4'h84cf;
         4'h7e80 	:	val_out <= 4'h84b6;
         4'h7e81 	:	val_out <= 4'h84b6;
         4'h7e82 	:	val_out <= 4'h84b6;
         4'h7e83 	:	val_out <= 4'h84b6;
         4'h7e88 	:	val_out <= 4'h849c;
         4'h7e89 	:	val_out <= 4'h849c;
         4'h7e8a 	:	val_out <= 4'h849c;
         4'h7e8b 	:	val_out <= 4'h849c;
         4'h7e90 	:	val_out <= 4'h8483;
         4'h7e91 	:	val_out <= 4'h8483;
         4'h7e92 	:	val_out <= 4'h8483;
         4'h7e93 	:	val_out <= 4'h8483;
         4'h7e98 	:	val_out <= 4'h846a;
         4'h7e99 	:	val_out <= 4'h846a;
         4'h7e9a 	:	val_out <= 4'h846a;
         4'h7e9b 	:	val_out <= 4'h846a;
         4'h7ea0 	:	val_out <= 4'h8451;
         4'h7ea1 	:	val_out <= 4'h8451;
         4'h7ea2 	:	val_out <= 4'h8451;
         4'h7ea3 	:	val_out <= 4'h8451;
         4'h7ea8 	:	val_out <= 4'h8438;
         4'h7ea9 	:	val_out <= 4'h8438;
         4'h7eaa 	:	val_out <= 4'h8438;
         4'h7eab 	:	val_out <= 4'h8438;
         4'h7eb0 	:	val_out <= 4'h841f;
         4'h7eb1 	:	val_out <= 4'h841f;
         4'h7eb2 	:	val_out <= 4'h841f;
         4'h7eb3 	:	val_out <= 4'h841f;
         4'h7eb8 	:	val_out <= 4'h8406;
         4'h7eb9 	:	val_out <= 4'h8406;
         4'h7eba 	:	val_out <= 4'h8406;
         4'h7ebb 	:	val_out <= 4'h8406;
         4'h7ec0 	:	val_out <= 4'h83ed;
         4'h7ec1 	:	val_out <= 4'h83ed;
         4'h7ec2 	:	val_out <= 4'h83ed;
         4'h7ec3 	:	val_out <= 4'h83ed;
         4'h7ec8 	:	val_out <= 4'h83d4;
         4'h7ec9 	:	val_out <= 4'h83d4;
         4'h7eca 	:	val_out <= 4'h83d4;
         4'h7ecb 	:	val_out <= 4'h83d4;
         4'h7ed0 	:	val_out <= 4'h83ba;
         4'h7ed1 	:	val_out <= 4'h83ba;
         4'h7ed2 	:	val_out <= 4'h83ba;
         4'h7ed3 	:	val_out <= 4'h83ba;
         4'h7ed8 	:	val_out <= 4'h83a1;
         4'h7ed9 	:	val_out <= 4'h83a1;
         4'h7eda 	:	val_out <= 4'h83a1;
         4'h7edb 	:	val_out <= 4'h83a1;
         4'h7ee0 	:	val_out <= 4'h8388;
         4'h7ee1 	:	val_out <= 4'h8388;
         4'h7ee2 	:	val_out <= 4'h8388;
         4'h7ee3 	:	val_out <= 4'h8388;
         4'h7ee8 	:	val_out <= 4'h836f;
         4'h7ee9 	:	val_out <= 4'h836f;
         4'h7eea 	:	val_out <= 4'h836f;
         4'h7eeb 	:	val_out <= 4'h836f;
         4'h7ef0 	:	val_out <= 4'h8356;
         4'h7ef1 	:	val_out <= 4'h8356;
         4'h7ef2 	:	val_out <= 4'h8356;
         4'h7ef3 	:	val_out <= 4'h8356;
         4'h7ef8 	:	val_out <= 4'h833d;
         4'h7ef9 	:	val_out <= 4'h833d;
         4'h7efa 	:	val_out <= 4'h833d;
         4'h7efb 	:	val_out <= 4'h833d;
         4'h7f00 	:	val_out <= 4'h8324;
         4'h7f01 	:	val_out <= 4'h8324;
         4'h7f02 	:	val_out <= 4'h8324;
         4'h7f03 	:	val_out <= 4'h8324;
         4'h7f08 	:	val_out <= 4'h830b;
         4'h7f09 	:	val_out <= 4'h830b;
         4'h7f0a 	:	val_out <= 4'h830b;
         4'h7f0b 	:	val_out <= 4'h830b;
         4'h7f10 	:	val_out <= 4'h82f1;
         4'h7f11 	:	val_out <= 4'h82f1;
         4'h7f12 	:	val_out <= 4'h82f1;
         4'h7f13 	:	val_out <= 4'h82f1;
         4'h7f18 	:	val_out <= 4'h82d8;
         4'h7f19 	:	val_out <= 4'h82d8;
         4'h7f1a 	:	val_out <= 4'h82d8;
         4'h7f1b 	:	val_out <= 4'h82d8;
         4'h7f20 	:	val_out <= 4'h82bf;
         4'h7f21 	:	val_out <= 4'h82bf;
         4'h7f22 	:	val_out <= 4'h82bf;
         4'h7f23 	:	val_out <= 4'h82bf;
         4'h7f28 	:	val_out <= 4'h82a6;
         4'h7f29 	:	val_out <= 4'h82a6;
         4'h7f2a 	:	val_out <= 4'h82a6;
         4'h7f2b 	:	val_out <= 4'h82a6;
         4'h7f30 	:	val_out <= 4'h828d;
         4'h7f31 	:	val_out <= 4'h828d;
         4'h7f32 	:	val_out <= 4'h828d;
         4'h7f33 	:	val_out <= 4'h828d;
         4'h7f38 	:	val_out <= 4'h8274;
         4'h7f39 	:	val_out <= 4'h8274;
         4'h7f3a 	:	val_out <= 4'h8274;
         4'h7f3b 	:	val_out <= 4'h8274;
         4'h7f40 	:	val_out <= 4'h825b;
         4'h7f41 	:	val_out <= 4'h825b;
         4'h7f42 	:	val_out <= 4'h825b;
         4'h7f43 	:	val_out <= 4'h825b;
         4'h7f48 	:	val_out <= 4'h8242;
         4'h7f49 	:	val_out <= 4'h8242;
         4'h7f4a 	:	val_out <= 4'h8242;
         4'h7f4b 	:	val_out <= 4'h8242;
         4'h7f50 	:	val_out <= 4'h8228;
         4'h7f51 	:	val_out <= 4'h8228;
         4'h7f52 	:	val_out <= 4'h8228;
         4'h7f53 	:	val_out <= 4'h8228;
         4'h7f58 	:	val_out <= 4'h820f;
         4'h7f59 	:	val_out <= 4'h820f;
         4'h7f5a 	:	val_out <= 4'h820f;
         4'h7f5b 	:	val_out <= 4'h820f;
         4'h7f60 	:	val_out <= 4'h81f6;
         4'h7f61 	:	val_out <= 4'h81f6;
         4'h7f62 	:	val_out <= 4'h81f6;
         4'h7f63 	:	val_out <= 4'h81f6;
         4'h7f68 	:	val_out <= 4'h81dd;
         4'h7f69 	:	val_out <= 4'h81dd;
         4'h7f6a 	:	val_out <= 4'h81dd;
         4'h7f6b 	:	val_out <= 4'h81dd;
         4'h7f70 	:	val_out <= 4'h81c4;
         4'h7f71 	:	val_out <= 4'h81c4;
         4'h7f72 	:	val_out <= 4'h81c4;
         4'h7f73 	:	val_out <= 4'h81c4;
         4'h7f78 	:	val_out <= 4'h81ab;
         4'h7f79 	:	val_out <= 4'h81ab;
         4'h7f7a 	:	val_out <= 4'h81ab;
         4'h7f7b 	:	val_out <= 4'h81ab;
         4'h7f80 	:	val_out <= 4'h8192;
         4'h7f81 	:	val_out <= 4'h8192;
         4'h7f82 	:	val_out <= 4'h8192;
         4'h7f83 	:	val_out <= 4'h8192;
         4'h7f88 	:	val_out <= 4'h8178;
         4'h7f89 	:	val_out <= 4'h8178;
         4'h7f8a 	:	val_out <= 4'h8178;
         4'h7f8b 	:	val_out <= 4'h8178;
         4'h7f90 	:	val_out <= 4'h815f;
         4'h7f91 	:	val_out <= 4'h815f;
         4'h7f92 	:	val_out <= 4'h815f;
         4'h7f93 	:	val_out <= 4'h815f;
         4'h7f98 	:	val_out <= 4'h8146;
         4'h7f99 	:	val_out <= 4'h8146;
         4'h7f9a 	:	val_out <= 4'h8146;
         4'h7f9b 	:	val_out <= 4'h8146;
         4'h7fa0 	:	val_out <= 4'h812d;
         4'h7fa1 	:	val_out <= 4'h812d;
         4'h7fa2 	:	val_out <= 4'h812d;
         4'h7fa3 	:	val_out <= 4'h812d;
         4'h7fa8 	:	val_out <= 4'h8114;
         4'h7fa9 	:	val_out <= 4'h8114;
         4'h7faa 	:	val_out <= 4'h8114;
         4'h7fab 	:	val_out <= 4'h8114;
         4'h7fb0 	:	val_out <= 4'h80fb;
         4'h7fb1 	:	val_out <= 4'h80fb;
         4'h7fb2 	:	val_out <= 4'h80fb;
         4'h7fb3 	:	val_out <= 4'h80fb;
         4'h7fb8 	:	val_out <= 4'h80e2;
         4'h7fb9 	:	val_out <= 4'h80e2;
         4'h7fba 	:	val_out <= 4'h80e2;
         4'h7fbb 	:	val_out <= 4'h80e2;
         4'h7fc0 	:	val_out <= 4'h80c9;
         4'h7fc1 	:	val_out <= 4'h80c9;
         4'h7fc2 	:	val_out <= 4'h80c9;
         4'h7fc3 	:	val_out <= 4'h80c9;
         4'h7fc8 	:	val_out <= 4'h80af;
         4'h7fc9 	:	val_out <= 4'h80af;
         4'h7fca 	:	val_out <= 4'h80af;
         4'h7fcb 	:	val_out <= 4'h80af;
         4'h7fd0 	:	val_out <= 4'h8096;
         4'h7fd1 	:	val_out <= 4'h8096;
         4'h7fd2 	:	val_out <= 4'h8096;
         4'h7fd3 	:	val_out <= 4'h8096;
         4'h7fd8 	:	val_out <= 4'h807d;
         4'h7fd9 	:	val_out <= 4'h807d;
         4'h7fda 	:	val_out <= 4'h807d;
         4'h7fdb 	:	val_out <= 4'h807d;
         4'h7fe0 	:	val_out <= 4'h8064;
         4'h7fe1 	:	val_out <= 4'h8064;
         4'h7fe2 	:	val_out <= 4'h8064;
         4'h7fe3 	:	val_out <= 4'h8064;
         4'h7fe8 	:	val_out <= 4'h804b;
         4'h7fe9 	:	val_out <= 4'h804b;
         4'h7fea 	:	val_out <= 4'h804b;
         4'h7feb 	:	val_out <= 4'h804b;
         4'h7ff0 	:	val_out <= 4'h8032;
         4'h7ff1 	:	val_out <= 4'h8032;
         4'h7ff2 	:	val_out <= 4'h8032;
         4'h7ff3 	:	val_out <= 4'h8032;
         4'h7ff8 	:	val_out <= 4'h8019;
         4'h7ff9 	:	val_out <= 4'h8019;
         4'h7ffa 	:	val_out <= 4'h8019;
         4'h7ffb 	:	val_out <= 4'h8019;
         4'h8000 	:	val_out <= 4'h8000;
         4'h8001 	:	val_out <= 4'h8000;
         4'h8002 	:	val_out <= 4'h8000;
         4'h8003 	:	val_out <= 4'h8000;
         4'h8008 	:	val_out <= 4'h7fe6;
         4'h8009 	:	val_out <= 4'h7fe6;
         4'h800a 	:	val_out <= 4'h7fe6;
         4'h800b 	:	val_out <= 4'h7fe6;
         4'h8010 	:	val_out <= 4'h7fcd;
         4'h8011 	:	val_out <= 4'h7fcd;
         4'h8012 	:	val_out <= 4'h7fcd;
         4'h8013 	:	val_out <= 4'h7fcd;
         4'h8018 	:	val_out <= 4'h7fb4;
         4'h8019 	:	val_out <= 4'h7fb4;
         4'h801a 	:	val_out <= 4'h7fb4;
         4'h801b 	:	val_out <= 4'h7fb4;
         4'h8020 	:	val_out <= 4'h7f9b;
         4'h8021 	:	val_out <= 4'h7f9b;
         4'h8022 	:	val_out <= 4'h7f9b;
         4'h8023 	:	val_out <= 4'h7f9b;
         4'h8028 	:	val_out <= 4'h7f82;
         4'h8029 	:	val_out <= 4'h7f82;
         4'h802a 	:	val_out <= 4'h7f82;
         4'h802b 	:	val_out <= 4'h7f82;
         4'h8030 	:	val_out <= 4'h7f69;
         4'h8031 	:	val_out <= 4'h7f69;
         4'h8032 	:	val_out <= 4'h7f69;
         4'h8033 	:	val_out <= 4'h7f69;
         4'h8038 	:	val_out <= 4'h7f50;
         4'h8039 	:	val_out <= 4'h7f50;
         4'h803a 	:	val_out <= 4'h7f50;
         4'h803b 	:	val_out <= 4'h7f50;
         4'h8040 	:	val_out <= 4'h7f36;
         4'h8041 	:	val_out <= 4'h7f36;
         4'h8042 	:	val_out <= 4'h7f36;
         4'h8043 	:	val_out <= 4'h7f36;
         4'h8048 	:	val_out <= 4'h7f1d;
         4'h8049 	:	val_out <= 4'h7f1d;
         4'h804a 	:	val_out <= 4'h7f1d;
         4'h804b 	:	val_out <= 4'h7f1d;
         4'h8050 	:	val_out <= 4'h7f04;
         4'h8051 	:	val_out <= 4'h7f04;
         4'h8052 	:	val_out <= 4'h7f04;
         4'h8053 	:	val_out <= 4'h7f04;
         4'h8058 	:	val_out <= 4'h7eeb;
         4'h8059 	:	val_out <= 4'h7eeb;
         4'h805a 	:	val_out <= 4'h7eeb;
         4'h805b 	:	val_out <= 4'h7eeb;
         4'h8060 	:	val_out <= 4'h7ed2;
         4'h8061 	:	val_out <= 4'h7ed2;
         4'h8062 	:	val_out <= 4'h7ed2;
         4'h8063 	:	val_out <= 4'h7ed2;
         4'h8068 	:	val_out <= 4'h7eb9;
         4'h8069 	:	val_out <= 4'h7eb9;
         4'h806a 	:	val_out <= 4'h7eb9;
         4'h806b 	:	val_out <= 4'h7eb9;
         4'h8070 	:	val_out <= 4'h7ea0;
         4'h8071 	:	val_out <= 4'h7ea0;
         4'h8072 	:	val_out <= 4'h7ea0;
         4'h8073 	:	val_out <= 4'h7ea0;
         4'h8078 	:	val_out <= 4'h7e87;
         4'h8079 	:	val_out <= 4'h7e87;
         4'h807a 	:	val_out <= 4'h7e87;
         4'h807b 	:	val_out <= 4'h7e87;
         4'h8080 	:	val_out <= 4'h7e6d;
         4'h8081 	:	val_out <= 4'h7e6d;
         4'h8082 	:	val_out <= 4'h7e6d;
         4'h8083 	:	val_out <= 4'h7e6d;
         4'h8088 	:	val_out <= 4'h7e54;
         4'h8089 	:	val_out <= 4'h7e54;
         4'h808a 	:	val_out <= 4'h7e54;
         4'h808b 	:	val_out <= 4'h7e54;
         4'h8090 	:	val_out <= 4'h7e3b;
         4'h8091 	:	val_out <= 4'h7e3b;
         4'h8092 	:	val_out <= 4'h7e3b;
         4'h8093 	:	val_out <= 4'h7e3b;
         4'h8098 	:	val_out <= 4'h7e22;
         4'h8099 	:	val_out <= 4'h7e22;
         4'h809a 	:	val_out <= 4'h7e22;
         4'h809b 	:	val_out <= 4'h7e22;
         4'h80a0 	:	val_out <= 4'h7e09;
         4'h80a1 	:	val_out <= 4'h7e09;
         4'h80a2 	:	val_out <= 4'h7e09;
         4'h80a3 	:	val_out <= 4'h7e09;
         4'h80a8 	:	val_out <= 4'h7df0;
         4'h80a9 	:	val_out <= 4'h7df0;
         4'h80aa 	:	val_out <= 4'h7df0;
         4'h80ab 	:	val_out <= 4'h7df0;
         4'h80b0 	:	val_out <= 4'h7dd7;
         4'h80b1 	:	val_out <= 4'h7dd7;
         4'h80b2 	:	val_out <= 4'h7dd7;
         4'h80b3 	:	val_out <= 4'h7dd7;
         4'h80b8 	:	val_out <= 4'h7dbd;
         4'h80b9 	:	val_out <= 4'h7dbd;
         4'h80ba 	:	val_out <= 4'h7dbd;
         4'h80bb 	:	val_out <= 4'h7dbd;
         4'h80c0 	:	val_out <= 4'h7da4;
         4'h80c1 	:	val_out <= 4'h7da4;
         4'h80c2 	:	val_out <= 4'h7da4;
         4'h80c3 	:	val_out <= 4'h7da4;
         4'h80c8 	:	val_out <= 4'h7d8b;
         4'h80c9 	:	val_out <= 4'h7d8b;
         4'h80ca 	:	val_out <= 4'h7d8b;
         4'h80cb 	:	val_out <= 4'h7d8b;
         4'h80d0 	:	val_out <= 4'h7d72;
         4'h80d1 	:	val_out <= 4'h7d72;
         4'h80d2 	:	val_out <= 4'h7d72;
         4'h80d3 	:	val_out <= 4'h7d72;
         4'h80d8 	:	val_out <= 4'h7d59;
         4'h80d9 	:	val_out <= 4'h7d59;
         4'h80da 	:	val_out <= 4'h7d59;
         4'h80db 	:	val_out <= 4'h7d59;
         4'h80e0 	:	val_out <= 4'h7d40;
         4'h80e1 	:	val_out <= 4'h7d40;
         4'h80e2 	:	val_out <= 4'h7d40;
         4'h80e3 	:	val_out <= 4'h7d40;
         4'h80e8 	:	val_out <= 4'h7d27;
         4'h80e9 	:	val_out <= 4'h7d27;
         4'h80ea 	:	val_out <= 4'h7d27;
         4'h80eb 	:	val_out <= 4'h7d27;
         4'h80f0 	:	val_out <= 4'h7d0e;
         4'h80f1 	:	val_out <= 4'h7d0e;
         4'h80f2 	:	val_out <= 4'h7d0e;
         4'h80f3 	:	val_out <= 4'h7d0e;
         4'h80f8 	:	val_out <= 4'h7cf4;
         4'h80f9 	:	val_out <= 4'h7cf4;
         4'h80fa 	:	val_out <= 4'h7cf4;
         4'h80fb 	:	val_out <= 4'h7cf4;
         4'h8100 	:	val_out <= 4'h7cdb;
         4'h8101 	:	val_out <= 4'h7cdb;
         4'h8102 	:	val_out <= 4'h7cdb;
         4'h8103 	:	val_out <= 4'h7cdb;
         4'h8108 	:	val_out <= 4'h7cc2;
         4'h8109 	:	val_out <= 4'h7cc2;
         4'h810a 	:	val_out <= 4'h7cc2;
         4'h810b 	:	val_out <= 4'h7cc2;
         4'h8110 	:	val_out <= 4'h7ca9;
         4'h8111 	:	val_out <= 4'h7ca9;
         4'h8112 	:	val_out <= 4'h7ca9;
         4'h8113 	:	val_out <= 4'h7ca9;
         4'h8118 	:	val_out <= 4'h7c90;
         4'h8119 	:	val_out <= 4'h7c90;
         4'h811a 	:	val_out <= 4'h7c90;
         4'h811b 	:	val_out <= 4'h7c90;
         4'h8120 	:	val_out <= 4'h7c77;
         4'h8121 	:	val_out <= 4'h7c77;
         4'h8122 	:	val_out <= 4'h7c77;
         4'h8123 	:	val_out <= 4'h7c77;
         4'h8128 	:	val_out <= 4'h7c5e;
         4'h8129 	:	val_out <= 4'h7c5e;
         4'h812a 	:	val_out <= 4'h7c5e;
         4'h812b 	:	val_out <= 4'h7c5e;
         4'h8130 	:	val_out <= 4'h7c45;
         4'h8131 	:	val_out <= 4'h7c45;
         4'h8132 	:	val_out <= 4'h7c45;
         4'h8133 	:	val_out <= 4'h7c45;
         4'h8138 	:	val_out <= 4'h7c2b;
         4'h8139 	:	val_out <= 4'h7c2b;
         4'h813a 	:	val_out <= 4'h7c2b;
         4'h813b 	:	val_out <= 4'h7c2b;
         4'h8140 	:	val_out <= 4'h7c12;
         4'h8141 	:	val_out <= 4'h7c12;
         4'h8142 	:	val_out <= 4'h7c12;
         4'h8143 	:	val_out <= 4'h7c12;
         4'h8148 	:	val_out <= 4'h7bf9;
         4'h8149 	:	val_out <= 4'h7bf9;
         4'h814a 	:	val_out <= 4'h7bf9;
         4'h814b 	:	val_out <= 4'h7bf9;
         4'h8150 	:	val_out <= 4'h7be0;
         4'h8151 	:	val_out <= 4'h7be0;
         4'h8152 	:	val_out <= 4'h7be0;
         4'h8153 	:	val_out <= 4'h7be0;
         4'h8158 	:	val_out <= 4'h7bc7;
         4'h8159 	:	val_out <= 4'h7bc7;
         4'h815a 	:	val_out <= 4'h7bc7;
         4'h815b 	:	val_out <= 4'h7bc7;
         4'h8160 	:	val_out <= 4'h7bae;
         4'h8161 	:	val_out <= 4'h7bae;
         4'h8162 	:	val_out <= 4'h7bae;
         4'h8163 	:	val_out <= 4'h7bae;
         4'h8168 	:	val_out <= 4'h7b95;
         4'h8169 	:	val_out <= 4'h7b95;
         4'h816a 	:	val_out <= 4'h7b95;
         4'h816b 	:	val_out <= 4'h7b95;
         4'h8170 	:	val_out <= 4'h7b7c;
         4'h8171 	:	val_out <= 4'h7b7c;
         4'h8172 	:	val_out <= 4'h7b7c;
         4'h8173 	:	val_out <= 4'h7b7c;
         4'h8178 	:	val_out <= 4'h7b63;
         4'h8179 	:	val_out <= 4'h7b63;
         4'h817a 	:	val_out <= 4'h7b63;
         4'h817b 	:	val_out <= 4'h7b63;
         4'h8180 	:	val_out <= 4'h7b49;
         4'h8181 	:	val_out <= 4'h7b49;
         4'h8182 	:	val_out <= 4'h7b49;
         4'h8183 	:	val_out <= 4'h7b49;
         4'h8188 	:	val_out <= 4'h7b30;
         4'h8189 	:	val_out <= 4'h7b30;
         4'h818a 	:	val_out <= 4'h7b30;
         4'h818b 	:	val_out <= 4'h7b30;
         4'h8190 	:	val_out <= 4'h7b17;
         4'h8191 	:	val_out <= 4'h7b17;
         4'h8192 	:	val_out <= 4'h7b17;
         4'h8193 	:	val_out <= 4'h7b17;
         4'h8198 	:	val_out <= 4'h7afe;
         4'h8199 	:	val_out <= 4'h7afe;
         4'h819a 	:	val_out <= 4'h7afe;
         4'h819b 	:	val_out <= 4'h7afe;
         4'h81a0 	:	val_out <= 4'h7ae5;
         4'h81a1 	:	val_out <= 4'h7ae5;
         4'h81a2 	:	val_out <= 4'h7ae5;
         4'h81a3 	:	val_out <= 4'h7ae5;
         4'h81a8 	:	val_out <= 4'h7acc;
         4'h81a9 	:	val_out <= 4'h7acc;
         4'h81aa 	:	val_out <= 4'h7acc;
         4'h81ab 	:	val_out <= 4'h7acc;
         4'h81b0 	:	val_out <= 4'h7ab3;
         4'h81b1 	:	val_out <= 4'h7ab3;
         4'h81b2 	:	val_out <= 4'h7ab3;
         4'h81b3 	:	val_out <= 4'h7ab3;
         4'h81b8 	:	val_out <= 4'h7a9a;
         4'h81b9 	:	val_out <= 4'h7a9a;
         4'h81ba 	:	val_out <= 4'h7a9a;
         4'h81bb 	:	val_out <= 4'h7a9a;
         4'h81c0 	:	val_out <= 4'h7a80;
         4'h81c1 	:	val_out <= 4'h7a80;
         4'h81c2 	:	val_out <= 4'h7a80;
         4'h81c3 	:	val_out <= 4'h7a80;
         4'h81c8 	:	val_out <= 4'h7a67;
         4'h81c9 	:	val_out <= 4'h7a67;
         4'h81ca 	:	val_out <= 4'h7a67;
         4'h81cb 	:	val_out <= 4'h7a67;
         4'h81d0 	:	val_out <= 4'h7a4e;
         4'h81d1 	:	val_out <= 4'h7a4e;
         4'h81d2 	:	val_out <= 4'h7a4e;
         4'h81d3 	:	val_out <= 4'h7a4e;
         4'h81d8 	:	val_out <= 4'h7a35;
         4'h81d9 	:	val_out <= 4'h7a35;
         4'h81da 	:	val_out <= 4'h7a35;
         4'h81db 	:	val_out <= 4'h7a35;
         4'h81e0 	:	val_out <= 4'h7a1c;
         4'h81e1 	:	val_out <= 4'h7a1c;
         4'h81e2 	:	val_out <= 4'h7a1c;
         4'h81e3 	:	val_out <= 4'h7a1c;
         4'h81e8 	:	val_out <= 4'h7a03;
         4'h81e9 	:	val_out <= 4'h7a03;
         4'h81ea 	:	val_out <= 4'h7a03;
         4'h81eb 	:	val_out <= 4'h7a03;
         4'h81f0 	:	val_out <= 4'h79ea;
         4'h81f1 	:	val_out <= 4'h79ea;
         4'h81f2 	:	val_out <= 4'h79ea;
         4'h81f3 	:	val_out <= 4'h79ea;
         4'h81f8 	:	val_out <= 4'h79d1;
         4'h81f9 	:	val_out <= 4'h79d1;
         4'h81fa 	:	val_out <= 4'h79d1;
         4'h81fb 	:	val_out <= 4'h79d1;
         4'h8200 	:	val_out <= 4'h79b8;
         4'h8201 	:	val_out <= 4'h79b8;
         4'h8202 	:	val_out <= 4'h79b8;
         4'h8203 	:	val_out <= 4'h79b8;
         4'h8208 	:	val_out <= 4'h799f;
         4'h8209 	:	val_out <= 4'h799f;
         4'h820a 	:	val_out <= 4'h799f;
         4'h820b 	:	val_out <= 4'h799f;
         4'h8210 	:	val_out <= 4'h7985;
         4'h8211 	:	val_out <= 4'h7985;
         4'h8212 	:	val_out <= 4'h7985;
         4'h8213 	:	val_out <= 4'h7985;
         4'h8218 	:	val_out <= 4'h796c;
         4'h8219 	:	val_out <= 4'h796c;
         4'h821a 	:	val_out <= 4'h796c;
         4'h821b 	:	val_out <= 4'h796c;
         4'h8220 	:	val_out <= 4'h7953;
         4'h8221 	:	val_out <= 4'h7953;
         4'h8222 	:	val_out <= 4'h7953;
         4'h8223 	:	val_out <= 4'h7953;
         4'h8228 	:	val_out <= 4'h793a;
         4'h8229 	:	val_out <= 4'h793a;
         4'h822a 	:	val_out <= 4'h793a;
         4'h822b 	:	val_out <= 4'h793a;
         4'h8230 	:	val_out <= 4'h7921;
         4'h8231 	:	val_out <= 4'h7921;
         4'h8232 	:	val_out <= 4'h7921;
         4'h8233 	:	val_out <= 4'h7921;
         4'h8238 	:	val_out <= 4'h7908;
         4'h8239 	:	val_out <= 4'h7908;
         4'h823a 	:	val_out <= 4'h7908;
         4'h823b 	:	val_out <= 4'h7908;
         4'h8240 	:	val_out <= 4'h78ef;
         4'h8241 	:	val_out <= 4'h78ef;
         4'h8242 	:	val_out <= 4'h78ef;
         4'h8243 	:	val_out <= 4'h78ef;
         4'h8248 	:	val_out <= 4'h78d6;
         4'h8249 	:	val_out <= 4'h78d6;
         4'h824a 	:	val_out <= 4'h78d6;
         4'h824b 	:	val_out <= 4'h78d6;
         4'h8250 	:	val_out <= 4'h78bd;
         4'h8251 	:	val_out <= 4'h78bd;
         4'h8252 	:	val_out <= 4'h78bd;
         4'h8253 	:	val_out <= 4'h78bd;
         4'h8258 	:	val_out <= 4'h78a4;
         4'h8259 	:	val_out <= 4'h78a4;
         4'h825a 	:	val_out <= 4'h78a4;
         4'h825b 	:	val_out <= 4'h78a4;
         4'h8260 	:	val_out <= 4'h788a;
         4'h8261 	:	val_out <= 4'h788a;
         4'h8262 	:	val_out <= 4'h788a;
         4'h8263 	:	val_out <= 4'h788a;
         4'h8268 	:	val_out <= 4'h7871;
         4'h8269 	:	val_out <= 4'h7871;
         4'h826a 	:	val_out <= 4'h7871;
         4'h826b 	:	val_out <= 4'h7871;
         4'h8270 	:	val_out <= 4'h7858;
         4'h8271 	:	val_out <= 4'h7858;
         4'h8272 	:	val_out <= 4'h7858;
         4'h8273 	:	val_out <= 4'h7858;
         4'h8278 	:	val_out <= 4'h783f;
         4'h8279 	:	val_out <= 4'h783f;
         4'h827a 	:	val_out <= 4'h783f;
         4'h827b 	:	val_out <= 4'h783f;
         4'h8280 	:	val_out <= 4'h7826;
         4'h8281 	:	val_out <= 4'h7826;
         4'h8282 	:	val_out <= 4'h7826;
         4'h8283 	:	val_out <= 4'h7826;
         4'h8288 	:	val_out <= 4'h780d;
         4'h8289 	:	val_out <= 4'h780d;
         4'h828a 	:	val_out <= 4'h780d;
         4'h828b 	:	val_out <= 4'h780d;
         4'h8290 	:	val_out <= 4'h77f4;
         4'h8291 	:	val_out <= 4'h77f4;
         4'h8292 	:	val_out <= 4'h77f4;
         4'h8293 	:	val_out <= 4'h77f4;
         4'h8298 	:	val_out <= 4'h77db;
         4'h8299 	:	val_out <= 4'h77db;
         4'h829a 	:	val_out <= 4'h77db;
         4'h829b 	:	val_out <= 4'h77db;
         4'h82a0 	:	val_out <= 4'h77c2;
         4'h82a1 	:	val_out <= 4'h77c2;
         4'h82a2 	:	val_out <= 4'h77c2;
         4'h82a3 	:	val_out <= 4'h77c2;
         4'h82a8 	:	val_out <= 4'h77a9;
         4'h82a9 	:	val_out <= 4'h77a9;
         4'h82aa 	:	val_out <= 4'h77a9;
         4'h82ab 	:	val_out <= 4'h77a9;
         4'h82b0 	:	val_out <= 4'h7790;
         4'h82b1 	:	val_out <= 4'h7790;
         4'h82b2 	:	val_out <= 4'h7790;
         4'h82b3 	:	val_out <= 4'h7790;
         4'h82b8 	:	val_out <= 4'h7777;
         4'h82b9 	:	val_out <= 4'h7777;
         4'h82ba 	:	val_out <= 4'h7777;
         4'h82bb 	:	val_out <= 4'h7777;
         4'h82c0 	:	val_out <= 4'h775d;
         4'h82c1 	:	val_out <= 4'h775d;
         4'h82c2 	:	val_out <= 4'h775d;
         4'h82c3 	:	val_out <= 4'h775d;
         4'h82c8 	:	val_out <= 4'h7744;
         4'h82c9 	:	val_out <= 4'h7744;
         4'h82ca 	:	val_out <= 4'h7744;
         4'h82cb 	:	val_out <= 4'h7744;
         4'h82d0 	:	val_out <= 4'h772b;
         4'h82d1 	:	val_out <= 4'h772b;
         4'h82d2 	:	val_out <= 4'h772b;
         4'h82d3 	:	val_out <= 4'h772b;
         4'h82d8 	:	val_out <= 4'h7712;
         4'h82d9 	:	val_out <= 4'h7712;
         4'h82da 	:	val_out <= 4'h7712;
         4'h82db 	:	val_out <= 4'h7712;
         4'h82e0 	:	val_out <= 4'h76f9;
         4'h82e1 	:	val_out <= 4'h76f9;
         4'h82e2 	:	val_out <= 4'h76f9;
         4'h82e3 	:	val_out <= 4'h76f9;
         4'h82e8 	:	val_out <= 4'h76e0;
         4'h82e9 	:	val_out <= 4'h76e0;
         4'h82ea 	:	val_out <= 4'h76e0;
         4'h82eb 	:	val_out <= 4'h76e0;
         4'h82f0 	:	val_out <= 4'h76c7;
         4'h82f1 	:	val_out <= 4'h76c7;
         4'h82f2 	:	val_out <= 4'h76c7;
         4'h82f3 	:	val_out <= 4'h76c7;
         4'h82f8 	:	val_out <= 4'h76ae;
         4'h82f9 	:	val_out <= 4'h76ae;
         4'h82fa 	:	val_out <= 4'h76ae;
         4'h82fb 	:	val_out <= 4'h76ae;
         4'h8300 	:	val_out <= 4'h7695;
         4'h8301 	:	val_out <= 4'h7695;
         4'h8302 	:	val_out <= 4'h7695;
         4'h8303 	:	val_out <= 4'h7695;
         4'h8308 	:	val_out <= 4'h767c;
         4'h8309 	:	val_out <= 4'h767c;
         4'h830a 	:	val_out <= 4'h767c;
         4'h830b 	:	val_out <= 4'h767c;
         4'h8310 	:	val_out <= 4'h7663;
         4'h8311 	:	val_out <= 4'h7663;
         4'h8312 	:	val_out <= 4'h7663;
         4'h8313 	:	val_out <= 4'h7663;
         4'h8318 	:	val_out <= 4'h764a;
         4'h8319 	:	val_out <= 4'h764a;
         4'h831a 	:	val_out <= 4'h764a;
         4'h831b 	:	val_out <= 4'h764a;
         4'h8320 	:	val_out <= 4'h7631;
         4'h8321 	:	val_out <= 4'h7631;
         4'h8322 	:	val_out <= 4'h7631;
         4'h8323 	:	val_out <= 4'h7631;
         4'h8328 	:	val_out <= 4'h7618;
         4'h8329 	:	val_out <= 4'h7618;
         4'h832a 	:	val_out <= 4'h7618;
         4'h832b 	:	val_out <= 4'h7618;
         4'h8330 	:	val_out <= 4'h75ff;
         4'h8331 	:	val_out <= 4'h75ff;
         4'h8332 	:	val_out <= 4'h75ff;
         4'h8333 	:	val_out <= 4'h75ff;
         4'h8338 	:	val_out <= 4'h75e6;
         4'h8339 	:	val_out <= 4'h75e6;
         4'h833a 	:	val_out <= 4'h75e6;
         4'h833b 	:	val_out <= 4'h75e6;
         4'h8340 	:	val_out <= 4'h75cc;
         4'h8341 	:	val_out <= 4'h75cc;
         4'h8342 	:	val_out <= 4'h75cc;
         4'h8343 	:	val_out <= 4'h75cc;
         4'h8348 	:	val_out <= 4'h75b3;
         4'h8349 	:	val_out <= 4'h75b3;
         4'h834a 	:	val_out <= 4'h75b3;
         4'h834b 	:	val_out <= 4'h75b3;
         4'h8350 	:	val_out <= 4'h759a;
         4'h8351 	:	val_out <= 4'h759a;
         4'h8352 	:	val_out <= 4'h759a;
         4'h8353 	:	val_out <= 4'h759a;
         4'h8358 	:	val_out <= 4'h7581;
         4'h8359 	:	val_out <= 4'h7581;
         4'h835a 	:	val_out <= 4'h7581;
         4'h835b 	:	val_out <= 4'h7581;
         4'h8360 	:	val_out <= 4'h7568;
         4'h8361 	:	val_out <= 4'h7568;
         4'h8362 	:	val_out <= 4'h7568;
         4'h8363 	:	val_out <= 4'h7568;
         4'h8368 	:	val_out <= 4'h754f;
         4'h8369 	:	val_out <= 4'h754f;
         4'h836a 	:	val_out <= 4'h754f;
         4'h836b 	:	val_out <= 4'h754f;
         4'h8370 	:	val_out <= 4'h7536;
         4'h8371 	:	val_out <= 4'h7536;
         4'h8372 	:	val_out <= 4'h7536;
         4'h8373 	:	val_out <= 4'h7536;
         4'h8378 	:	val_out <= 4'h751d;
         4'h8379 	:	val_out <= 4'h751d;
         4'h837a 	:	val_out <= 4'h751d;
         4'h837b 	:	val_out <= 4'h751d;
         4'h8380 	:	val_out <= 4'h7504;
         4'h8381 	:	val_out <= 4'h7504;
         4'h8382 	:	val_out <= 4'h7504;
         4'h8383 	:	val_out <= 4'h7504;
         4'h8388 	:	val_out <= 4'h74eb;
         4'h8389 	:	val_out <= 4'h74eb;
         4'h838a 	:	val_out <= 4'h74eb;
         4'h838b 	:	val_out <= 4'h74eb;
         4'h8390 	:	val_out <= 4'h74d2;
         4'h8391 	:	val_out <= 4'h74d2;
         4'h8392 	:	val_out <= 4'h74d2;
         4'h8393 	:	val_out <= 4'h74d2;
         4'h8398 	:	val_out <= 4'h74b9;
         4'h8399 	:	val_out <= 4'h74b9;
         4'h839a 	:	val_out <= 4'h74b9;
         4'h839b 	:	val_out <= 4'h74b9;
         4'h83a0 	:	val_out <= 4'h74a0;
         4'h83a1 	:	val_out <= 4'h74a0;
         4'h83a2 	:	val_out <= 4'h74a0;
         4'h83a3 	:	val_out <= 4'h74a0;
         4'h83a8 	:	val_out <= 4'h7487;
         4'h83a9 	:	val_out <= 4'h7487;
         4'h83aa 	:	val_out <= 4'h7487;
         4'h83ab 	:	val_out <= 4'h7487;
         4'h83b0 	:	val_out <= 4'h746e;
         4'h83b1 	:	val_out <= 4'h746e;
         4'h83b2 	:	val_out <= 4'h746e;
         4'h83b3 	:	val_out <= 4'h746e;
         4'h83b8 	:	val_out <= 4'h7455;
         4'h83b9 	:	val_out <= 4'h7455;
         4'h83ba 	:	val_out <= 4'h7455;
         4'h83bb 	:	val_out <= 4'h7455;
         4'h83c0 	:	val_out <= 4'h743c;
         4'h83c1 	:	val_out <= 4'h743c;
         4'h83c2 	:	val_out <= 4'h743c;
         4'h83c3 	:	val_out <= 4'h743c;
         4'h83c8 	:	val_out <= 4'h7423;
         4'h83c9 	:	val_out <= 4'h7423;
         4'h83ca 	:	val_out <= 4'h7423;
         4'h83cb 	:	val_out <= 4'h7423;
         4'h83d0 	:	val_out <= 4'h740a;
         4'h83d1 	:	val_out <= 4'h740a;
         4'h83d2 	:	val_out <= 4'h740a;
         4'h83d3 	:	val_out <= 4'h740a;
         4'h83d8 	:	val_out <= 4'h73f1;
         4'h83d9 	:	val_out <= 4'h73f1;
         4'h83da 	:	val_out <= 4'h73f1;
         4'h83db 	:	val_out <= 4'h73f1;
         4'h83e0 	:	val_out <= 4'h73d8;
         4'h83e1 	:	val_out <= 4'h73d8;
         4'h83e2 	:	val_out <= 4'h73d8;
         4'h83e3 	:	val_out <= 4'h73d8;
         4'h83e8 	:	val_out <= 4'h73bf;
         4'h83e9 	:	val_out <= 4'h73bf;
         4'h83ea 	:	val_out <= 4'h73bf;
         4'h83eb 	:	val_out <= 4'h73bf;
         4'h83f0 	:	val_out <= 4'h73a6;
         4'h83f1 	:	val_out <= 4'h73a6;
         4'h83f2 	:	val_out <= 4'h73a6;
         4'h83f3 	:	val_out <= 4'h73a6;
         4'h83f8 	:	val_out <= 4'h738d;
         4'h83f9 	:	val_out <= 4'h738d;
         4'h83fa 	:	val_out <= 4'h738d;
         4'h83fb 	:	val_out <= 4'h738d;
         4'h8400 	:	val_out <= 4'h7374;
         4'h8401 	:	val_out <= 4'h7374;
         4'h8402 	:	val_out <= 4'h7374;
         4'h8403 	:	val_out <= 4'h7374;
         4'h8408 	:	val_out <= 4'h735b;
         4'h8409 	:	val_out <= 4'h735b;
         4'h840a 	:	val_out <= 4'h735b;
         4'h840b 	:	val_out <= 4'h735b;
         4'h8410 	:	val_out <= 4'h7342;
         4'h8411 	:	val_out <= 4'h7342;
         4'h8412 	:	val_out <= 4'h7342;
         4'h8413 	:	val_out <= 4'h7342;
         4'h8418 	:	val_out <= 4'h7329;
         4'h8419 	:	val_out <= 4'h7329;
         4'h841a 	:	val_out <= 4'h7329;
         4'h841b 	:	val_out <= 4'h7329;
         4'h8420 	:	val_out <= 4'h7310;
         4'h8421 	:	val_out <= 4'h7310;
         4'h8422 	:	val_out <= 4'h7310;
         4'h8423 	:	val_out <= 4'h7310;
         4'h8428 	:	val_out <= 4'h72f7;
         4'h8429 	:	val_out <= 4'h72f7;
         4'h842a 	:	val_out <= 4'h72f7;
         4'h842b 	:	val_out <= 4'h72f7;
         4'h8430 	:	val_out <= 4'h72de;
         4'h8431 	:	val_out <= 4'h72de;
         4'h8432 	:	val_out <= 4'h72de;
         4'h8433 	:	val_out <= 4'h72de;
         4'h8438 	:	val_out <= 4'h72c5;
         4'h8439 	:	val_out <= 4'h72c5;
         4'h843a 	:	val_out <= 4'h72c5;
         4'h843b 	:	val_out <= 4'h72c5;
         4'h8440 	:	val_out <= 4'h72ac;
         4'h8441 	:	val_out <= 4'h72ac;
         4'h8442 	:	val_out <= 4'h72ac;
         4'h8443 	:	val_out <= 4'h72ac;
         4'h8448 	:	val_out <= 4'h7293;
         4'h8449 	:	val_out <= 4'h7293;
         4'h844a 	:	val_out <= 4'h7293;
         4'h844b 	:	val_out <= 4'h7293;
         4'h8450 	:	val_out <= 4'h727a;
         4'h8451 	:	val_out <= 4'h727a;
         4'h8452 	:	val_out <= 4'h727a;
         4'h8453 	:	val_out <= 4'h727a;
         4'h8458 	:	val_out <= 4'h7261;
         4'h8459 	:	val_out <= 4'h7261;
         4'h845a 	:	val_out <= 4'h7261;
         4'h845b 	:	val_out <= 4'h7261;
         4'h8460 	:	val_out <= 4'h7248;
         4'h8461 	:	val_out <= 4'h7248;
         4'h8462 	:	val_out <= 4'h7248;
         4'h8463 	:	val_out <= 4'h7248;
         4'h8468 	:	val_out <= 4'h722f;
         4'h8469 	:	val_out <= 4'h722f;
         4'h846a 	:	val_out <= 4'h722f;
         4'h846b 	:	val_out <= 4'h722f;
         4'h8470 	:	val_out <= 4'h7216;
         4'h8471 	:	val_out <= 4'h7216;
         4'h8472 	:	val_out <= 4'h7216;
         4'h8473 	:	val_out <= 4'h7216;
         4'h8478 	:	val_out <= 4'h71fd;
         4'h8479 	:	val_out <= 4'h71fd;
         4'h847a 	:	val_out <= 4'h71fd;
         4'h847b 	:	val_out <= 4'h71fd;
         4'h8480 	:	val_out <= 4'h71e4;
         4'h8481 	:	val_out <= 4'h71e4;
         4'h8482 	:	val_out <= 4'h71e4;
         4'h8483 	:	val_out <= 4'h71e4;
         4'h8488 	:	val_out <= 4'h71cb;
         4'h8489 	:	val_out <= 4'h71cb;
         4'h848a 	:	val_out <= 4'h71cb;
         4'h848b 	:	val_out <= 4'h71cb;
         4'h8490 	:	val_out <= 4'h71b2;
         4'h8491 	:	val_out <= 4'h71b2;
         4'h8492 	:	val_out <= 4'h71b2;
         4'h8493 	:	val_out <= 4'h71b2;
         4'h8498 	:	val_out <= 4'h7199;
         4'h8499 	:	val_out <= 4'h7199;
         4'h849a 	:	val_out <= 4'h7199;
         4'h849b 	:	val_out <= 4'h7199;
         4'h84a0 	:	val_out <= 4'h7180;
         4'h84a1 	:	val_out <= 4'h7180;
         4'h84a2 	:	val_out <= 4'h7180;
         4'h84a3 	:	val_out <= 4'h7180;
         4'h84a8 	:	val_out <= 4'h7167;
         4'h84a9 	:	val_out <= 4'h7167;
         4'h84aa 	:	val_out <= 4'h7167;
         4'h84ab 	:	val_out <= 4'h7167;
         4'h84b0 	:	val_out <= 4'h714e;
         4'h84b1 	:	val_out <= 4'h714e;
         4'h84b2 	:	val_out <= 4'h714e;
         4'h84b3 	:	val_out <= 4'h714e;
         4'h84b8 	:	val_out <= 4'h7135;
         4'h84b9 	:	val_out <= 4'h7135;
         4'h84ba 	:	val_out <= 4'h7135;
         4'h84bb 	:	val_out <= 4'h7135;
         4'h84c0 	:	val_out <= 4'h711c;
         4'h84c1 	:	val_out <= 4'h711c;
         4'h84c2 	:	val_out <= 4'h711c;
         4'h84c3 	:	val_out <= 4'h711c;
         4'h84c8 	:	val_out <= 4'h7103;
         4'h84c9 	:	val_out <= 4'h7103;
         4'h84ca 	:	val_out <= 4'h7103;
         4'h84cb 	:	val_out <= 4'h7103;
         4'h84d0 	:	val_out <= 4'h70ea;
         4'h84d1 	:	val_out <= 4'h70ea;
         4'h84d2 	:	val_out <= 4'h70ea;
         4'h84d3 	:	val_out <= 4'h70ea;
         4'h84d8 	:	val_out <= 4'h70d1;
         4'h84d9 	:	val_out <= 4'h70d1;
         4'h84da 	:	val_out <= 4'h70d1;
         4'h84db 	:	val_out <= 4'h70d1;
         4'h84e0 	:	val_out <= 4'h70b8;
         4'h84e1 	:	val_out <= 4'h70b8;
         4'h84e2 	:	val_out <= 4'h70b8;
         4'h84e3 	:	val_out <= 4'h70b8;
         4'h84e8 	:	val_out <= 4'h709f;
         4'h84e9 	:	val_out <= 4'h709f;
         4'h84ea 	:	val_out <= 4'h709f;
         4'h84eb 	:	val_out <= 4'h709f;
         4'h84f0 	:	val_out <= 4'h7086;
         4'h84f1 	:	val_out <= 4'h7086;
         4'h84f2 	:	val_out <= 4'h7086;
         4'h84f3 	:	val_out <= 4'h7086;
         4'h84f8 	:	val_out <= 4'h706d;
         4'h84f9 	:	val_out <= 4'h706d;
         4'h84fa 	:	val_out <= 4'h706d;
         4'h84fb 	:	val_out <= 4'h706d;
         4'h8500 	:	val_out <= 4'h7054;
         4'h8501 	:	val_out <= 4'h7054;
         4'h8502 	:	val_out <= 4'h7054;
         4'h8503 	:	val_out <= 4'h7054;
         4'h8508 	:	val_out <= 4'h703b;
         4'h8509 	:	val_out <= 4'h703b;
         4'h850a 	:	val_out <= 4'h703b;
         4'h850b 	:	val_out <= 4'h703b;
         4'h8510 	:	val_out <= 4'h7022;
         4'h8511 	:	val_out <= 4'h7022;
         4'h8512 	:	val_out <= 4'h7022;
         4'h8513 	:	val_out <= 4'h7022;
         4'h8518 	:	val_out <= 4'h700a;
         4'h8519 	:	val_out <= 4'h700a;
         4'h851a 	:	val_out <= 4'h700a;
         4'h851b 	:	val_out <= 4'h700a;
         4'h8520 	:	val_out <= 4'h6ff1;
         4'h8521 	:	val_out <= 4'h6ff1;
         4'h8522 	:	val_out <= 4'h6ff1;
         4'h8523 	:	val_out <= 4'h6ff1;
         4'h8528 	:	val_out <= 4'h6fd8;
         4'h8529 	:	val_out <= 4'h6fd8;
         4'h852a 	:	val_out <= 4'h6fd8;
         4'h852b 	:	val_out <= 4'h6fd8;
         4'h8530 	:	val_out <= 4'h6fbf;
         4'h8531 	:	val_out <= 4'h6fbf;
         4'h8532 	:	val_out <= 4'h6fbf;
         4'h8533 	:	val_out <= 4'h6fbf;
         4'h8538 	:	val_out <= 4'h6fa6;
         4'h8539 	:	val_out <= 4'h6fa6;
         4'h853a 	:	val_out <= 4'h6fa6;
         4'h853b 	:	val_out <= 4'h6fa6;
         4'h8540 	:	val_out <= 4'h6f8d;
         4'h8541 	:	val_out <= 4'h6f8d;
         4'h8542 	:	val_out <= 4'h6f8d;
         4'h8543 	:	val_out <= 4'h6f8d;
         4'h8548 	:	val_out <= 4'h6f74;
         4'h8549 	:	val_out <= 4'h6f74;
         4'h854a 	:	val_out <= 4'h6f74;
         4'h854b 	:	val_out <= 4'h6f74;
         4'h8550 	:	val_out <= 4'h6f5b;
         4'h8551 	:	val_out <= 4'h6f5b;
         4'h8552 	:	val_out <= 4'h6f5b;
         4'h8553 	:	val_out <= 4'h6f5b;
         4'h8558 	:	val_out <= 4'h6f42;
         4'h8559 	:	val_out <= 4'h6f42;
         4'h855a 	:	val_out <= 4'h6f42;
         4'h855b 	:	val_out <= 4'h6f42;
         4'h8560 	:	val_out <= 4'h6f29;
         4'h8561 	:	val_out <= 4'h6f29;
         4'h8562 	:	val_out <= 4'h6f29;
         4'h8563 	:	val_out <= 4'h6f29;
         4'h8568 	:	val_out <= 4'h6f10;
         4'h8569 	:	val_out <= 4'h6f10;
         4'h856a 	:	val_out <= 4'h6f10;
         4'h856b 	:	val_out <= 4'h6f10;
         4'h8570 	:	val_out <= 4'h6ef7;
         4'h8571 	:	val_out <= 4'h6ef7;
         4'h8572 	:	val_out <= 4'h6ef7;
         4'h8573 	:	val_out <= 4'h6ef7;
         4'h8578 	:	val_out <= 4'h6ede;
         4'h8579 	:	val_out <= 4'h6ede;
         4'h857a 	:	val_out <= 4'h6ede;
         4'h857b 	:	val_out <= 4'h6ede;
         4'h8580 	:	val_out <= 4'h6ec6;
         4'h8581 	:	val_out <= 4'h6ec6;
         4'h8582 	:	val_out <= 4'h6ec6;
         4'h8583 	:	val_out <= 4'h6ec6;
         4'h8588 	:	val_out <= 4'h6ead;
         4'h8589 	:	val_out <= 4'h6ead;
         4'h858a 	:	val_out <= 4'h6ead;
         4'h858b 	:	val_out <= 4'h6ead;
         4'h8590 	:	val_out <= 4'h6e94;
         4'h8591 	:	val_out <= 4'h6e94;
         4'h8592 	:	val_out <= 4'h6e94;
         4'h8593 	:	val_out <= 4'h6e94;
         4'h8598 	:	val_out <= 4'h6e7b;
         4'h8599 	:	val_out <= 4'h6e7b;
         4'h859a 	:	val_out <= 4'h6e7b;
         4'h859b 	:	val_out <= 4'h6e7b;
         4'h85a0 	:	val_out <= 4'h6e62;
         4'h85a1 	:	val_out <= 4'h6e62;
         4'h85a2 	:	val_out <= 4'h6e62;
         4'h85a3 	:	val_out <= 4'h6e62;
         4'h85a8 	:	val_out <= 4'h6e49;
         4'h85a9 	:	val_out <= 4'h6e49;
         4'h85aa 	:	val_out <= 4'h6e49;
         4'h85ab 	:	val_out <= 4'h6e49;
         4'h85b0 	:	val_out <= 4'h6e30;
         4'h85b1 	:	val_out <= 4'h6e30;
         4'h85b2 	:	val_out <= 4'h6e30;
         4'h85b3 	:	val_out <= 4'h6e30;
         4'h85b8 	:	val_out <= 4'h6e17;
         4'h85b9 	:	val_out <= 4'h6e17;
         4'h85ba 	:	val_out <= 4'h6e17;
         4'h85bb 	:	val_out <= 4'h6e17;
         4'h85c0 	:	val_out <= 4'h6dfe;
         4'h85c1 	:	val_out <= 4'h6dfe;
         4'h85c2 	:	val_out <= 4'h6dfe;
         4'h85c3 	:	val_out <= 4'h6dfe;
         4'h85c8 	:	val_out <= 4'h6de6;
         4'h85c9 	:	val_out <= 4'h6de6;
         4'h85ca 	:	val_out <= 4'h6de6;
         4'h85cb 	:	val_out <= 4'h6de6;
         4'h85d0 	:	val_out <= 4'h6dcd;
         4'h85d1 	:	val_out <= 4'h6dcd;
         4'h85d2 	:	val_out <= 4'h6dcd;
         4'h85d3 	:	val_out <= 4'h6dcd;
         4'h85d8 	:	val_out <= 4'h6db4;
         4'h85d9 	:	val_out <= 4'h6db4;
         4'h85da 	:	val_out <= 4'h6db4;
         4'h85db 	:	val_out <= 4'h6db4;
         4'h85e0 	:	val_out <= 4'h6d9b;
         4'h85e1 	:	val_out <= 4'h6d9b;
         4'h85e2 	:	val_out <= 4'h6d9b;
         4'h85e3 	:	val_out <= 4'h6d9b;
         4'h85e8 	:	val_out <= 4'h6d82;
         4'h85e9 	:	val_out <= 4'h6d82;
         4'h85ea 	:	val_out <= 4'h6d82;
         4'h85eb 	:	val_out <= 4'h6d82;
         4'h85f0 	:	val_out <= 4'h6d69;
         4'h85f1 	:	val_out <= 4'h6d69;
         4'h85f2 	:	val_out <= 4'h6d69;
         4'h85f3 	:	val_out <= 4'h6d69;
         4'h85f8 	:	val_out <= 4'h6d50;
         4'h85f9 	:	val_out <= 4'h6d50;
         4'h85fa 	:	val_out <= 4'h6d50;
         4'h85fb 	:	val_out <= 4'h6d50;
         4'h8600 	:	val_out <= 4'h6d37;
         4'h8601 	:	val_out <= 4'h6d37;
         4'h8602 	:	val_out <= 4'h6d37;
         4'h8603 	:	val_out <= 4'h6d37;
         4'h8608 	:	val_out <= 4'h6d1f;
         4'h8609 	:	val_out <= 4'h6d1f;
         4'h860a 	:	val_out <= 4'h6d1f;
         4'h860b 	:	val_out <= 4'h6d1f;
         4'h8610 	:	val_out <= 4'h6d06;
         4'h8611 	:	val_out <= 4'h6d06;
         4'h8612 	:	val_out <= 4'h6d06;
         4'h8613 	:	val_out <= 4'h6d06;
         4'h8618 	:	val_out <= 4'h6ced;
         4'h8619 	:	val_out <= 4'h6ced;
         4'h861a 	:	val_out <= 4'h6ced;
         4'h861b 	:	val_out <= 4'h6ced;
         4'h8620 	:	val_out <= 4'h6cd4;
         4'h8621 	:	val_out <= 4'h6cd4;
         4'h8622 	:	val_out <= 4'h6cd4;
         4'h8623 	:	val_out <= 4'h6cd4;
         4'h8628 	:	val_out <= 4'h6cbb;
         4'h8629 	:	val_out <= 4'h6cbb;
         4'h862a 	:	val_out <= 4'h6cbb;
         4'h862b 	:	val_out <= 4'h6cbb;
         4'h8630 	:	val_out <= 4'h6ca2;
         4'h8631 	:	val_out <= 4'h6ca2;
         4'h8632 	:	val_out <= 4'h6ca2;
         4'h8633 	:	val_out <= 4'h6ca2;
         4'h8638 	:	val_out <= 4'h6c89;
         4'h8639 	:	val_out <= 4'h6c89;
         4'h863a 	:	val_out <= 4'h6c89;
         4'h863b 	:	val_out <= 4'h6c89;
         4'h8640 	:	val_out <= 4'h6c71;
         4'h8641 	:	val_out <= 4'h6c71;
         4'h8642 	:	val_out <= 4'h6c71;
         4'h8643 	:	val_out <= 4'h6c71;
         4'h8648 	:	val_out <= 4'h6c58;
         4'h8649 	:	val_out <= 4'h6c58;
         4'h864a 	:	val_out <= 4'h6c58;
         4'h864b 	:	val_out <= 4'h6c58;
         4'h8650 	:	val_out <= 4'h6c3f;
         4'h8651 	:	val_out <= 4'h6c3f;
         4'h8652 	:	val_out <= 4'h6c3f;
         4'h8653 	:	val_out <= 4'h6c3f;
         4'h8658 	:	val_out <= 4'h6c26;
         4'h8659 	:	val_out <= 4'h6c26;
         4'h865a 	:	val_out <= 4'h6c26;
         4'h865b 	:	val_out <= 4'h6c26;
         4'h8660 	:	val_out <= 4'h6c0d;
         4'h8661 	:	val_out <= 4'h6c0d;
         4'h8662 	:	val_out <= 4'h6c0d;
         4'h8663 	:	val_out <= 4'h6c0d;
         4'h8668 	:	val_out <= 4'h6bf4;
         4'h8669 	:	val_out <= 4'h6bf4;
         4'h866a 	:	val_out <= 4'h6bf4;
         4'h866b 	:	val_out <= 4'h6bf4;
         4'h8670 	:	val_out <= 4'h6bdc;
         4'h8671 	:	val_out <= 4'h6bdc;
         4'h8672 	:	val_out <= 4'h6bdc;
         4'h8673 	:	val_out <= 4'h6bdc;
         4'h8678 	:	val_out <= 4'h6bc3;
         4'h8679 	:	val_out <= 4'h6bc3;
         4'h867a 	:	val_out <= 4'h6bc3;
         4'h867b 	:	val_out <= 4'h6bc3;
         4'h8680 	:	val_out <= 4'h6baa;
         4'h8681 	:	val_out <= 4'h6baa;
         4'h8682 	:	val_out <= 4'h6baa;
         4'h8683 	:	val_out <= 4'h6baa;
         4'h8688 	:	val_out <= 4'h6b91;
         4'h8689 	:	val_out <= 4'h6b91;
         4'h868a 	:	val_out <= 4'h6b91;
         4'h868b 	:	val_out <= 4'h6b91;
         4'h8690 	:	val_out <= 4'h6b78;
         4'h8691 	:	val_out <= 4'h6b78;
         4'h8692 	:	val_out <= 4'h6b78;
         4'h8693 	:	val_out <= 4'h6b78;
         4'h8698 	:	val_out <= 4'h6b60;
         4'h8699 	:	val_out <= 4'h6b60;
         4'h869a 	:	val_out <= 4'h6b60;
         4'h869b 	:	val_out <= 4'h6b60;
         4'h86a0 	:	val_out <= 4'h6b47;
         4'h86a1 	:	val_out <= 4'h6b47;
         4'h86a2 	:	val_out <= 4'h6b47;
         4'h86a3 	:	val_out <= 4'h6b47;
         4'h86a8 	:	val_out <= 4'h6b2e;
         4'h86a9 	:	val_out <= 4'h6b2e;
         4'h86aa 	:	val_out <= 4'h6b2e;
         4'h86ab 	:	val_out <= 4'h6b2e;
         4'h86b0 	:	val_out <= 4'h6b15;
         4'h86b1 	:	val_out <= 4'h6b15;
         4'h86b2 	:	val_out <= 4'h6b15;
         4'h86b3 	:	val_out <= 4'h6b15;
         4'h86b8 	:	val_out <= 4'h6afc;
         4'h86b9 	:	val_out <= 4'h6afc;
         4'h86ba 	:	val_out <= 4'h6afc;
         4'h86bb 	:	val_out <= 4'h6afc;
         4'h86c0 	:	val_out <= 4'h6ae4;
         4'h86c1 	:	val_out <= 4'h6ae4;
         4'h86c2 	:	val_out <= 4'h6ae4;
         4'h86c3 	:	val_out <= 4'h6ae4;
         4'h86c8 	:	val_out <= 4'h6acb;
         4'h86c9 	:	val_out <= 4'h6acb;
         4'h86ca 	:	val_out <= 4'h6acb;
         4'h86cb 	:	val_out <= 4'h6acb;
         4'h86d0 	:	val_out <= 4'h6ab2;
         4'h86d1 	:	val_out <= 4'h6ab2;
         4'h86d2 	:	val_out <= 4'h6ab2;
         4'h86d3 	:	val_out <= 4'h6ab2;
         4'h86d8 	:	val_out <= 4'h6a99;
         4'h86d9 	:	val_out <= 4'h6a99;
         4'h86da 	:	val_out <= 4'h6a99;
         4'h86db 	:	val_out <= 4'h6a99;
         4'h86e0 	:	val_out <= 4'h6a80;
         4'h86e1 	:	val_out <= 4'h6a80;
         4'h86e2 	:	val_out <= 4'h6a80;
         4'h86e3 	:	val_out <= 4'h6a80;
         4'h86e8 	:	val_out <= 4'h6a68;
         4'h86e9 	:	val_out <= 4'h6a68;
         4'h86ea 	:	val_out <= 4'h6a68;
         4'h86eb 	:	val_out <= 4'h6a68;
         4'h86f0 	:	val_out <= 4'h6a4f;
         4'h86f1 	:	val_out <= 4'h6a4f;
         4'h86f2 	:	val_out <= 4'h6a4f;
         4'h86f3 	:	val_out <= 4'h6a4f;
         4'h86f8 	:	val_out <= 4'h6a36;
         4'h86f9 	:	val_out <= 4'h6a36;
         4'h86fa 	:	val_out <= 4'h6a36;
         4'h86fb 	:	val_out <= 4'h6a36;
         4'h8700 	:	val_out <= 4'h6a1d;
         4'h8701 	:	val_out <= 4'h6a1d;
         4'h8702 	:	val_out <= 4'h6a1d;
         4'h8703 	:	val_out <= 4'h6a1d;
         4'h8708 	:	val_out <= 4'h6a05;
         4'h8709 	:	val_out <= 4'h6a05;
         4'h870a 	:	val_out <= 4'h6a05;
         4'h870b 	:	val_out <= 4'h6a05;
         4'h8710 	:	val_out <= 4'h69ec;
         4'h8711 	:	val_out <= 4'h69ec;
         4'h8712 	:	val_out <= 4'h69ec;
         4'h8713 	:	val_out <= 4'h69ec;
         4'h8718 	:	val_out <= 4'h69d3;
         4'h8719 	:	val_out <= 4'h69d3;
         4'h871a 	:	val_out <= 4'h69d3;
         4'h871b 	:	val_out <= 4'h69d3;
         4'h8720 	:	val_out <= 4'h69ba;
         4'h8721 	:	val_out <= 4'h69ba;
         4'h8722 	:	val_out <= 4'h69ba;
         4'h8723 	:	val_out <= 4'h69ba;
         4'h8728 	:	val_out <= 4'h69a2;
         4'h8729 	:	val_out <= 4'h69a2;
         4'h872a 	:	val_out <= 4'h69a2;
         4'h872b 	:	val_out <= 4'h69a2;
         4'h8730 	:	val_out <= 4'h6989;
         4'h8731 	:	val_out <= 4'h6989;
         4'h8732 	:	val_out <= 4'h6989;
         4'h8733 	:	val_out <= 4'h6989;
         4'h8738 	:	val_out <= 4'h6970;
         4'h8739 	:	val_out <= 4'h6970;
         4'h873a 	:	val_out <= 4'h6970;
         4'h873b 	:	val_out <= 4'h6970;
         4'h8740 	:	val_out <= 4'h6957;
         4'h8741 	:	val_out <= 4'h6957;
         4'h8742 	:	val_out <= 4'h6957;
         4'h8743 	:	val_out <= 4'h6957;
         4'h8748 	:	val_out <= 4'h693f;
         4'h8749 	:	val_out <= 4'h693f;
         4'h874a 	:	val_out <= 4'h693f;
         4'h874b 	:	val_out <= 4'h693f;
         4'h8750 	:	val_out <= 4'h6926;
         4'h8751 	:	val_out <= 4'h6926;
         4'h8752 	:	val_out <= 4'h6926;
         4'h8753 	:	val_out <= 4'h6926;
         4'h8758 	:	val_out <= 4'h690d;
         4'h8759 	:	val_out <= 4'h690d;
         4'h875a 	:	val_out <= 4'h690d;
         4'h875b 	:	val_out <= 4'h690d;
         4'h8760 	:	val_out <= 4'h68f5;
         4'h8761 	:	val_out <= 4'h68f5;
         4'h8762 	:	val_out <= 4'h68f5;
         4'h8763 	:	val_out <= 4'h68f5;
         4'h8768 	:	val_out <= 4'h68dc;
         4'h8769 	:	val_out <= 4'h68dc;
         4'h876a 	:	val_out <= 4'h68dc;
         4'h876b 	:	val_out <= 4'h68dc;
         4'h8770 	:	val_out <= 4'h68c3;
         4'h8771 	:	val_out <= 4'h68c3;
         4'h8772 	:	val_out <= 4'h68c3;
         4'h8773 	:	val_out <= 4'h68c3;
         4'h8778 	:	val_out <= 4'h68aa;
         4'h8779 	:	val_out <= 4'h68aa;
         4'h877a 	:	val_out <= 4'h68aa;
         4'h877b 	:	val_out <= 4'h68aa;
         4'h8780 	:	val_out <= 4'h6892;
         4'h8781 	:	val_out <= 4'h6892;
         4'h8782 	:	val_out <= 4'h6892;
         4'h8783 	:	val_out <= 4'h6892;
         4'h8788 	:	val_out <= 4'h6879;
         4'h8789 	:	val_out <= 4'h6879;
         4'h878a 	:	val_out <= 4'h6879;
         4'h878b 	:	val_out <= 4'h6879;
         4'h8790 	:	val_out <= 4'h6860;
         4'h8791 	:	val_out <= 4'h6860;
         4'h8792 	:	val_out <= 4'h6860;
         4'h8793 	:	val_out <= 4'h6860;
         4'h8798 	:	val_out <= 4'h6848;
         4'h8799 	:	val_out <= 4'h6848;
         4'h879a 	:	val_out <= 4'h6848;
         4'h879b 	:	val_out <= 4'h6848;
         4'h87a0 	:	val_out <= 4'h682f;
         4'h87a1 	:	val_out <= 4'h682f;
         4'h87a2 	:	val_out <= 4'h682f;
         4'h87a3 	:	val_out <= 4'h682f;
         4'h87a8 	:	val_out <= 4'h6816;
         4'h87a9 	:	val_out <= 4'h6816;
         4'h87aa 	:	val_out <= 4'h6816;
         4'h87ab 	:	val_out <= 4'h6816;
         4'h87b0 	:	val_out <= 4'h67fd;
         4'h87b1 	:	val_out <= 4'h67fd;
         4'h87b2 	:	val_out <= 4'h67fd;
         4'h87b3 	:	val_out <= 4'h67fd;
         4'h87b8 	:	val_out <= 4'h67e5;
         4'h87b9 	:	val_out <= 4'h67e5;
         4'h87ba 	:	val_out <= 4'h67e5;
         4'h87bb 	:	val_out <= 4'h67e5;
         4'h87c0 	:	val_out <= 4'h67cc;
         4'h87c1 	:	val_out <= 4'h67cc;
         4'h87c2 	:	val_out <= 4'h67cc;
         4'h87c3 	:	val_out <= 4'h67cc;
         4'h87c8 	:	val_out <= 4'h67b3;
         4'h87c9 	:	val_out <= 4'h67b3;
         4'h87ca 	:	val_out <= 4'h67b3;
         4'h87cb 	:	val_out <= 4'h67b3;
         4'h87d0 	:	val_out <= 4'h679b;
         4'h87d1 	:	val_out <= 4'h679b;
         4'h87d2 	:	val_out <= 4'h679b;
         4'h87d3 	:	val_out <= 4'h679b;
         4'h87d8 	:	val_out <= 4'h6782;
         4'h87d9 	:	val_out <= 4'h6782;
         4'h87da 	:	val_out <= 4'h6782;
         4'h87db 	:	val_out <= 4'h6782;
         4'h87e0 	:	val_out <= 4'h6769;
         4'h87e1 	:	val_out <= 4'h6769;
         4'h87e2 	:	val_out <= 4'h6769;
         4'h87e3 	:	val_out <= 4'h6769;
         4'h87e8 	:	val_out <= 4'h6751;
         4'h87e9 	:	val_out <= 4'h6751;
         4'h87ea 	:	val_out <= 4'h6751;
         4'h87eb 	:	val_out <= 4'h6751;
         4'h87f0 	:	val_out <= 4'h6738;
         4'h87f1 	:	val_out <= 4'h6738;
         4'h87f2 	:	val_out <= 4'h6738;
         4'h87f3 	:	val_out <= 4'h6738;
         4'h87f8 	:	val_out <= 4'h671f;
         4'h87f9 	:	val_out <= 4'h671f;
         4'h87fa 	:	val_out <= 4'h671f;
         4'h87fb 	:	val_out <= 4'h671f;
         4'h8800 	:	val_out <= 4'h6707;
         4'h8801 	:	val_out <= 4'h6707;
         4'h8802 	:	val_out <= 4'h6707;
         4'h8803 	:	val_out <= 4'h6707;
         4'h8808 	:	val_out <= 4'h66ee;
         4'h8809 	:	val_out <= 4'h66ee;
         4'h880a 	:	val_out <= 4'h66ee;
         4'h880b 	:	val_out <= 4'h66ee;
         4'h8810 	:	val_out <= 4'h66d5;
         4'h8811 	:	val_out <= 4'h66d5;
         4'h8812 	:	val_out <= 4'h66d5;
         4'h8813 	:	val_out <= 4'h66d5;
         4'h8818 	:	val_out <= 4'h66bd;
         4'h8819 	:	val_out <= 4'h66bd;
         4'h881a 	:	val_out <= 4'h66bd;
         4'h881b 	:	val_out <= 4'h66bd;
         4'h8820 	:	val_out <= 4'h66a4;
         4'h8821 	:	val_out <= 4'h66a4;
         4'h8822 	:	val_out <= 4'h66a4;
         4'h8823 	:	val_out <= 4'h66a4;
         4'h8828 	:	val_out <= 4'h668c;
         4'h8829 	:	val_out <= 4'h668c;
         4'h882a 	:	val_out <= 4'h668c;
         4'h882b 	:	val_out <= 4'h668c;
         4'h8830 	:	val_out <= 4'h6673;
         4'h8831 	:	val_out <= 4'h6673;
         4'h8832 	:	val_out <= 4'h6673;
         4'h8833 	:	val_out <= 4'h6673;
         4'h8838 	:	val_out <= 4'h665a;
         4'h8839 	:	val_out <= 4'h665a;
         4'h883a 	:	val_out <= 4'h665a;
         4'h883b 	:	val_out <= 4'h665a;
         4'h8840 	:	val_out <= 4'h6642;
         4'h8841 	:	val_out <= 4'h6642;
         4'h8842 	:	val_out <= 4'h6642;
         4'h8843 	:	val_out <= 4'h6642;
         4'h8848 	:	val_out <= 4'h6629;
         4'h8849 	:	val_out <= 4'h6629;
         4'h884a 	:	val_out <= 4'h6629;
         4'h884b 	:	val_out <= 4'h6629;
         4'h8850 	:	val_out <= 4'h6610;
         4'h8851 	:	val_out <= 4'h6610;
         4'h8852 	:	val_out <= 4'h6610;
         4'h8853 	:	val_out <= 4'h6610;
         4'h8858 	:	val_out <= 4'h65f8;
         4'h8859 	:	val_out <= 4'h65f8;
         4'h885a 	:	val_out <= 4'h65f8;
         4'h885b 	:	val_out <= 4'h65f8;
         4'h8860 	:	val_out <= 4'h65df;
         4'h8861 	:	val_out <= 4'h65df;
         4'h8862 	:	val_out <= 4'h65df;
         4'h8863 	:	val_out <= 4'h65df;
         4'h8868 	:	val_out <= 4'h65c7;
         4'h8869 	:	val_out <= 4'h65c7;
         4'h886a 	:	val_out <= 4'h65c7;
         4'h886b 	:	val_out <= 4'h65c7;
         4'h8870 	:	val_out <= 4'h65ae;
         4'h8871 	:	val_out <= 4'h65ae;
         4'h8872 	:	val_out <= 4'h65ae;
         4'h8873 	:	val_out <= 4'h65ae;
         4'h8878 	:	val_out <= 4'h6595;
         4'h8879 	:	val_out <= 4'h6595;
         4'h887a 	:	val_out <= 4'h6595;
         4'h887b 	:	val_out <= 4'h6595;
         4'h8880 	:	val_out <= 4'h657d;
         4'h8881 	:	val_out <= 4'h657d;
         4'h8882 	:	val_out <= 4'h657d;
         4'h8883 	:	val_out <= 4'h657d;
         4'h8888 	:	val_out <= 4'h6564;
         4'h8889 	:	val_out <= 4'h6564;
         4'h888a 	:	val_out <= 4'h6564;
         4'h888b 	:	val_out <= 4'h6564;
         4'h8890 	:	val_out <= 4'h654c;
         4'h8891 	:	val_out <= 4'h654c;
         4'h8892 	:	val_out <= 4'h654c;
         4'h8893 	:	val_out <= 4'h654c;
         4'h8898 	:	val_out <= 4'h6533;
         4'h8899 	:	val_out <= 4'h6533;
         4'h889a 	:	val_out <= 4'h6533;
         4'h889b 	:	val_out <= 4'h6533;
         4'h88a0 	:	val_out <= 4'h651b;
         4'h88a1 	:	val_out <= 4'h651b;
         4'h88a2 	:	val_out <= 4'h651b;
         4'h88a3 	:	val_out <= 4'h651b;
         4'h88a8 	:	val_out <= 4'h6502;
         4'h88a9 	:	val_out <= 4'h6502;
         4'h88aa 	:	val_out <= 4'h6502;
         4'h88ab 	:	val_out <= 4'h6502;
         4'h88b0 	:	val_out <= 4'h64e9;
         4'h88b1 	:	val_out <= 4'h64e9;
         4'h88b2 	:	val_out <= 4'h64e9;
         4'h88b3 	:	val_out <= 4'h64e9;
         4'h88b8 	:	val_out <= 4'h64d1;
         4'h88b9 	:	val_out <= 4'h64d1;
         4'h88ba 	:	val_out <= 4'h64d1;
         4'h88bb 	:	val_out <= 4'h64d1;
         4'h88c0 	:	val_out <= 4'h64b8;
         4'h88c1 	:	val_out <= 4'h64b8;
         4'h88c2 	:	val_out <= 4'h64b8;
         4'h88c3 	:	val_out <= 4'h64b8;
         4'h88c8 	:	val_out <= 4'h64a0;
         4'h88c9 	:	val_out <= 4'h64a0;
         4'h88ca 	:	val_out <= 4'h64a0;
         4'h88cb 	:	val_out <= 4'h64a0;
         4'h88d0 	:	val_out <= 4'h6487;
         4'h88d1 	:	val_out <= 4'h6487;
         4'h88d2 	:	val_out <= 4'h6487;
         4'h88d3 	:	val_out <= 4'h6487;
         4'h88d8 	:	val_out <= 4'h646f;
         4'h88d9 	:	val_out <= 4'h646f;
         4'h88da 	:	val_out <= 4'h646f;
         4'h88db 	:	val_out <= 4'h646f;
         4'h88e0 	:	val_out <= 4'h6456;
         4'h88e1 	:	val_out <= 4'h6456;
         4'h88e2 	:	val_out <= 4'h6456;
         4'h88e3 	:	val_out <= 4'h6456;
         4'h88e8 	:	val_out <= 4'h643e;
         4'h88e9 	:	val_out <= 4'h643e;
         4'h88ea 	:	val_out <= 4'h643e;
         4'h88eb 	:	val_out <= 4'h643e;
         4'h88f0 	:	val_out <= 4'h6425;
         4'h88f1 	:	val_out <= 4'h6425;
         4'h88f2 	:	val_out <= 4'h6425;
         4'h88f3 	:	val_out <= 4'h6425;
         4'h88f8 	:	val_out <= 4'h640d;
         4'h88f9 	:	val_out <= 4'h640d;
         4'h88fa 	:	val_out <= 4'h640d;
         4'h88fb 	:	val_out <= 4'h640d;
         4'h8900 	:	val_out <= 4'h63f4;
         4'h8901 	:	val_out <= 4'h63f4;
         4'h8902 	:	val_out <= 4'h63f4;
         4'h8903 	:	val_out <= 4'h63f4;
         4'h8908 	:	val_out <= 4'h63db;
         4'h8909 	:	val_out <= 4'h63db;
         4'h890a 	:	val_out <= 4'h63db;
         4'h890b 	:	val_out <= 4'h63db;
         4'h8910 	:	val_out <= 4'h63c3;
         4'h8911 	:	val_out <= 4'h63c3;
         4'h8912 	:	val_out <= 4'h63c3;
         4'h8913 	:	val_out <= 4'h63c3;
         4'h8918 	:	val_out <= 4'h63aa;
         4'h8919 	:	val_out <= 4'h63aa;
         4'h891a 	:	val_out <= 4'h63aa;
         4'h891b 	:	val_out <= 4'h63aa;
         4'h8920 	:	val_out <= 4'h6392;
         4'h8921 	:	val_out <= 4'h6392;
         4'h8922 	:	val_out <= 4'h6392;
         4'h8923 	:	val_out <= 4'h6392;
         4'h8928 	:	val_out <= 4'h6379;
         4'h8929 	:	val_out <= 4'h6379;
         4'h892a 	:	val_out <= 4'h6379;
         4'h892b 	:	val_out <= 4'h6379;
         4'h8930 	:	val_out <= 4'h6361;
         4'h8931 	:	val_out <= 4'h6361;
         4'h8932 	:	val_out <= 4'h6361;
         4'h8933 	:	val_out <= 4'h6361;
         4'h8938 	:	val_out <= 4'h6348;
         4'h8939 	:	val_out <= 4'h6348;
         4'h893a 	:	val_out <= 4'h6348;
         4'h893b 	:	val_out <= 4'h6348;
         4'h8940 	:	val_out <= 4'h6330;
         4'h8941 	:	val_out <= 4'h6330;
         4'h8942 	:	val_out <= 4'h6330;
         4'h8943 	:	val_out <= 4'h6330;
         4'h8948 	:	val_out <= 4'h6317;
         4'h8949 	:	val_out <= 4'h6317;
         4'h894a 	:	val_out <= 4'h6317;
         4'h894b 	:	val_out <= 4'h6317;
         4'h8950 	:	val_out <= 4'h62ff;
         4'h8951 	:	val_out <= 4'h62ff;
         4'h8952 	:	val_out <= 4'h62ff;
         4'h8953 	:	val_out <= 4'h62ff;
         4'h8958 	:	val_out <= 4'h62e7;
         4'h8959 	:	val_out <= 4'h62e7;
         4'h895a 	:	val_out <= 4'h62e7;
         4'h895b 	:	val_out <= 4'h62e7;
         4'h8960 	:	val_out <= 4'h62ce;
         4'h8961 	:	val_out <= 4'h62ce;
         4'h8962 	:	val_out <= 4'h62ce;
         4'h8963 	:	val_out <= 4'h62ce;
         4'h8968 	:	val_out <= 4'h62b6;
         4'h8969 	:	val_out <= 4'h62b6;
         4'h896a 	:	val_out <= 4'h62b6;
         4'h896b 	:	val_out <= 4'h62b6;
         4'h8970 	:	val_out <= 4'h629d;
         4'h8971 	:	val_out <= 4'h629d;
         4'h8972 	:	val_out <= 4'h629d;
         4'h8973 	:	val_out <= 4'h629d;
         4'h8978 	:	val_out <= 4'h6285;
         4'h8979 	:	val_out <= 4'h6285;
         4'h897a 	:	val_out <= 4'h6285;
         4'h897b 	:	val_out <= 4'h6285;
         4'h8980 	:	val_out <= 4'h626c;
         4'h8981 	:	val_out <= 4'h626c;
         4'h8982 	:	val_out <= 4'h626c;
         4'h8983 	:	val_out <= 4'h626c;
         4'h8988 	:	val_out <= 4'h6254;
         4'h8989 	:	val_out <= 4'h6254;
         4'h898a 	:	val_out <= 4'h6254;
         4'h898b 	:	val_out <= 4'h6254;
         4'h8990 	:	val_out <= 4'h623b;
         4'h8991 	:	val_out <= 4'h623b;
         4'h8992 	:	val_out <= 4'h623b;
         4'h8993 	:	val_out <= 4'h623b;
         4'h8998 	:	val_out <= 4'h6223;
         4'h8999 	:	val_out <= 4'h6223;
         4'h899a 	:	val_out <= 4'h6223;
         4'h899b 	:	val_out <= 4'h6223;
         4'h89a0 	:	val_out <= 4'h620a;
         4'h89a1 	:	val_out <= 4'h620a;
         4'h89a2 	:	val_out <= 4'h620a;
         4'h89a3 	:	val_out <= 4'h620a;
         4'h89a8 	:	val_out <= 4'h61f2;
         4'h89a9 	:	val_out <= 4'h61f2;
         4'h89aa 	:	val_out <= 4'h61f2;
         4'h89ab 	:	val_out <= 4'h61f2;
         4'h89b0 	:	val_out <= 4'h61da;
         4'h89b1 	:	val_out <= 4'h61da;
         4'h89b2 	:	val_out <= 4'h61da;
         4'h89b3 	:	val_out <= 4'h61da;
         4'h89b8 	:	val_out <= 4'h61c1;
         4'h89b9 	:	val_out <= 4'h61c1;
         4'h89ba 	:	val_out <= 4'h61c1;
         4'h89bb 	:	val_out <= 4'h61c1;
         4'h89c0 	:	val_out <= 4'h61a9;
         4'h89c1 	:	val_out <= 4'h61a9;
         4'h89c2 	:	val_out <= 4'h61a9;
         4'h89c3 	:	val_out <= 4'h61a9;
         4'h89c8 	:	val_out <= 4'h6190;
         4'h89c9 	:	val_out <= 4'h6190;
         4'h89ca 	:	val_out <= 4'h6190;
         4'h89cb 	:	val_out <= 4'h6190;
         4'h89d0 	:	val_out <= 4'h6178;
         4'h89d1 	:	val_out <= 4'h6178;
         4'h89d2 	:	val_out <= 4'h6178;
         4'h89d3 	:	val_out <= 4'h6178;
         4'h89d8 	:	val_out <= 4'h615f;
         4'h89d9 	:	val_out <= 4'h615f;
         4'h89da 	:	val_out <= 4'h615f;
         4'h89db 	:	val_out <= 4'h615f;
         4'h89e0 	:	val_out <= 4'h6147;
         4'h89e1 	:	val_out <= 4'h6147;
         4'h89e2 	:	val_out <= 4'h6147;
         4'h89e3 	:	val_out <= 4'h6147;
         4'h89e8 	:	val_out <= 4'h612f;
         4'h89e9 	:	val_out <= 4'h612f;
         4'h89ea 	:	val_out <= 4'h612f;
         4'h89eb 	:	val_out <= 4'h612f;
         4'h89f0 	:	val_out <= 4'h6116;
         4'h89f1 	:	val_out <= 4'h6116;
         4'h89f2 	:	val_out <= 4'h6116;
         4'h89f3 	:	val_out <= 4'h6116;
         4'h89f8 	:	val_out <= 4'h60fe;
         4'h89f9 	:	val_out <= 4'h60fe;
         4'h89fa 	:	val_out <= 4'h60fe;
         4'h89fb 	:	val_out <= 4'h60fe;
         4'h8a00 	:	val_out <= 4'h60e6;
         4'h8a01 	:	val_out <= 4'h60e6;
         4'h8a02 	:	val_out <= 4'h60e6;
         4'h8a03 	:	val_out <= 4'h60e6;
         4'h8a08 	:	val_out <= 4'h60cd;
         4'h8a09 	:	val_out <= 4'h60cd;
         4'h8a0a 	:	val_out <= 4'h60cd;
         4'h8a0b 	:	val_out <= 4'h60cd;
         4'h8a10 	:	val_out <= 4'h60b5;
         4'h8a11 	:	val_out <= 4'h60b5;
         4'h8a12 	:	val_out <= 4'h60b5;
         4'h8a13 	:	val_out <= 4'h60b5;
         4'h8a18 	:	val_out <= 4'h609c;
         4'h8a19 	:	val_out <= 4'h609c;
         4'h8a1a 	:	val_out <= 4'h609c;
         4'h8a1b 	:	val_out <= 4'h609c;
         4'h8a20 	:	val_out <= 4'h6084;
         4'h8a21 	:	val_out <= 4'h6084;
         4'h8a22 	:	val_out <= 4'h6084;
         4'h8a23 	:	val_out <= 4'h6084;
         4'h8a28 	:	val_out <= 4'h606c;
         4'h8a29 	:	val_out <= 4'h606c;
         4'h8a2a 	:	val_out <= 4'h606c;
         4'h8a2b 	:	val_out <= 4'h606c;
         4'h8a30 	:	val_out <= 4'h6053;
         4'h8a31 	:	val_out <= 4'h6053;
         4'h8a32 	:	val_out <= 4'h6053;
         4'h8a33 	:	val_out <= 4'h6053;
         4'h8a38 	:	val_out <= 4'h603b;
         4'h8a39 	:	val_out <= 4'h603b;
         4'h8a3a 	:	val_out <= 4'h603b;
         4'h8a3b 	:	val_out <= 4'h603b;
         4'h8a40 	:	val_out <= 4'h6023;
         4'h8a41 	:	val_out <= 4'h6023;
         4'h8a42 	:	val_out <= 4'h6023;
         4'h8a43 	:	val_out <= 4'h6023;
         4'h8a48 	:	val_out <= 4'h600a;
         4'h8a49 	:	val_out <= 4'h600a;
         4'h8a4a 	:	val_out <= 4'h600a;
         4'h8a4b 	:	val_out <= 4'h600a;
         4'h8a50 	:	val_out <= 4'h5ff2;
         4'h8a51 	:	val_out <= 4'h5ff2;
         4'h8a52 	:	val_out <= 4'h5ff2;
         4'h8a53 	:	val_out <= 4'h5ff2;
         4'h8a58 	:	val_out <= 4'h5fda;
         4'h8a59 	:	val_out <= 4'h5fda;
         4'h8a5a 	:	val_out <= 4'h5fda;
         4'h8a5b 	:	val_out <= 4'h5fda;
         4'h8a60 	:	val_out <= 4'h5fc1;
         4'h8a61 	:	val_out <= 4'h5fc1;
         4'h8a62 	:	val_out <= 4'h5fc1;
         4'h8a63 	:	val_out <= 4'h5fc1;
         4'h8a68 	:	val_out <= 4'h5fa9;
         4'h8a69 	:	val_out <= 4'h5fa9;
         4'h8a6a 	:	val_out <= 4'h5fa9;
         4'h8a6b 	:	val_out <= 4'h5fa9;
         4'h8a70 	:	val_out <= 4'h5f91;
         4'h8a71 	:	val_out <= 4'h5f91;
         4'h8a72 	:	val_out <= 4'h5f91;
         4'h8a73 	:	val_out <= 4'h5f91;
         4'h8a78 	:	val_out <= 4'h5f78;
         4'h8a79 	:	val_out <= 4'h5f78;
         4'h8a7a 	:	val_out <= 4'h5f78;
         4'h8a7b 	:	val_out <= 4'h5f78;
         4'h8a80 	:	val_out <= 4'h5f60;
         4'h8a81 	:	val_out <= 4'h5f60;
         4'h8a82 	:	val_out <= 4'h5f60;
         4'h8a83 	:	val_out <= 4'h5f60;
         4'h8a88 	:	val_out <= 4'h5f48;
         4'h8a89 	:	val_out <= 4'h5f48;
         4'h8a8a 	:	val_out <= 4'h5f48;
         4'h8a8b 	:	val_out <= 4'h5f48;
         4'h8a90 	:	val_out <= 4'h5f2f;
         4'h8a91 	:	val_out <= 4'h5f2f;
         4'h8a92 	:	val_out <= 4'h5f2f;
         4'h8a93 	:	val_out <= 4'h5f2f;
         4'h8a98 	:	val_out <= 4'h5f17;
         4'h8a99 	:	val_out <= 4'h5f17;
         4'h8a9a 	:	val_out <= 4'h5f17;
         4'h8a9b 	:	val_out <= 4'h5f17;
         4'h8aa0 	:	val_out <= 4'h5eff;
         4'h8aa1 	:	val_out <= 4'h5eff;
         4'h8aa2 	:	val_out <= 4'h5eff;
         4'h8aa3 	:	val_out <= 4'h5eff;
         4'h8aa8 	:	val_out <= 4'h5ee7;
         4'h8aa9 	:	val_out <= 4'h5ee7;
         4'h8aaa 	:	val_out <= 4'h5ee7;
         4'h8aab 	:	val_out <= 4'h5ee7;
         4'h8ab0 	:	val_out <= 4'h5ece;
         4'h8ab1 	:	val_out <= 4'h5ece;
         4'h8ab2 	:	val_out <= 4'h5ece;
         4'h8ab3 	:	val_out <= 4'h5ece;
         4'h8ab8 	:	val_out <= 4'h5eb6;
         4'h8ab9 	:	val_out <= 4'h5eb6;
         4'h8aba 	:	val_out <= 4'h5eb6;
         4'h8abb 	:	val_out <= 4'h5eb6;
         4'h8ac0 	:	val_out <= 4'h5e9e;
         4'h8ac1 	:	val_out <= 4'h5e9e;
         4'h8ac2 	:	val_out <= 4'h5e9e;
         4'h8ac3 	:	val_out <= 4'h5e9e;
         4'h8ac8 	:	val_out <= 4'h5e86;
         4'h8ac9 	:	val_out <= 4'h5e86;
         4'h8aca 	:	val_out <= 4'h5e86;
         4'h8acb 	:	val_out <= 4'h5e86;
         4'h8ad0 	:	val_out <= 4'h5e6d;
         4'h8ad1 	:	val_out <= 4'h5e6d;
         4'h8ad2 	:	val_out <= 4'h5e6d;
         4'h8ad3 	:	val_out <= 4'h5e6d;
         4'h8ad8 	:	val_out <= 4'h5e55;
         4'h8ad9 	:	val_out <= 4'h5e55;
         4'h8ada 	:	val_out <= 4'h5e55;
         4'h8adb 	:	val_out <= 4'h5e55;
         4'h8ae0 	:	val_out <= 4'h5e3d;
         4'h8ae1 	:	val_out <= 4'h5e3d;
         4'h8ae2 	:	val_out <= 4'h5e3d;
         4'h8ae3 	:	val_out <= 4'h5e3d;
         4'h8ae8 	:	val_out <= 4'h5e25;
         4'h8ae9 	:	val_out <= 4'h5e25;
         4'h8aea 	:	val_out <= 4'h5e25;
         4'h8aeb 	:	val_out <= 4'h5e25;
         4'h8af0 	:	val_out <= 4'h5e0c;
         4'h8af1 	:	val_out <= 4'h5e0c;
         4'h8af2 	:	val_out <= 4'h5e0c;
         4'h8af3 	:	val_out <= 4'h5e0c;
         4'h8af8 	:	val_out <= 4'h5df4;
         4'h8af9 	:	val_out <= 4'h5df4;
         4'h8afa 	:	val_out <= 4'h5df4;
         4'h8afb 	:	val_out <= 4'h5df4;
         4'h8b00 	:	val_out <= 4'h5ddc;
         4'h8b01 	:	val_out <= 4'h5ddc;
         4'h8b02 	:	val_out <= 4'h5ddc;
         4'h8b03 	:	val_out <= 4'h5ddc;
         4'h8b08 	:	val_out <= 4'h5dc4;
         4'h8b09 	:	val_out <= 4'h5dc4;
         4'h8b0a 	:	val_out <= 4'h5dc4;
         4'h8b0b 	:	val_out <= 4'h5dc4;
         4'h8b10 	:	val_out <= 4'h5dab;
         4'h8b11 	:	val_out <= 4'h5dab;
         4'h8b12 	:	val_out <= 4'h5dab;
         4'h8b13 	:	val_out <= 4'h5dab;
         4'h8b18 	:	val_out <= 4'h5d93;
         4'h8b19 	:	val_out <= 4'h5d93;
         4'h8b1a 	:	val_out <= 4'h5d93;
         4'h8b1b 	:	val_out <= 4'h5d93;
         4'h8b20 	:	val_out <= 4'h5d7b;
         4'h8b21 	:	val_out <= 4'h5d7b;
         4'h8b22 	:	val_out <= 4'h5d7b;
         4'h8b23 	:	val_out <= 4'h5d7b;
         4'h8b28 	:	val_out <= 4'h5d63;
         4'h8b29 	:	val_out <= 4'h5d63;
         4'h8b2a 	:	val_out <= 4'h5d63;
         4'h8b2b 	:	val_out <= 4'h5d63;
         4'h8b30 	:	val_out <= 4'h5d4b;
         4'h8b31 	:	val_out <= 4'h5d4b;
         4'h8b32 	:	val_out <= 4'h5d4b;
         4'h8b33 	:	val_out <= 4'h5d4b;
         4'h8b38 	:	val_out <= 4'h5d32;
         4'h8b39 	:	val_out <= 4'h5d32;
         4'h8b3a 	:	val_out <= 4'h5d32;
         4'h8b3b 	:	val_out <= 4'h5d32;
         4'h8b40 	:	val_out <= 4'h5d1a;
         4'h8b41 	:	val_out <= 4'h5d1a;
         4'h8b42 	:	val_out <= 4'h5d1a;
         4'h8b43 	:	val_out <= 4'h5d1a;
         4'h8b48 	:	val_out <= 4'h5d02;
         4'h8b49 	:	val_out <= 4'h5d02;
         4'h8b4a 	:	val_out <= 4'h5d02;
         4'h8b4b 	:	val_out <= 4'h5d02;
         4'h8b50 	:	val_out <= 4'h5cea;
         4'h8b51 	:	val_out <= 4'h5cea;
         4'h8b52 	:	val_out <= 4'h5cea;
         4'h8b53 	:	val_out <= 4'h5cea;
         4'h8b58 	:	val_out <= 4'h5cd2;
         4'h8b59 	:	val_out <= 4'h5cd2;
         4'h8b5a 	:	val_out <= 4'h5cd2;
         4'h8b5b 	:	val_out <= 4'h5cd2;
         4'h8b60 	:	val_out <= 4'h5cba;
         4'h8b61 	:	val_out <= 4'h5cba;
         4'h8b62 	:	val_out <= 4'h5cba;
         4'h8b63 	:	val_out <= 4'h5cba;
         4'h8b68 	:	val_out <= 4'h5ca1;
         4'h8b69 	:	val_out <= 4'h5ca1;
         4'h8b6a 	:	val_out <= 4'h5ca1;
         4'h8b6b 	:	val_out <= 4'h5ca1;
         4'h8b70 	:	val_out <= 4'h5c89;
         4'h8b71 	:	val_out <= 4'h5c89;
         4'h8b72 	:	val_out <= 4'h5c89;
         4'h8b73 	:	val_out <= 4'h5c89;
         4'h8b78 	:	val_out <= 4'h5c71;
         4'h8b79 	:	val_out <= 4'h5c71;
         4'h8b7a 	:	val_out <= 4'h5c71;
         4'h8b7b 	:	val_out <= 4'h5c71;
         4'h8b80 	:	val_out <= 4'h5c59;
         4'h8b81 	:	val_out <= 4'h5c59;
         4'h8b82 	:	val_out <= 4'h5c59;
         4'h8b83 	:	val_out <= 4'h5c59;
         4'h8b88 	:	val_out <= 4'h5c41;
         4'h8b89 	:	val_out <= 4'h5c41;
         4'h8b8a 	:	val_out <= 4'h5c41;
         4'h8b8b 	:	val_out <= 4'h5c41;
         4'h8b90 	:	val_out <= 4'h5c29;
         4'h8b91 	:	val_out <= 4'h5c29;
         4'h8b92 	:	val_out <= 4'h5c29;
         4'h8b93 	:	val_out <= 4'h5c29;
         4'h8b98 	:	val_out <= 4'h5c11;
         4'h8b99 	:	val_out <= 4'h5c11;
         4'h8b9a 	:	val_out <= 4'h5c11;
         4'h8b9b 	:	val_out <= 4'h5c11;
         4'h8ba0 	:	val_out <= 4'h5bf8;
         4'h8ba1 	:	val_out <= 4'h5bf8;
         4'h8ba2 	:	val_out <= 4'h5bf8;
         4'h8ba3 	:	val_out <= 4'h5bf8;
         4'h8ba8 	:	val_out <= 4'h5be0;
         4'h8ba9 	:	val_out <= 4'h5be0;
         4'h8baa 	:	val_out <= 4'h5be0;
         4'h8bab 	:	val_out <= 4'h5be0;
         4'h8bb0 	:	val_out <= 4'h5bc8;
         4'h8bb1 	:	val_out <= 4'h5bc8;
         4'h8bb2 	:	val_out <= 4'h5bc8;
         4'h8bb3 	:	val_out <= 4'h5bc8;
         4'h8bb8 	:	val_out <= 4'h5bb0;
         4'h8bb9 	:	val_out <= 4'h5bb0;
         4'h8bba 	:	val_out <= 4'h5bb0;
         4'h8bbb 	:	val_out <= 4'h5bb0;
         4'h8bc0 	:	val_out <= 4'h5b98;
         4'h8bc1 	:	val_out <= 4'h5b98;
         4'h8bc2 	:	val_out <= 4'h5b98;
         4'h8bc3 	:	val_out <= 4'h5b98;
         4'h8bc8 	:	val_out <= 4'h5b80;
         4'h8bc9 	:	val_out <= 4'h5b80;
         4'h8bca 	:	val_out <= 4'h5b80;
         4'h8bcb 	:	val_out <= 4'h5b80;
         4'h8bd0 	:	val_out <= 4'h5b68;
         4'h8bd1 	:	val_out <= 4'h5b68;
         4'h8bd2 	:	val_out <= 4'h5b68;
         4'h8bd3 	:	val_out <= 4'h5b68;
         4'h8bd8 	:	val_out <= 4'h5b50;
         4'h8bd9 	:	val_out <= 4'h5b50;
         4'h8bda 	:	val_out <= 4'h5b50;
         4'h8bdb 	:	val_out <= 4'h5b50;
         4'h8be0 	:	val_out <= 4'h5b38;
         4'h8be1 	:	val_out <= 4'h5b38;
         4'h8be2 	:	val_out <= 4'h5b38;
         4'h8be3 	:	val_out <= 4'h5b38;
         4'h8be8 	:	val_out <= 4'h5b20;
         4'h8be9 	:	val_out <= 4'h5b20;
         4'h8bea 	:	val_out <= 4'h5b20;
         4'h8beb 	:	val_out <= 4'h5b20;
         4'h8bf0 	:	val_out <= 4'h5b08;
         4'h8bf1 	:	val_out <= 4'h5b08;
         4'h8bf2 	:	val_out <= 4'h5b08;
         4'h8bf3 	:	val_out <= 4'h5b08;
         4'h8bf8 	:	val_out <= 4'h5af0;
         4'h8bf9 	:	val_out <= 4'h5af0;
         4'h8bfa 	:	val_out <= 4'h5af0;
         4'h8bfb 	:	val_out <= 4'h5af0;
         4'h8c00 	:	val_out <= 4'h5ad7;
         4'h8c01 	:	val_out <= 4'h5ad7;
         4'h8c02 	:	val_out <= 4'h5ad7;
         4'h8c03 	:	val_out <= 4'h5ad7;
         4'h8c08 	:	val_out <= 4'h5abf;
         4'h8c09 	:	val_out <= 4'h5abf;
         4'h8c0a 	:	val_out <= 4'h5abf;
         4'h8c0b 	:	val_out <= 4'h5abf;
         4'h8c10 	:	val_out <= 4'h5aa7;
         4'h8c11 	:	val_out <= 4'h5aa7;
         4'h8c12 	:	val_out <= 4'h5aa7;
         4'h8c13 	:	val_out <= 4'h5aa7;
         4'h8c18 	:	val_out <= 4'h5a8f;
         4'h8c19 	:	val_out <= 4'h5a8f;
         4'h8c1a 	:	val_out <= 4'h5a8f;
         4'h8c1b 	:	val_out <= 4'h5a8f;
         4'h8c20 	:	val_out <= 4'h5a77;
         4'h8c21 	:	val_out <= 4'h5a77;
         4'h8c22 	:	val_out <= 4'h5a77;
         4'h8c23 	:	val_out <= 4'h5a77;
         4'h8c28 	:	val_out <= 4'h5a5f;
         4'h8c29 	:	val_out <= 4'h5a5f;
         4'h8c2a 	:	val_out <= 4'h5a5f;
         4'h8c2b 	:	val_out <= 4'h5a5f;
         4'h8c30 	:	val_out <= 4'h5a47;
         4'h8c31 	:	val_out <= 4'h5a47;
         4'h8c32 	:	val_out <= 4'h5a47;
         4'h8c33 	:	val_out <= 4'h5a47;
         4'h8c38 	:	val_out <= 4'h5a2f;
         4'h8c39 	:	val_out <= 4'h5a2f;
         4'h8c3a 	:	val_out <= 4'h5a2f;
         4'h8c3b 	:	val_out <= 4'h5a2f;
         4'h8c40 	:	val_out <= 4'h5a17;
         4'h8c41 	:	val_out <= 4'h5a17;
         4'h8c42 	:	val_out <= 4'h5a17;
         4'h8c43 	:	val_out <= 4'h5a17;
         4'h8c48 	:	val_out <= 4'h59ff;
         4'h8c49 	:	val_out <= 4'h59ff;
         4'h8c4a 	:	val_out <= 4'h59ff;
         4'h8c4b 	:	val_out <= 4'h59ff;
         4'h8c50 	:	val_out <= 4'h59e7;
         4'h8c51 	:	val_out <= 4'h59e7;
         4'h8c52 	:	val_out <= 4'h59e7;
         4'h8c53 	:	val_out <= 4'h59e7;
         4'h8c58 	:	val_out <= 4'h59cf;
         4'h8c59 	:	val_out <= 4'h59cf;
         4'h8c5a 	:	val_out <= 4'h59cf;
         4'h8c5b 	:	val_out <= 4'h59cf;
         4'h8c60 	:	val_out <= 4'h59b7;
         4'h8c61 	:	val_out <= 4'h59b7;
         4'h8c62 	:	val_out <= 4'h59b7;
         4'h8c63 	:	val_out <= 4'h59b7;
         4'h8c68 	:	val_out <= 4'h599f;
         4'h8c69 	:	val_out <= 4'h599f;
         4'h8c6a 	:	val_out <= 4'h599f;
         4'h8c6b 	:	val_out <= 4'h599f;
         4'h8c70 	:	val_out <= 4'h5987;
         4'h8c71 	:	val_out <= 4'h5987;
         4'h8c72 	:	val_out <= 4'h5987;
         4'h8c73 	:	val_out <= 4'h5987;
         4'h8c78 	:	val_out <= 4'h596f;
         4'h8c79 	:	val_out <= 4'h596f;
         4'h8c7a 	:	val_out <= 4'h596f;
         4'h8c7b 	:	val_out <= 4'h596f;
         4'h8c80 	:	val_out <= 4'h5957;
         4'h8c81 	:	val_out <= 4'h5957;
         4'h8c82 	:	val_out <= 4'h5957;
         4'h8c83 	:	val_out <= 4'h5957;
         4'h8c88 	:	val_out <= 4'h593f;
         4'h8c89 	:	val_out <= 4'h593f;
         4'h8c8a 	:	val_out <= 4'h593f;
         4'h8c8b 	:	val_out <= 4'h593f;
         4'h8c90 	:	val_out <= 4'h5927;
         4'h8c91 	:	val_out <= 4'h5927;
         4'h8c92 	:	val_out <= 4'h5927;
         4'h8c93 	:	val_out <= 4'h5927;
         4'h8c98 	:	val_out <= 4'h5910;
         4'h8c99 	:	val_out <= 4'h5910;
         4'h8c9a 	:	val_out <= 4'h5910;
         4'h8c9b 	:	val_out <= 4'h5910;
         4'h8ca0 	:	val_out <= 4'h58f8;
         4'h8ca1 	:	val_out <= 4'h58f8;
         4'h8ca2 	:	val_out <= 4'h58f8;
         4'h8ca3 	:	val_out <= 4'h58f8;
         4'h8ca8 	:	val_out <= 4'h58e0;
         4'h8ca9 	:	val_out <= 4'h58e0;
         4'h8caa 	:	val_out <= 4'h58e0;
         4'h8cab 	:	val_out <= 4'h58e0;
         4'h8cb0 	:	val_out <= 4'h58c8;
         4'h8cb1 	:	val_out <= 4'h58c8;
         4'h8cb2 	:	val_out <= 4'h58c8;
         4'h8cb3 	:	val_out <= 4'h58c8;
         4'h8cb8 	:	val_out <= 4'h58b0;
         4'h8cb9 	:	val_out <= 4'h58b0;
         4'h8cba 	:	val_out <= 4'h58b0;
         4'h8cbb 	:	val_out <= 4'h58b0;
         4'h8cc0 	:	val_out <= 4'h5898;
         4'h8cc1 	:	val_out <= 4'h5898;
         4'h8cc2 	:	val_out <= 4'h5898;
         4'h8cc3 	:	val_out <= 4'h5898;
         4'h8cc8 	:	val_out <= 4'h5880;
         4'h8cc9 	:	val_out <= 4'h5880;
         4'h8cca 	:	val_out <= 4'h5880;
         4'h8ccb 	:	val_out <= 4'h5880;
         4'h8cd0 	:	val_out <= 4'h5868;
         4'h8cd1 	:	val_out <= 4'h5868;
         4'h8cd2 	:	val_out <= 4'h5868;
         4'h8cd3 	:	val_out <= 4'h5868;
         4'h8cd8 	:	val_out <= 4'h5850;
         4'h8cd9 	:	val_out <= 4'h5850;
         4'h8cda 	:	val_out <= 4'h5850;
         4'h8cdb 	:	val_out <= 4'h5850;
         4'h8ce0 	:	val_out <= 4'h5838;
         4'h8ce1 	:	val_out <= 4'h5838;
         4'h8ce2 	:	val_out <= 4'h5838;
         4'h8ce3 	:	val_out <= 4'h5838;
         4'h8ce8 	:	val_out <= 4'h5820;
         4'h8ce9 	:	val_out <= 4'h5820;
         4'h8cea 	:	val_out <= 4'h5820;
         4'h8ceb 	:	val_out <= 4'h5820;
         4'h8cf0 	:	val_out <= 4'h5809;
         4'h8cf1 	:	val_out <= 4'h5809;
         4'h8cf2 	:	val_out <= 4'h5809;
         4'h8cf3 	:	val_out <= 4'h5809;
         4'h8cf8 	:	val_out <= 4'h57f1;
         4'h8cf9 	:	val_out <= 4'h57f1;
         4'h8cfa 	:	val_out <= 4'h57f1;
         4'h8cfb 	:	val_out <= 4'h57f1;
         4'h8d00 	:	val_out <= 4'h57d9;
         4'h8d01 	:	val_out <= 4'h57d9;
         4'h8d02 	:	val_out <= 4'h57d9;
         4'h8d03 	:	val_out <= 4'h57d9;
         4'h8d08 	:	val_out <= 4'h57c1;
         4'h8d09 	:	val_out <= 4'h57c1;
         4'h8d0a 	:	val_out <= 4'h57c1;
         4'h8d0b 	:	val_out <= 4'h57c1;
         4'h8d10 	:	val_out <= 4'h57a9;
         4'h8d11 	:	val_out <= 4'h57a9;
         4'h8d12 	:	val_out <= 4'h57a9;
         4'h8d13 	:	val_out <= 4'h57a9;
         4'h8d18 	:	val_out <= 4'h5791;
         4'h8d19 	:	val_out <= 4'h5791;
         4'h8d1a 	:	val_out <= 4'h5791;
         4'h8d1b 	:	val_out <= 4'h5791;
         4'h8d20 	:	val_out <= 4'h5779;
         4'h8d21 	:	val_out <= 4'h5779;
         4'h8d22 	:	val_out <= 4'h5779;
         4'h8d23 	:	val_out <= 4'h5779;
         4'h8d28 	:	val_out <= 4'h5762;
         4'h8d29 	:	val_out <= 4'h5762;
         4'h8d2a 	:	val_out <= 4'h5762;
         4'h8d2b 	:	val_out <= 4'h5762;
         4'h8d30 	:	val_out <= 4'h574a;
         4'h8d31 	:	val_out <= 4'h574a;
         4'h8d32 	:	val_out <= 4'h574a;
         4'h8d33 	:	val_out <= 4'h574a;
         4'h8d38 	:	val_out <= 4'h5732;
         4'h8d39 	:	val_out <= 4'h5732;
         4'h8d3a 	:	val_out <= 4'h5732;
         4'h8d3b 	:	val_out <= 4'h5732;
         4'h8d40 	:	val_out <= 4'h571a;
         4'h8d41 	:	val_out <= 4'h571a;
         4'h8d42 	:	val_out <= 4'h571a;
         4'h8d43 	:	val_out <= 4'h571a;
         4'h8d48 	:	val_out <= 4'h5702;
         4'h8d49 	:	val_out <= 4'h5702;
         4'h8d4a 	:	val_out <= 4'h5702;
         4'h8d4b 	:	val_out <= 4'h5702;
         4'h8d50 	:	val_out <= 4'h56ea;
         4'h8d51 	:	val_out <= 4'h56ea;
         4'h8d52 	:	val_out <= 4'h56ea;
         4'h8d53 	:	val_out <= 4'h56ea;
         4'h8d58 	:	val_out <= 4'h56d3;
         4'h8d59 	:	val_out <= 4'h56d3;
         4'h8d5a 	:	val_out <= 4'h56d3;
         4'h8d5b 	:	val_out <= 4'h56d3;
         4'h8d60 	:	val_out <= 4'h56bb;
         4'h8d61 	:	val_out <= 4'h56bb;
         4'h8d62 	:	val_out <= 4'h56bb;
         4'h8d63 	:	val_out <= 4'h56bb;
         4'h8d68 	:	val_out <= 4'h56a3;
         4'h8d69 	:	val_out <= 4'h56a3;
         4'h8d6a 	:	val_out <= 4'h56a3;
         4'h8d6b 	:	val_out <= 4'h56a3;
         4'h8d70 	:	val_out <= 4'h568b;
         4'h8d71 	:	val_out <= 4'h568b;
         4'h8d72 	:	val_out <= 4'h568b;
         4'h8d73 	:	val_out <= 4'h568b;
         4'h8d78 	:	val_out <= 4'h5674;
         4'h8d79 	:	val_out <= 4'h5674;
         4'h8d7a 	:	val_out <= 4'h5674;
         4'h8d7b 	:	val_out <= 4'h5674;
         4'h8d80 	:	val_out <= 4'h565c;
         4'h8d81 	:	val_out <= 4'h565c;
         4'h8d82 	:	val_out <= 4'h565c;
         4'h8d83 	:	val_out <= 4'h565c;
         4'h8d88 	:	val_out <= 4'h5644;
         4'h8d89 	:	val_out <= 4'h5644;
         4'h8d8a 	:	val_out <= 4'h5644;
         4'h8d8b 	:	val_out <= 4'h5644;
         4'h8d90 	:	val_out <= 4'h562c;
         4'h8d91 	:	val_out <= 4'h562c;
         4'h8d92 	:	val_out <= 4'h562c;
         4'h8d93 	:	val_out <= 4'h562c;
         4'h8d98 	:	val_out <= 4'h5614;
         4'h8d99 	:	val_out <= 4'h5614;
         4'h8d9a 	:	val_out <= 4'h5614;
         4'h8d9b 	:	val_out <= 4'h5614;
         4'h8da0 	:	val_out <= 4'h55fd;
         4'h8da1 	:	val_out <= 4'h55fd;
         4'h8da2 	:	val_out <= 4'h55fd;
         4'h8da3 	:	val_out <= 4'h55fd;
         4'h8da8 	:	val_out <= 4'h55e5;
         4'h8da9 	:	val_out <= 4'h55e5;
         4'h8daa 	:	val_out <= 4'h55e5;
         4'h8dab 	:	val_out <= 4'h55e5;
         4'h8db0 	:	val_out <= 4'h55cd;
         4'h8db1 	:	val_out <= 4'h55cd;
         4'h8db2 	:	val_out <= 4'h55cd;
         4'h8db3 	:	val_out <= 4'h55cd;
         4'h8db8 	:	val_out <= 4'h55b6;
         4'h8db9 	:	val_out <= 4'h55b6;
         4'h8dba 	:	val_out <= 4'h55b6;
         4'h8dbb 	:	val_out <= 4'h55b6;
         4'h8dc0 	:	val_out <= 4'h559e;
         4'h8dc1 	:	val_out <= 4'h559e;
         4'h8dc2 	:	val_out <= 4'h559e;
         4'h8dc3 	:	val_out <= 4'h559e;
         4'h8dc8 	:	val_out <= 4'h5586;
         4'h8dc9 	:	val_out <= 4'h5586;
         4'h8dca 	:	val_out <= 4'h5586;
         4'h8dcb 	:	val_out <= 4'h5586;
         4'h8dd0 	:	val_out <= 4'h556e;
         4'h8dd1 	:	val_out <= 4'h556e;
         4'h8dd2 	:	val_out <= 4'h556e;
         4'h8dd3 	:	val_out <= 4'h556e;
         4'h8dd8 	:	val_out <= 4'h5557;
         4'h8dd9 	:	val_out <= 4'h5557;
         4'h8dda 	:	val_out <= 4'h5557;
         4'h8ddb 	:	val_out <= 4'h5557;
         4'h8de0 	:	val_out <= 4'h553f;
         4'h8de1 	:	val_out <= 4'h553f;
         4'h8de2 	:	val_out <= 4'h553f;
         4'h8de3 	:	val_out <= 4'h553f;
         4'h8de8 	:	val_out <= 4'h5527;
         4'h8de9 	:	val_out <= 4'h5527;
         4'h8dea 	:	val_out <= 4'h5527;
         4'h8deb 	:	val_out <= 4'h5527;
         4'h8df0 	:	val_out <= 4'h5510;
         4'h8df1 	:	val_out <= 4'h5510;
         4'h8df2 	:	val_out <= 4'h5510;
         4'h8df3 	:	val_out <= 4'h5510;
         4'h8df8 	:	val_out <= 4'h54f8;
         4'h8df9 	:	val_out <= 4'h54f8;
         4'h8dfa 	:	val_out <= 4'h54f8;
         4'h8dfb 	:	val_out <= 4'h54f8;
         4'h8e00 	:	val_out <= 4'h54e0;
         4'h8e01 	:	val_out <= 4'h54e0;
         4'h8e02 	:	val_out <= 4'h54e0;
         4'h8e03 	:	val_out <= 4'h54e0;
         4'h8e08 	:	val_out <= 4'h54c9;
         4'h8e09 	:	val_out <= 4'h54c9;
         4'h8e0a 	:	val_out <= 4'h54c9;
         4'h8e0b 	:	val_out <= 4'h54c9;
         4'h8e10 	:	val_out <= 4'h54b1;
         4'h8e11 	:	val_out <= 4'h54b1;
         4'h8e12 	:	val_out <= 4'h54b1;
         4'h8e13 	:	val_out <= 4'h54b1;
         4'h8e18 	:	val_out <= 4'h5499;
         4'h8e19 	:	val_out <= 4'h5499;
         4'h8e1a 	:	val_out <= 4'h5499;
         4'h8e1b 	:	val_out <= 4'h5499;
         4'h8e20 	:	val_out <= 4'h5482;
         4'h8e21 	:	val_out <= 4'h5482;
         4'h8e22 	:	val_out <= 4'h5482;
         4'h8e23 	:	val_out <= 4'h5482;
         4'h8e28 	:	val_out <= 4'h546a;
         4'h8e29 	:	val_out <= 4'h546a;
         4'h8e2a 	:	val_out <= 4'h546a;
         4'h8e2b 	:	val_out <= 4'h546a;
         4'h8e30 	:	val_out <= 4'h5452;
         4'h8e31 	:	val_out <= 4'h5452;
         4'h8e32 	:	val_out <= 4'h5452;
         4'h8e33 	:	val_out <= 4'h5452;
         4'h8e38 	:	val_out <= 4'h543b;
         4'h8e39 	:	val_out <= 4'h543b;
         4'h8e3a 	:	val_out <= 4'h543b;
         4'h8e3b 	:	val_out <= 4'h543b;
         4'h8e40 	:	val_out <= 4'h5423;
         4'h8e41 	:	val_out <= 4'h5423;
         4'h8e42 	:	val_out <= 4'h5423;
         4'h8e43 	:	val_out <= 4'h5423;
         4'h8e48 	:	val_out <= 4'h540c;
         4'h8e49 	:	val_out <= 4'h540c;
         4'h8e4a 	:	val_out <= 4'h540c;
         4'h8e4b 	:	val_out <= 4'h540c;
         4'h8e50 	:	val_out <= 4'h53f4;
         4'h8e51 	:	val_out <= 4'h53f4;
         4'h8e52 	:	val_out <= 4'h53f4;
         4'h8e53 	:	val_out <= 4'h53f4;
         4'h8e58 	:	val_out <= 4'h53dc;
         4'h8e59 	:	val_out <= 4'h53dc;
         4'h8e5a 	:	val_out <= 4'h53dc;
         4'h8e5b 	:	val_out <= 4'h53dc;
         4'h8e60 	:	val_out <= 4'h53c5;
         4'h8e61 	:	val_out <= 4'h53c5;
         4'h8e62 	:	val_out <= 4'h53c5;
         4'h8e63 	:	val_out <= 4'h53c5;
         4'h8e68 	:	val_out <= 4'h53ad;
         4'h8e69 	:	val_out <= 4'h53ad;
         4'h8e6a 	:	val_out <= 4'h53ad;
         4'h8e6b 	:	val_out <= 4'h53ad;
         4'h8e70 	:	val_out <= 4'h5396;
         4'h8e71 	:	val_out <= 4'h5396;
         4'h8e72 	:	val_out <= 4'h5396;
         4'h8e73 	:	val_out <= 4'h5396;
         4'h8e78 	:	val_out <= 4'h537e;
         4'h8e79 	:	val_out <= 4'h537e;
         4'h8e7a 	:	val_out <= 4'h537e;
         4'h8e7b 	:	val_out <= 4'h537e;
         4'h8e80 	:	val_out <= 4'h5367;
         4'h8e81 	:	val_out <= 4'h5367;
         4'h8e82 	:	val_out <= 4'h5367;
         4'h8e83 	:	val_out <= 4'h5367;
         4'h8e88 	:	val_out <= 4'h534f;
         4'h8e89 	:	val_out <= 4'h534f;
         4'h8e8a 	:	val_out <= 4'h534f;
         4'h8e8b 	:	val_out <= 4'h534f;
         4'h8e90 	:	val_out <= 4'h5337;
         4'h8e91 	:	val_out <= 4'h5337;
         4'h8e92 	:	val_out <= 4'h5337;
         4'h8e93 	:	val_out <= 4'h5337;
         4'h8e98 	:	val_out <= 4'h5320;
         4'h8e99 	:	val_out <= 4'h5320;
         4'h8e9a 	:	val_out <= 4'h5320;
         4'h8e9b 	:	val_out <= 4'h5320;
         4'h8ea0 	:	val_out <= 4'h5308;
         4'h8ea1 	:	val_out <= 4'h5308;
         4'h8ea2 	:	val_out <= 4'h5308;
         4'h8ea3 	:	val_out <= 4'h5308;
         4'h8ea8 	:	val_out <= 4'h52f1;
         4'h8ea9 	:	val_out <= 4'h52f1;
         4'h8eaa 	:	val_out <= 4'h52f1;
         4'h8eab 	:	val_out <= 4'h52f1;
         4'h8eb0 	:	val_out <= 4'h52d9;
         4'h8eb1 	:	val_out <= 4'h52d9;
         4'h8eb2 	:	val_out <= 4'h52d9;
         4'h8eb3 	:	val_out <= 4'h52d9;
         4'h8eb8 	:	val_out <= 4'h52c2;
         4'h8eb9 	:	val_out <= 4'h52c2;
         4'h8eba 	:	val_out <= 4'h52c2;
         4'h8ebb 	:	val_out <= 4'h52c2;
         4'h8ec0 	:	val_out <= 4'h52aa;
         4'h8ec1 	:	val_out <= 4'h52aa;
         4'h8ec2 	:	val_out <= 4'h52aa;
         4'h8ec3 	:	val_out <= 4'h52aa;
         4'h8ec8 	:	val_out <= 4'h5293;
         4'h8ec9 	:	val_out <= 4'h5293;
         4'h8eca 	:	val_out <= 4'h5293;
         4'h8ecb 	:	val_out <= 4'h5293;
         4'h8ed0 	:	val_out <= 4'h527b;
         4'h8ed1 	:	val_out <= 4'h527b;
         4'h8ed2 	:	val_out <= 4'h527b;
         4'h8ed3 	:	val_out <= 4'h527b;
         4'h8ed8 	:	val_out <= 4'h5264;
         4'h8ed9 	:	val_out <= 4'h5264;
         4'h8eda 	:	val_out <= 4'h5264;
         4'h8edb 	:	val_out <= 4'h5264;
         4'h8ee0 	:	val_out <= 4'h524c;
         4'h8ee1 	:	val_out <= 4'h524c;
         4'h8ee2 	:	val_out <= 4'h524c;
         4'h8ee3 	:	val_out <= 4'h524c;
         4'h8ee8 	:	val_out <= 4'h5235;
         4'h8ee9 	:	val_out <= 4'h5235;
         4'h8eea 	:	val_out <= 4'h5235;
         4'h8eeb 	:	val_out <= 4'h5235;
         4'h8ef0 	:	val_out <= 4'h521d;
         4'h8ef1 	:	val_out <= 4'h521d;
         4'h8ef2 	:	val_out <= 4'h521d;
         4'h8ef3 	:	val_out <= 4'h521d;
         4'h8ef8 	:	val_out <= 4'h5206;
         4'h8ef9 	:	val_out <= 4'h5206;
         4'h8efa 	:	val_out <= 4'h5206;
         4'h8efb 	:	val_out <= 4'h5206;
         4'h8f00 	:	val_out <= 4'h51ee;
         4'h8f01 	:	val_out <= 4'h51ee;
         4'h8f02 	:	val_out <= 4'h51ee;
         4'h8f03 	:	val_out <= 4'h51ee;
         4'h8f08 	:	val_out <= 4'h51d7;
         4'h8f09 	:	val_out <= 4'h51d7;
         4'h8f0a 	:	val_out <= 4'h51d7;
         4'h8f0b 	:	val_out <= 4'h51d7;
         4'h8f10 	:	val_out <= 4'h51c0;
         4'h8f11 	:	val_out <= 4'h51c0;
         4'h8f12 	:	val_out <= 4'h51c0;
         4'h8f13 	:	val_out <= 4'h51c0;
         4'h8f18 	:	val_out <= 4'h51a8;
         4'h8f19 	:	val_out <= 4'h51a8;
         4'h8f1a 	:	val_out <= 4'h51a8;
         4'h8f1b 	:	val_out <= 4'h51a8;
         4'h8f20 	:	val_out <= 4'h5191;
         4'h8f21 	:	val_out <= 4'h5191;
         4'h8f22 	:	val_out <= 4'h5191;
         4'h8f23 	:	val_out <= 4'h5191;
         4'h8f28 	:	val_out <= 4'h5179;
         4'h8f29 	:	val_out <= 4'h5179;
         4'h8f2a 	:	val_out <= 4'h5179;
         4'h8f2b 	:	val_out <= 4'h5179;
         4'h8f30 	:	val_out <= 4'h5162;
         4'h8f31 	:	val_out <= 4'h5162;
         4'h8f32 	:	val_out <= 4'h5162;
         4'h8f33 	:	val_out <= 4'h5162;
         4'h8f38 	:	val_out <= 4'h514a;
         4'h8f39 	:	val_out <= 4'h514a;
         4'h8f3a 	:	val_out <= 4'h514a;
         4'h8f3b 	:	val_out <= 4'h514a;
         4'h8f40 	:	val_out <= 4'h5133;
         4'h8f41 	:	val_out <= 4'h5133;
         4'h8f42 	:	val_out <= 4'h5133;
         4'h8f43 	:	val_out <= 4'h5133;
         4'h8f48 	:	val_out <= 4'h511c;
         4'h8f49 	:	val_out <= 4'h511c;
         4'h8f4a 	:	val_out <= 4'h511c;
         4'h8f4b 	:	val_out <= 4'h511c;
         4'h8f50 	:	val_out <= 4'h5104;
         4'h8f51 	:	val_out <= 4'h5104;
         4'h8f52 	:	val_out <= 4'h5104;
         4'h8f53 	:	val_out <= 4'h5104;
         4'h8f58 	:	val_out <= 4'h50ed;
         4'h8f59 	:	val_out <= 4'h50ed;
         4'h8f5a 	:	val_out <= 4'h50ed;
         4'h8f5b 	:	val_out <= 4'h50ed;
         4'h8f60 	:	val_out <= 4'h50d6;
         4'h8f61 	:	val_out <= 4'h50d6;
         4'h8f62 	:	val_out <= 4'h50d6;
         4'h8f63 	:	val_out <= 4'h50d6;
         4'h8f68 	:	val_out <= 4'h50be;
         4'h8f69 	:	val_out <= 4'h50be;
         4'h8f6a 	:	val_out <= 4'h50be;
         4'h8f6b 	:	val_out <= 4'h50be;
         4'h8f70 	:	val_out <= 4'h50a7;
         4'h8f71 	:	val_out <= 4'h50a7;
         4'h8f72 	:	val_out <= 4'h50a7;
         4'h8f73 	:	val_out <= 4'h50a7;
         4'h8f78 	:	val_out <= 4'h5090;
         4'h8f79 	:	val_out <= 4'h5090;
         4'h8f7a 	:	val_out <= 4'h5090;
         4'h8f7b 	:	val_out <= 4'h5090;
         4'h8f80 	:	val_out <= 4'h5078;
         4'h8f81 	:	val_out <= 4'h5078;
         4'h8f82 	:	val_out <= 4'h5078;
         4'h8f83 	:	val_out <= 4'h5078;
         4'h8f88 	:	val_out <= 4'h5061;
         4'h8f89 	:	val_out <= 4'h5061;
         4'h8f8a 	:	val_out <= 4'h5061;
         4'h8f8b 	:	val_out <= 4'h5061;
         4'h8f90 	:	val_out <= 4'h504a;
         4'h8f91 	:	val_out <= 4'h504a;
         4'h8f92 	:	val_out <= 4'h504a;
         4'h8f93 	:	val_out <= 4'h504a;
         4'h8f98 	:	val_out <= 4'h5032;
         4'h8f99 	:	val_out <= 4'h5032;
         4'h8f9a 	:	val_out <= 4'h5032;
         4'h8f9b 	:	val_out <= 4'h5032;
         4'h8fa0 	:	val_out <= 4'h501b;
         4'h8fa1 	:	val_out <= 4'h501b;
         4'h8fa2 	:	val_out <= 4'h501b;
         4'h8fa3 	:	val_out <= 4'h501b;
         4'h8fa8 	:	val_out <= 4'h5004;
         4'h8fa9 	:	val_out <= 4'h5004;
         4'h8faa 	:	val_out <= 4'h5004;
         4'h8fab 	:	val_out <= 4'h5004;
         4'h8fb0 	:	val_out <= 4'h4fec;
         4'h8fb1 	:	val_out <= 4'h4fec;
         4'h8fb2 	:	val_out <= 4'h4fec;
         4'h8fb3 	:	val_out <= 4'h4fec;
         4'h8fb8 	:	val_out <= 4'h4fd5;
         4'h8fb9 	:	val_out <= 4'h4fd5;
         4'h8fba 	:	val_out <= 4'h4fd5;
         4'h8fbb 	:	val_out <= 4'h4fd5;
         4'h8fc0 	:	val_out <= 4'h4fbe;
         4'h8fc1 	:	val_out <= 4'h4fbe;
         4'h8fc2 	:	val_out <= 4'h4fbe;
         4'h8fc3 	:	val_out <= 4'h4fbe;
         4'h8fc8 	:	val_out <= 4'h4fa6;
         4'h8fc9 	:	val_out <= 4'h4fa6;
         4'h8fca 	:	val_out <= 4'h4fa6;
         4'h8fcb 	:	val_out <= 4'h4fa6;
         4'h8fd0 	:	val_out <= 4'h4f8f;
         4'h8fd1 	:	val_out <= 4'h4f8f;
         4'h8fd2 	:	val_out <= 4'h4f8f;
         4'h8fd3 	:	val_out <= 4'h4f8f;
         4'h8fd8 	:	val_out <= 4'h4f78;
         4'h8fd9 	:	val_out <= 4'h4f78;
         4'h8fda 	:	val_out <= 4'h4f78;
         4'h8fdb 	:	val_out <= 4'h4f78;
         4'h8fe0 	:	val_out <= 4'h4f61;
         4'h8fe1 	:	val_out <= 4'h4f61;
         4'h8fe2 	:	val_out <= 4'h4f61;
         4'h8fe3 	:	val_out <= 4'h4f61;
         4'h8fe8 	:	val_out <= 4'h4f49;
         4'h8fe9 	:	val_out <= 4'h4f49;
         4'h8fea 	:	val_out <= 4'h4f49;
         4'h8feb 	:	val_out <= 4'h4f49;
         4'h8ff0 	:	val_out <= 4'h4f32;
         4'h8ff1 	:	val_out <= 4'h4f32;
         4'h8ff2 	:	val_out <= 4'h4f32;
         4'h8ff3 	:	val_out <= 4'h4f32;
         4'h8ff8 	:	val_out <= 4'h4f1b;
         4'h8ff9 	:	val_out <= 4'h4f1b;
         4'h8ffa 	:	val_out <= 4'h4f1b;
         4'h8ffb 	:	val_out <= 4'h4f1b;
         4'h9000 	:	val_out <= 4'h4f04;
         4'h9001 	:	val_out <= 4'h4f04;
         4'h9002 	:	val_out <= 4'h4f04;
         4'h9003 	:	val_out <= 4'h4f04;
         4'h9008 	:	val_out <= 4'h4eed;
         4'h9009 	:	val_out <= 4'h4eed;
         4'h900a 	:	val_out <= 4'h4eed;
         4'h900b 	:	val_out <= 4'h4eed;
         4'h9010 	:	val_out <= 4'h4ed5;
         4'h9011 	:	val_out <= 4'h4ed5;
         4'h9012 	:	val_out <= 4'h4ed5;
         4'h9013 	:	val_out <= 4'h4ed5;
         4'h9018 	:	val_out <= 4'h4ebe;
         4'h9019 	:	val_out <= 4'h4ebe;
         4'h901a 	:	val_out <= 4'h4ebe;
         4'h901b 	:	val_out <= 4'h4ebe;
         4'h9020 	:	val_out <= 4'h4ea7;
         4'h9021 	:	val_out <= 4'h4ea7;
         4'h9022 	:	val_out <= 4'h4ea7;
         4'h9023 	:	val_out <= 4'h4ea7;
         4'h9028 	:	val_out <= 4'h4e90;
         4'h9029 	:	val_out <= 4'h4e90;
         4'h902a 	:	val_out <= 4'h4e90;
         4'h902b 	:	val_out <= 4'h4e90;
         4'h9030 	:	val_out <= 4'h4e79;
         4'h9031 	:	val_out <= 4'h4e79;
         4'h9032 	:	val_out <= 4'h4e79;
         4'h9033 	:	val_out <= 4'h4e79;
         4'h9038 	:	val_out <= 4'h4e61;
         4'h9039 	:	val_out <= 4'h4e61;
         4'h903a 	:	val_out <= 4'h4e61;
         4'h903b 	:	val_out <= 4'h4e61;
         4'h9040 	:	val_out <= 4'h4e4a;
         4'h9041 	:	val_out <= 4'h4e4a;
         4'h9042 	:	val_out <= 4'h4e4a;
         4'h9043 	:	val_out <= 4'h4e4a;
         4'h9048 	:	val_out <= 4'h4e33;
         4'h9049 	:	val_out <= 4'h4e33;
         4'h904a 	:	val_out <= 4'h4e33;
         4'h904b 	:	val_out <= 4'h4e33;
         4'h9050 	:	val_out <= 4'h4e1c;
         4'h9051 	:	val_out <= 4'h4e1c;
         4'h9052 	:	val_out <= 4'h4e1c;
         4'h9053 	:	val_out <= 4'h4e1c;
         4'h9058 	:	val_out <= 4'h4e05;
         4'h9059 	:	val_out <= 4'h4e05;
         4'h905a 	:	val_out <= 4'h4e05;
         4'h905b 	:	val_out <= 4'h4e05;
         4'h9060 	:	val_out <= 4'h4dee;
         4'h9061 	:	val_out <= 4'h4dee;
         4'h9062 	:	val_out <= 4'h4dee;
         4'h9063 	:	val_out <= 4'h4dee;
         4'h9068 	:	val_out <= 4'h4dd7;
         4'h9069 	:	val_out <= 4'h4dd7;
         4'h906a 	:	val_out <= 4'h4dd7;
         4'h906b 	:	val_out <= 4'h4dd7;
         4'h9070 	:	val_out <= 4'h4dbf;
         4'h9071 	:	val_out <= 4'h4dbf;
         4'h9072 	:	val_out <= 4'h4dbf;
         4'h9073 	:	val_out <= 4'h4dbf;
         4'h9078 	:	val_out <= 4'h4da8;
         4'h9079 	:	val_out <= 4'h4da8;
         4'h907a 	:	val_out <= 4'h4da8;
         4'h907b 	:	val_out <= 4'h4da8;
         4'h9080 	:	val_out <= 4'h4d91;
         4'h9081 	:	val_out <= 4'h4d91;
         4'h9082 	:	val_out <= 4'h4d91;
         4'h9083 	:	val_out <= 4'h4d91;
         4'h9088 	:	val_out <= 4'h4d7a;
         4'h9089 	:	val_out <= 4'h4d7a;
         4'h908a 	:	val_out <= 4'h4d7a;
         4'h908b 	:	val_out <= 4'h4d7a;
         4'h9090 	:	val_out <= 4'h4d63;
         4'h9091 	:	val_out <= 4'h4d63;
         4'h9092 	:	val_out <= 4'h4d63;
         4'h9093 	:	val_out <= 4'h4d63;
         4'h9098 	:	val_out <= 4'h4d4c;
         4'h9099 	:	val_out <= 4'h4d4c;
         4'h909a 	:	val_out <= 4'h4d4c;
         4'h909b 	:	val_out <= 4'h4d4c;
         4'h90a0 	:	val_out <= 4'h4d35;
         4'h90a1 	:	val_out <= 4'h4d35;
         4'h90a2 	:	val_out <= 4'h4d35;
         4'h90a3 	:	val_out <= 4'h4d35;
         4'h90a8 	:	val_out <= 4'h4d1e;
         4'h90a9 	:	val_out <= 4'h4d1e;
         4'h90aa 	:	val_out <= 4'h4d1e;
         4'h90ab 	:	val_out <= 4'h4d1e;
         4'h90b0 	:	val_out <= 4'h4d07;
         4'h90b1 	:	val_out <= 4'h4d07;
         4'h90b2 	:	val_out <= 4'h4d07;
         4'h90b3 	:	val_out <= 4'h4d07;
         4'h90b8 	:	val_out <= 4'h4cf0;
         4'h90b9 	:	val_out <= 4'h4cf0;
         4'h90ba 	:	val_out <= 4'h4cf0;
         4'h90bb 	:	val_out <= 4'h4cf0;
         4'h90c0 	:	val_out <= 4'h4cd9;
         4'h90c1 	:	val_out <= 4'h4cd9;
         4'h90c2 	:	val_out <= 4'h4cd9;
         4'h90c3 	:	val_out <= 4'h4cd9;
         4'h90c8 	:	val_out <= 4'h4cc2;
         4'h90c9 	:	val_out <= 4'h4cc2;
         4'h90ca 	:	val_out <= 4'h4cc2;
         4'h90cb 	:	val_out <= 4'h4cc2;
         4'h90d0 	:	val_out <= 4'h4cab;
         4'h90d1 	:	val_out <= 4'h4cab;
         4'h90d2 	:	val_out <= 4'h4cab;
         4'h90d3 	:	val_out <= 4'h4cab;
         4'h90d8 	:	val_out <= 4'h4c94;
         4'h90d9 	:	val_out <= 4'h4c94;
         4'h90da 	:	val_out <= 4'h4c94;
         4'h90db 	:	val_out <= 4'h4c94;
         4'h90e0 	:	val_out <= 4'h4c7d;
         4'h90e1 	:	val_out <= 4'h4c7d;
         4'h90e2 	:	val_out <= 4'h4c7d;
         4'h90e3 	:	val_out <= 4'h4c7d;
         4'h90e8 	:	val_out <= 4'h4c66;
         4'h90e9 	:	val_out <= 4'h4c66;
         4'h90ea 	:	val_out <= 4'h4c66;
         4'h90eb 	:	val_out <= 4'h4c66;
         4'h90f0 	:	val_out <= 4'h4c4f;
         4'h90f1 	:	val_out <= 4'h4c4f;
         4'h90f2 	:	val_out <= 4'h4c4f;
         4'h90f3 	:	val_out <= 4'h4c4f;
         4'h90f8 	:	val_out <= 4'h4c38;
         4'h90f9 	:	val_out <= 4'h4c38;
         4'h90fa 	:	val_out <= 4'h4c38;
         4'h90fb 	:	val_out <= 4'h4c38;
         4'h9100 	:	val_out <= 4'h4c21;
         4'h9101 	:	val_out <= 4'h4c21;
         4'h9102 	:	val_out <= 4'h4c21;
         4'h9103 	:	val_out <= 4'h4c21;
         4'h9108 	:	val_out <= 4'h4c0a;
         4'h9109 	:	val_out <= 4'h4c0a;
         4'h910a 	:	val_out <= 4'h4c0a;
         4'h910b 	:	val_out <= 4'h4c0a;
         4'h9110 	:	val_out <= 4'h4bf3;
         4'h9111 	:	val_out <= 4'h4bf3;
         4'h9112 	:	val_out <= 4'h4bf3;
         4'h9113 	:	val_out <= 4'h4bf3;
         4'h9118 	:	val_out <= 4'h4bdc;
         4'h9119 	:	val_out <= 4'h4bdc;
         4'h911a 	:	val_out <= 4'h4bdc;
         4'h911b 	:	val_out <= 4'h4bdc;
         4'h9120 	:	val_out <= 4'h4bc5;
         4'h9121 	:	val_out <= 4'h4bc5;
         4'h9122 	:	val_out <= 4'h4bc5;
         4'h9123 	:	val_out <= 4'h4bc5;
         4'h9128 	:	val_out <= 4'h4bae;
         4'h9129 	:	val_out <= 4'h4bae;
         4'h912a 	:	val_out <= 4'h4bae;
         4'h912b 	:	val_out <= 4'h4bae;
         4'h9130 	:	val_out <= 4'h4b97;
         4'h9131 	:	val_out <= 4'h4b97;
         4'h9132 	:	val_out <= 4'h4b97;
         4'h9133 	:	val_out <= 4'h4b97;
         4'h9138 	:	val_out <= 4'h4b80;
         4'h9139 	:	val_out <= 4'h4b80;
         4'h913a 	:	val_out <= 4'h4b80;
         4'h913b 	:	val_out <= 4'h4b80;
         4'h9140 	:	val_out <= 4'h4b69;
         4'h9141 	:	val_out <= 4'h4b69;
         4'h9142 	:	val_out <= 4'h4b69;
         4'h9143 	:	val_out <= 4'h4b69;
         4'h9148 	:	val_out <= 4'h4b52;
         4'h9149 	:	val_out <= 4'h4b52;
         4'h914a 	:	val_out <= 4'h4b52;
         4'h914b 	:	val_out <= 4'h4b52;
         4'h9150 	:	val_out <= 4'h4b3b;
         4'h9151 	:	val_out <= 4'h4b3b;
         4'h9152 	:	val_out <= 4'h4b3b;
         4'h9153 	:	val_out <= 4'h4b3b;
         4'h9158 	:	val_out <= 4'h4b24;
         4'h9159 	:	val_out <= 4'h4b24;
         4'h915a 	:	val_out <= 4'h4b24;
         4'h915b 	:	val_out <= 4'h4b24;
         4'h9160 	:	val_out <= 4'h4b0d;
         4'h9161 	:	val_out <= 4'h4b0d;
         4'h9162 	:	val_out <= 4'h4b0d;
         4'h9163 	:	val_out <= 4'h4b0d;
         4'h9168 	:	val_out <= 4'h4af7;
         4'h9169 	:	val_out <= 4'h4af7;
         4'h916a 	:	val_out <= 4'h4af7;
         4'h916b 	:	val_out <= 4'h4af7;
         4'h9170 	:	val_out <= 4'h4ae0;
         4'h9171 	:	val_out <= 4'h4ae0;
         4'h9172 	:	val_out <= 4'h4ae0;
         4'h9173 	:	val_out <= 4'h4ae0;
         4'h9178 	:	val_out <= 4'h4ac9;
         4'h9179 	:	val_out <= 4'h4ac9;
         4'h917a 	:	val_out <= 4'h4ac9;
         4'h917b 	:	val_out <= 4'h4ac9;
         4'h9180 	:	val_out <= 4'h4ab2;
         4'h9181 	:	val_out <= 4'h4ab2;
         4'h9182 	:	val_out <= 4'h4ab2;
         4'h9183 	:	val_out <= 4'h4ab2;
         4'h9188 	:	val_out <= 4'h4a9b;
         4'h9189 	:	val_out <= 4'h4a9b;
         4'h918a 	:	val_out <= 4'h4a9b;
         4'h918b 	:	val_out <= 4'h4a9b;
         4'h9190 	:	val_out <= 4'h4a84;
         4'h9191 	:	val_out <= 4'h4a84;
         4'h9192 	:	val_out <= 4'h4a84;
         4'h9193 	:	val_out <= 4'h4a84;
         4'h9198 	:	val_out <= 4'h4a6d;
         4'h9199 	:	val_out <= 4'h4a6d;
         4'h919a 	:	val_out <= 4'h4a6d;
         4'h919b 	:	val_out <= 4'h4a6d;
         4'h91a0 	:	val_out <= 4'h4a57;
         4'h91a1 	:	val_out <= 4'h4a57;
         4'h91a2 	:	val_out <= 4'h4a57;
         4'h91a3 	:	val_out <= 4'h4a57;
         4'h91a8 	:	val_out <= 4'h4a40;
         4'h91a9 	:	val_out <= 4'h4a40;
         4'h91aa 	:	val_out <= 4'h4a40;
         4'h91ab 	:	val_out <= 4'h4a40;
         4'h91b0 	:	val_out <= 4'h4a29;
         4'h91b1 	:	val_out <= 4'h4a29;
         4'h91b2 	:	val_out <= 4'h4a29;
         4'h91b3 	:	val_out <= 4'h4a29;
         4'h91b8 	:	val_out <= 4'h4a12;
         4'h91b9 	:	val_out <= 4'h4a12;
         4'h91ba 	:	val_out <= 4'h4a12;
         4'h91bb 	:	val_out <= 4'h4a12;
         4'h91c0 	:	val_out <= 4'h49fb;
         4'h91c1 	:	val_out <= 4'h49fb;
         4'h91c2 	:	val_out <= 4'h49fb;
         4'h91c3 	:	val_out <= 4'h49fb;
         4'h91c8 	:	val_out <= 4'h49e5;
         4'h91c9 	:	val_out <= 4'h49e5;
         4'h91ca 	:	val_out <= 4'h49e5;
         4'h91cb 	:	val_out <= 4'h49e5;
         4'h91d0 	:	val_out <= 4'h49ce;
         4'h91d1 	:	val_out <= 4'h49ce;
         4'h91d2 	:	val_out <= 4'h49ce;
         4'h91d3 	:	val_out <= 4'h49ce;
         4'h91d8 	:	val_out <= 4'h49b7;
         4'h91d9 	:	val_out <= 4'h49b7;
         4'h91da 	:	val_out <= 4'h49b7;
         4'h91db 	:	val_out <= 4'h49b7;
         4'h91e0 	:	val_out <= 4'h49a0;
         4'h91e1 	:	val_out <= 4'h49a0;
         4'h91e2 	:	val_out <= 4'h49a0;
         4'h91e3 	:	val_out <= 4'h49a0;
         4'h91e8 	:	val_out <= 4'h498a;
         4'h91e9 	:	val_out <= 4'h498a;
         4'h91ea 	:	val_out <= 4'h498a;
         4'h91eb 	:	val_out <= 4'h498a;
         4'h91f0 	:	val_out <= 4'h4973;
         4'h91f1 	:	val_out <= 4'h4973;
         4'h91f2 	:	val_out <= 4'h4973;
         4'h91f3 	:	val_out <= 4'h4973;
         4'h91f8 	:	val_out <= 4'h495c;
         4'h91f9 	:	val_out <= 4'h495c;
         4'h91fa 	:	val_out <= 4'h495c;
         4'h91fb 	:	val_out <= 4'h495c;
         4'h9200 	:	val_out <= 4'h4945;
         4'h9201 	:	val_out <= 4'h4945;
         4'h9202 	:	val_out <= 4'h4945;
         4'h9203 	:	val_out <= 4'h4945;
         4'h9208 	:	val_out <= 4'h492f;
         4'h9209 	:	val_out <= 4'h492f;
         4'h920a 	:	val_out <= 4'h492f;
         4'h920b 	:	val_out <= 4'h492f;
         4'h9210 	:	val_out <= 4'h4918;
         4'h9211 	:	val_out <= 4'h4918;
         4'h9212 	:	val_out <= 4'h4918;
         4'h9213 	:	val_out <= 4'h4918;
         4'h9218 	:	val_out <= 4'h4901;
         4'h9219 	:	val_out <= 4'h4901;
         4'h921a 	:	val_out <= 4'h4901;
         4'h921b 	:	val_out <= 4'h4901;
         4'h9220 	:	val_out <= 4'h48eb;
         4'h9221 	:	val_out <= 4'h48eb;
         4'h9222 	:	val_out <= 4'h48eb;
         4'h9223 	:	val_out <= 4'h48eb;
         4'h9228 	:	val_out <= 4'h48d4;
         4'h9229 	:	val_out <= 4'h48d4;
         4'h922a 	:	val_out <= 4'h48d4;
         4'h922b 	:	val_out <= 4'h48d4;
         4'h9230 	:	val_out <= 4'h48bd;
         4'h9231 	:	val_out <= 4'h48bd;
         4'h9232 	:	val_out <= 4'h48bd;
         4'h9233 	:	val_out <= 4'h48bd;
         4'h9238 	:	val_out <= 4'h48a7;
         4'h9239 	:	val_out <= 4'h48a7;
         4'h923a 	:	val_out <= 4'h48a7;
         4'h923b 	:	val_out <= 4'h48a7;
         4'h9240 	:	val_out <= 4'h4890;
         4'h9241 	:	val_out <= 4'h4890;
         4'h9242 	:	val_out <= 4'h4890;
         4'h9243 	:	val_out <= 4'h4890;
         4'h9248 	:	val_out <= 4'h4879;
         4'h9249 	:	val_out <= 4'h4879;
         4'h924a 	:	val_out <= 4'h4879;
         4'h924b 	:	val_out <= 4'h4879;
         4'h9250 	:	val_out <= 4'h4863;
         4'h9251 	:	val_out <= 4'h4863;
         4'h9252 	:	val_out <= 4'h4863;
         4'h9253 	:	val_out <= 4'h4863;
         4'h9258 	:	val_out <= 4'h484c;
         4'h9259 	:	val_out <= 4'h484c;
         4'h925a 	:	val_out <= 4'h484c;
         4'h925b 	:	val_out <= 4'h484c;
         4'h9260 	:	val_out <= 4'h4835;
         4'h9261 	:	val_out <= 4'h4835;
         4'h9262 	:	val_out <= 4'h4835;
         4'h9263 	:	val_out <= 4'h4835;
         4'h9268 	:	val_out <= 4'h481f;
         4'h9269 	:	val_out <= 4'h481f;
         4'h926a 	:	val_out <= 4'h481f;
         4'h926b 	:	val_out <= 4'h481f;
         4'h9270 	:	val_out <= 4'h4808;
         4'h9271 	:	val_out <= 4'h4808;
         4'h9272 	:	val_out <= 4'h4808;
         4'h9273 	:	val_out <= 4'h4808;
         4'h9278 	:	val_out <= 4'h47f2;
         4'h9279 	:	val_out <= 4'h47f2;
         4'h927a 	:	val_out <= 4'h47f2;
         4'h927b 	:	val_out <= 4'h47f2;
         4'h9280 	:	val_out <= 4'h47db;
         4'h9281 	:	val_out <= 4'h47db;
         4'h9282 	:	val_out <= 4'h47db;
         4'h9283 	:	val_out <= 4'h47db;
         4'h9288 	:	val_out <= 4'h47c4;
         4'h9289 	:	val_out <= 4'h47c4;
         4'h928a 	:	val_out <= 4'h47c4;
         4'h928b 	:	val_out <= 4'h47c4;
         4'h9290 	:	val_out <= 4'h47ae;
         4'h9291 	:	val_out <= 4'h47ae;
         4'h9292 	:	val_out <= 4'h47ae;
         4'h9293 	:	val_out <= 4'h47ae;
         4'h9298 	:	val_out <= 4'h4797;
         4'h9299 	:	val_out <= 4'h4797;
         4'h929a 	:	val_out <= 4'h4797;
         4'h929b 	:	val_out <= 4'h4797;
         4'h92a0 	:	val_out <= 4'h4781;
         4'h92a1 	:	val_out <= 4'h4781;
         4'h92a2 	:	val_out <= 4'h4781;
         4'h92a3 	:	val_out <= 4'h4781;
         4'h92a8 	:	val_out <= 4'h476a;
         4'h92a9 	:	val_out <= 4'h476a;
         4'h92aa 	:	val_out <= 4'h476a;
         4'h92ab 	:	val_out <= 4'h476a;
         4'h92b0 	:	val_out <= 4'h4754;
         4'h92b1 	:	val_out <= 4'h4754;
         4'h92b2 	:	val_out <= 4'h4754;
         4'h92b3 	:	val_out <= 4'h4754;
         4'h92b8 	:	val_out <= 4'h473d;
         4'h92b9 	:	val_out <= 4'h473d;
         4'h92ba 	:	val_out <= 4'h473d;
         4'h92bb 	:	val_out <= 4'h473d;
         4'h92c0 	:	val_out <= 4'h4727;
         4'h92c1 	:	val_out <= 4'h4727;
         4'h92c2 	:	val_out <= 4'h4727;
         4'h92c3 	:	val_out <= 4'h4727;
         4'h92c8 	:	val_out <= 4'h4710;
         4'h92c9 	:	val_out <= 4'h4710;
         4'h92ca 	:	val_out <= 4'h4710;
         4'h92cb 	:	val_out <= 4'h4710;
         4'h92d0 	:	val_out <= 4'h46f9;
         4'h92d1 	:	val_out <= 4'h46f9;
         4'h92d2 	:	val_out <= 4'h46f9;
         4'h92d3 	:	val_out <= 4'h46f9;
         4'h92d8 	:	val_out <= 4'h46e3;
         4'h92d9 	:	val_out <= 4'h46e3;
         4'h92da 	:	val_out <= 4'h46e3;
         4'h92db 	:	val_out <= 4'h46e3;
         4'h92e0 	:	val_out <= 4'h46cd;
         4'h92e1 	:	val_out <= 4'h46cd;
         4'h92e2 	:	val_out <= 4'h46cd;
         4'h92e3 	:	val_out <= 4'h46cd;
         4'h92e8 	:	val_out <= 4'h46b6;
         4'h92e9 	:	val_out <= 4'h46b6;
         4'h92ea 	:	val_out <= 4'h46b6;
         4'h92eb 	:	val_out <= 4'h46b6;
         4'h92f0 	:	val_out <= 4'h46a0;
         4'h92f1 	:	val_out <= 4'h46a0;
         4'h92f2 	:	val_out <= 4'h46a0;
         4'h92f3 	:	val_out <= 4'h46a0;
         4'h92f8 	:	val_out <= 4'h4689;
         4'h92f9 	:	val_out <= 4'h4689;
         4'h92fa 	:	val_out <= 4'h4689;
         4'h92fb 	:	val_out <= 4'h4689;
         4'h9300 	:	val_out <= 4'h4673;
         4'h9301 	:	val_out <= 4'h4673;
         4'h9302 	:	val_out <= 4'h4673;
         4'h9303 	:	val_out <= 4'h4673;
         4'h9308 	:	val_out <= 4'h465c;
         4'h9309 	:	val_out <= 4'h465c;
         4'h930a 	:	val_out <= 4'h465c;
         4'h930b 	:	val_out <= 4'h465c;
         4'h9310 	:	val_out <= 4'h4646;
         4'h9311 	:	val_out <= 4'h4646;
         4'h9312 	:	val_out <= 4'h4646;
         4'h9313 	:	val_out <= 4'h4646;
         4'h9318 	:	val_out <= 4'h462f;
         4'h9319 	:	val_out <= 4'h462f;
         4'h931a 	:	val_out <= 4'h462f;
         4'h931b 	:	val_out <= 4'h462f;
         4'h9320 	:	val_out <= 4'h4619;
         4'h9321 	:	val_out <= 4'h4619;
         4'h9322 	:	val_out <= 4'h4619;
         4'h9323 	:	val_out <= 4'h4619;
         4'h9328 	:	val_out <= 4'h4602;
         4'h9329 	:	val_out <= 4'h4602;
         4'h932a 	:	val_out <= 4'h4602;
         4'h932b 	:	val_out <= 4'h4602;
         4'h9330 	:	val_out <= 4'h45ec;
         4'h9331 	:	val_out <= 4'h45ec;
         4'h9332 	:	val_out <= 4'h45ec;
         4'h9333 	:	val_out <= 4'h45ec;
         4'h9338 	:	val_out <= 4'h45d6;
         4'h9339 	:	val_out <= 4'h45d6;
         4'h933a 	:	val_out <= 4'h45d6;
         4'h933b 	:	val_out <= 4'h45d6;
         4'h9340 	:	val_out <= 4'h45bf;
         4'h9341 	:	val_out <= 4'h45bf;
         4'h9342 	:	val_out <= 4'h45bf;
         4'h9343 	:	val_out <= 4'h45bf;
         4'h9348 	:	val_out <= 4'h45a9;
         4'h9349 	:	val_out <= 4'h45a9;
         4'h934a 	:	val_out <= 4'h45a9;
         4'h934b 	:	val_out <= 4'h45a9;
         4'h9350 	:	val_out <= 4'h4593;
         4'h9351 	:	val_out <= 4'h4593;
         4'h9352 	:	val_out <= 4'h4593;
         4'h9353 	:	val_out <= 4'h4593;
         4'h9358 	:	val_out <= 4'h457c;
         4'h9359 	:	val_out <= 4'h457c;
         4'h935a 	:	val_out <= 4'h457c;
         4'h935b 	:	val_out <= 4'h457c;
         4'h9360 	:	val_out <= 4'h4566;
         4'h9361 	:	val_out <= 4'h4566;
         4'h9362 	:	val_out <= 4'h4566;
         4'h9363 	:	val_out <= 4'h4566;
         4'h9368 	:	val_out <= 4'h4550;
         4'h9369 	:	val_out <= 4'h4550;
         4'h936a 	:	val_out <= 4'h4550;
         4'h936b 	:	val_out <= 4'h4550;
         4'h9370 	:	val_out <= 4'h4539;
         4'h9371 	:	val_out <= 4'h4539;
         4'h9372 	:	val_out <= 4'h4539;
         4'h9373 	:	val_out <= 4'h4539;
         4'h9378 	:	val_out <= 4'h4523;
         4'h9379 	:	val_out <= 4'h4523;
         4'h937a 	:	val_out <= 4'h4523;
         4'h937b 	:	val_out <= 4'h4523;
         4'h9380 	:	val_out <= 4'h450d;
         4'h9381 	:	val_out <= 4'h450d;
         4'h9382 	:	val_out <= 4'h450d;
         4'h9383 	:	val_out <= 4'h450d;
         4'h9388 	:	val_out <= 4'h44f6;
         4'h9389 	:	val_out <= 4'h44f6;
         4'h938a 	:	val_out <= 4'h44f6;
         4'h938b 	:	val_out <= 4'h44f6;
         4'h9390 	:	val_out <= 4'h44e0;
         4'h9391 	:	val_out <= 4'h44e0;
         4'h9392 	:	val_out <= 4'h44e0;
         4'h9393 	:	val_out <= 4'h44e0;
         4'h9398 	:	val_out <= 4'h44ca;
         4'h9399 	:	val_out <= 4'h44ca;
         4'h939a 	:	val_out <= 4'h44ca;
         4'h939b 	:	val_out <= 4'h44ca;
         4'h93a0 	:	val_out <= 4'h44b3;
         4'h93a1 	:	val_out <= 4'h44b3;
         4'h93a2 	:	val_out <= 4'h44b3;
         4'h93a3 	:	val_out <= 4'h44b3;
         4'h93a8 	:	val_out <= 4'h449d;
         4'h93a9 	:	val_out <= 4'h449d;
         4'h93aa 	:	val_out <= 4'h449d;
         4'h93ab 	:	val_out <= 4'h449d;
         4'h93b0 	:	val_out <= 4'h4487;
         4'h93b1 	:	val_out <= 4'h4487;
         4'h93b2 	:	val_out <= 4'h4487;
         4'h93b3 	:	val_out <= 4'h4487;
         4'h93b8 	:	val_out <= 4'h4471;
         4'h93b9 	:	val_out <= 4'h4471;
         4'h93ba 	:	val_out <= 4'h4471;
         4'h93bb 	:	val_out <= 4'h4471;
         4'h93c0 	:	val_out <= 4'h445a;
         4'h93c1 	:	val_out <= 4'h445a;
         4'h93c2 	:	val_out <= 4'h445a;
         4'h93c3 	:	val_out <= 4'h445a;
         4'h93c8 	:	val_out <= 4'h4444;
         4'h93c9 	:	val_out <= 4'h4444;
         4'h93ca 	:	val_out <= 4'h4444;
         4'h93cb 	:	val_out <= 4'h4444;
         4'h93d0 	:	val_out <= 4'h442e;
         4'h93d1 	:	val_out <= 4'h442e;
         4'h93d2 	:	val_out <= 4'h442e;
         4'h93d3 	:	val_out <= 4'h442e;
         4'h93d8 	:	val_out <= 4'h4418;
         4'h93d9 	:	val_out <= 4'h4418;
         4'h93da 	:	val_out <= 4'h4418;
         4'h93db 	:	val_out <= 4'h4418;
         4'h93e0 	:	val_out <= 4'h4402;
         4'h93e1 	:	val_out <= 4'h4402;
         4'h93e2 	:	val_out <= 4'h4402;
         4'h93e3 	:	val_out <= 4'h4402;
         4'h93e8 	:	val_out <= 4'h43eb;
         4'h93e9 	:	val_out <= 4'h43eb;
         4'h93ea 	:	val_out <= 4'h43eb;
         4'h93eb 	:	val_out <= 4'h43eb;
         4'h93f0 	:	val_out <= 4'h43d5;
         4'h93f1 	:	val_out <= 4'h43d5;
         4'h93f2 	:	val_out <= 4'h43d5;
         4'h93f3 	:	val_out <= 4'h43d5;
         4'h93f8 	:	val_out <= 4'h43bf;
         4'h93f9 	:	val_out <= 4'h43bf;
         4'h93fa 	:	val_out <= 4'h43bf;
         4'h93fb 	:	val_out <= 4'h43bf;
         4'h9400 	:	val_out <= 4'h43a9;
         4'h9401 	:	val_out <= 4'h43a9;
         4'h9402 	:	val_out <= 4'h43a9;
         4'h9403 	:	val_out <= 4'h43a9;
         4'h9408 	:	val_out <= 4'h4393;
         4'h9409 	:	val_out <= 4'h4393;
         4'h940a 	:	val_out <= 4'h4393;
         4'h940b 	:	val_out <= 4'h4393;
         4'h9410 	:	val_out <= 4'h437c;
         4'h9411 	:	val_out <= 4'h437c;
         4'h9412 	:	val_out <= 4'h437c;
         4'h9413 	:	val_out <= 4'h437c;
         4'h9418 	:	val_out <= 4'h4366;
         4'h9419 	:	val_out <= 4'h4366;
         4'h941a 	:	val_out <= 4'h4366;
         4'h941b 	:	val_out <= 4'h4366;
         4'h9420 	:	val_out <= 4'h4350;
         4'h9421 	:	val_out <= 4'h4350;
         4'h9422 	:	val_out <= 4'h4350;
         4'h9423 	:	val_out <= 4'h4350;
         4'h9428 	:	val_out <= 4'h433a;
         4'h9429 	:	val_out <= 4'h433a;
         4'h942a 	:	val_out <= 4'h433a;
         4'h942b 	:	val_out <= 4'h433a;
         4'h9430 	:	val_out <= 4'h4324;
         4'h9431 	:	val_out <= 4'h4324;
         4'h9432 	:	val_out <= 4'h4324;
         4'h9433 	:	val_out <= 4'h4324;
         4'h9438 	:	val_out <= 4'h430e;
         4'h9439 	:	val_out <= 4'h430e;
         4'h943a 	:	val_out <= 4'h430e;
         4'h943b 	:	val_out <= 4'h430e;
         4'h9440 	:	val_out <= 4'h42f8;
         4'h9441 	:	val_out <= 4'h42f8;
         4'h9442 	:	val_out <= 4'h42f8;
         4'h9443 	:	val_out <= 4'h42f8;
         4'h9448 	:	val_out <= 4'h42e2;
         4'h9449 	:	val_out <= 4'h42e2;
         4'h944a 	:	val_out <= 4'h42e2;
         4'h944b 	:	val_out <= 4'h42e2;
         4'h9450 	:	val_out <= 4'h42cc;
         4'h9451 	:	val_out <= 4'h42cc;
         4'h9452 	:	val_out <= 4'h42cc;
         4'h9453 	:	val_out <= 4'h42cc;
         4'h9458 	:	val_out <= 4'h42b6;
         4'h9459 	:	val_out <= 4'h42b6;
         4'h945a 	:	val_out <= 4'h42b6;
         4'h945b 	:	val_out <= 4'h42b6;
         4'h9460 	:	val_out <= 4'h429f;
         4'h9461 	:	val_out <= 4'h429f;
         4'h9462 	:	val_out <= 4'h429f;
         4'h9463 	:	val_out <= 4'h429f;
         4'h9468 	:	val_out <= 4'h4289;
         4'h9469 	:	val_out <= 4'h4289;
         4'h946a 	:	val_out <= 4'h4289;
         4'h946b 	:	val_out <= 4'h4289;
         4'h9470 	:	val_out <= 4'h4273;
         4'h9471 	:	val_out <= 4'h4273;
         4'h9472 	:	val_out <= 4'h4273;
         4'h9473 	:	val_out <= 4'h4273;
         4'h9478 	:	val_out <= 4'h425d;
         4'h9479 	:	val_out <= 4'h425d;
         4'h947a 	:	val_out <= 4'h425d;
         4'h947b 	:	val_out <= 4'h425d;
         4'h9480 	:	val_out <= 4'h4247;
         4'h9481 	:	val_out <= 4'h4247;
         4'h9482 	:	val_out <= 4'h4247;
         4'h9483 	:	val_out <= 4'h4247;
         4'h9488 	:	val_out <= 4'h4231;
         4'h9489 	:	val_out <= 4'h4231;
         4'h948a 	:	val_out <= 4'h4231;
         4'h948b 	:	val_out <= 4'h4231;
         4'h9490 	:	val_out <= 4'h421b;
         4'h9491 	:	val_out <= 4'h421b;
         4'h9492 	:	val_out <= 4'h421b;
         4'h9493 	:	val_out <= 4'h421b;
         4'h9498 	:	val_out <= 4'h4205;
         4'h9499 	:	val_out <= 4'h4205;
         4'h949a 	:	val_out <= 4'h4205;
         4'h949b 	:	val_out <= 4'h4205;
         4'h94a0 	:	val_out <= 4'h41ef;
         4'h94a1 	:	val_out <= 4'h41ef;
         4'h94a2 	:	val_out <= 4'h41ef;
         4'h94a3 	:	val_out <= 4'h41ef;
         4'h94a8 	:	val_out <= 4'h41d9;
         4'h94a9 	:	val_out <= 4'h41d9;
         4'h94aa 	:	val_out <= 4'h41d9;
         4'h94ab 	:	val_out <= 4'h41d9;
         4'h94b0 	:	val_out <= 4'h41c3;
         4'h94b1 	:	val_out <= 4'h41c3;
         4'h94b2 	:	val_out <= 4'h41c3;
         4'h94b3 	:	val_out <= 4'h41c3;
         4'h94b8 	:	val_out <= 4'h41ad;
         4'h94b9 	:	val_out <= 4'h41ad;
         4'h94ba 	:	val_out <= 4'h41ad;
         4'h94bb 	:	val_out <= 4'h41ad;
         4'h94c0 	:	val_out <= 4'h4197;
         4'h94c1 	:	val_out <= 4'h4197;
         4'h94c2 	:	val_out <= 4'h4197;
         4'h94c3 	:	val_out <= 4'h4197;
         4'h94c8 	:	val_out <= 4'h4182;
         4'h94c9 	:	val_out <= 4'h4182;
         4'h94ca 	:	val_out <= 4'h4182;
         4'h94cb 	:	val_out <= 4'h4182;
         4'h94d0 	:	val_out <= 4'h416c;
         4'h94d1 	:	val_out <= 4'h416c;
         4'h94d2 	:	val_out <= 4'h416c;
         4'h94d3 	:	val_out <= 4'h416c;
         4'h94d8 	:	val_out <= 4'h4156;
         4'h94d9 	:	val_out <= 4'h4156;
         4'h94da 	:	val_out <= 4'h4156;
         4'h94db 	:	val_out <= 4'h4156;
         4'h94e0 	:	val_out <= 4'h4140;
         4'h94e1 	:	val_out <= 4'h4140;
         4'h94e2 	:	val_out <= 4'h4140;
         4'h94e3 	:	val_out <= 4'h4140;
         4'h94e8 	:	val_out <= 4'h412a;
         4'h94e9 	:	val_out <= 4'h412a;
         4'h94ea 	:	val_out <= 4'h412a;
         4'h94eb 	:	val_out <= 4'h412a;
         4'h94f0 	:	val_out <= 4'h4114;
         4'h94f1 	:	val_out <= 4'h4114;
         4'h94f2 	:	val_out <= 4'h4114;
         4'h94f3 	:	val_out <= 4'h4114;
         4'h94f8 	:	val_out <= 4'h40fe;
         4'h94f9 	:	val_out <= 4'h40fe;
         4'h94fa 	:	val_out <= 4'h40fe;
         4'h94fb 	:	val_out <= 4'h40fe;
         4'h9500 	:	val_out <= 4'h40e8;
         4'h9501 	:	val_out <= 4'h40e8;
         4'h9502 	:	val_out <= 4'h40e8;
         4'h9503 	:	val_out <= 4'h40e8;
         4'h9508 	:	val_out <= 4'h40d2;
         4'h9509 	:	val_out <= 4'h40d2;
         4'h950a 	:	val_out <= 4'h40d2;
         4'h950b 	:	val_out <= 4'h40d2;
         4'h9510 	:	val_out <= 4'h40bc;
         4'h9511 	:	val_out <= 4'h40bc;
         4'h9512 	:	val_out <= 4'h40bc;
         4'h9513 	:	val_out <= 4'h40bc;
         4'h9518 	:	val_out <= 4'h40a7;
         4'h9519 	:	val_out <= 4'h40a7;
         4'h951a 	:	val_out <= 4'h40a7;
         4'h951b 	:	val_out <= 4'h40a7;
         4'h9520 	:	val_out <= 4'h4091;
         4'h9521 	:	val_out <= 4'h4091;
         4'h9522 	:	val_out <= 4'h4091;
         4'h9523 	:	val_out <= 4'h4091;
         4'h9528 	:	val_out <= 4'h407b;
         4'h9529 	:	val_out <= 4'h407b;
         4'h952a 	:	val_out <= 4'h407b;
         4'h952b 	:	val_out <= 4'h407b;
         4'h9530 	:	val_out <= 4'h4065;
         4'h9531 	:	val_out <= 4'h4065;
         4'h9532 	:	val_out <= 4'h4065;
         4'h9533 	:	val_out <= 4'h4065;
         4'h9538 	:	val_out <= 4'h404f;
         4'h9539 	:	val_out <= 4'h404f;
         4'h953a 	:	val_out <= 4'h404f;
         4'h953b 	:	val_out <= 4'h404f;
         4'h9540 	:	val_out <= 4'h403a;
         4'h9541 	:	val_out <= 4'h403a;
         4'h9542 	:	val_out <= 4'h403a;
         4'h9543 	:	val_out <= 4'h403a;
         4'h9548 	:	val_out <= 4'h4024;
         4'h9549 	:	val_out <= 4'h4024;
         4'h954a 	:	val_out <= 4'h4024;
         4'h954b 	:	val_out <= 4'h4024;
         4'h9550 	:	val_out <= 4'h400e;
         4'h9551 	:	val_out <= 4'h400e;
         4'h9552 	:	val_out <= 4'h400e;
         4'h9553 	:	val_out <= 4'h400e;
         4'h9558 	:	val_out <= 4'h3ff8;
         4'h9559 	:	val_out <= 4'h3ff8;
         4'h955a 	:	val_out <= 4'h3ff8;
         4'h955b 	:	val_out <= 4'h3ff8;
         4'h9560 	:	val_out <= 4'h3fe2;
         4'h9561 	:	val_out <= 4'h3fe2;
         4'h9562 	:	val_out <= 4'h3fe2;
         4'h9563 	:	val_out <= 4'h3fe2;
         4'h9568 	:	val_out <= 4'h3fcd;
         4'h9569 	:	val_out <= 4'h3fcd;
         4'h956a 	:	val_out <= 4'h3fcd;
         4'h956b 	:	val_out <= 4'h3fcd;
         4'h9570 	:	val_out <= 4'h3fb7;
         4'h9571 	:	val_out <= 4'h3fb7;
         4'h9572 	:	val_out <= 4'h3fb7;
         4'h9573 	:	val_out <= 4'h3fb7;
         4'h9578 	:	val_out <= 4'h3fa1;
         4'h9579 	:	val_out <= 4'h3fa1;
         4'h957a 	:	val_out <= 4'h3fa1;
         4'h957b 	:	val_out <= 4'h3fa1;
         4'h9580 	:	val_out <= 4'h3f8c;
         4'h9581 	:	val_out <= 4'h3f8c;
         4'h9582 	:	val_out <= 4'h3f8c;
         4'h9583 	:	val_out <= 4'h3f8c;
         4'h9588 	:	val_out <= 4'h3f76;
         4'h9589 	:	val_out <= 4'h3f76;
         4'h958a 	:	val_out <= 4'h3f76;
         4'h958b 	:	val_out <= 4'h3f76;
         4'h9590 	:	val_out <= 4'h3f60;
         4'h9591 	:	val_out <= 4'h3f60;
         4'h9592 	:	val_out <= 4'h3f60;
         4'h9593 	:	val_out <= 4'h3f60;
         4'h9598 	:	val_out <= 4'h3f4a;
         4'h9599 	:	val_out <= 4'h3f4a;
         4'h959a 	:	val_out <= 4'h3f4a;
         4'h959b 	:	val_out <= 4'h3f4a;
         4'h95a0 	:	val_out <= 4'h3f35;
         4'h95a1 	:	val_out <= 4'h3f35;
         4'h95a2 	:	val_out <= 4'h3f35;
         4'h95a3 	:	val_out <= 4'h3f35;
         4'h95a8 	:	val_out <= 4'h3f1f;
         4'h95a9 	:	val_out <= 4'h3f1f;
         4'h95aa 	:	val_out <= 4'h3f1f;
         4'h95ab 	:	val_out <= 4'h3f1f;
         4'h95b0 	:	val_out <= 4'h3f09;
         4'h95b1 	:	val_out <= 4'h3f09;
         4'h95b2 	:	val_out <= 4'h3f09;
         4'h95b3 	:	val_out <= 4'h3f09;
         4'h95b8 	:	val_out <= 4'h3ef4;
         4'h95b9 	:	val_out <= 4'h3ef4;
         4'h95ba 	:	val_out <= 4'h3ef4;
         4'h95bb 	:	val_out <= 4'h3ef4;
         4'h95c0 	:	val_out <= 4'h3ede;
         4'h95c1 	:	val_out <= 4'h3ede;
         4'h95c2 	:	val_out <= 4'h3ede;
         4'h95c3 	:	val_out <= 4'h3ede;
         4'h95c8 	:	val_out <= 4'h3ec9;
         4'h95c9 	:	val_out <= 4'h3ec9;
         4'h95ca 	:	val_out <= 4'h3ec9;
         4'h95cb 	:	val_out <= 4'h3ec9;
         4'h95d0 	:	val_out <= 4'h3eb3;
         4'h95d1 	:	val_out <= 4'h3eb3;
         4'h95d2 	:	val_out <= 4'h3eb3;
         4'h95d3 	:	val_out <= 4'h3eb3;
         4'h95d8 	:	val_out <= 4'h3e9d;
         4'h95d9 	:	val_out <= 4'h3e9d;
         4'h95da 	:	val_out <= 4'h3e9d;
         4'h95db 	:	val_out <= 4'h3e9d;
         4'h95e0 	:	val_out <= 4'h3e88;
         4'h95e1 	:	val_out <= 4'h3e88;
         4'h95e2 	:	val_out <= 4'h3e88;
         4'h95e3 	:	val_out <= 4'h3e88;
         4'h95e8 	:	val_out <= 4'h3e72;
         4'h95e9 	:	val_out <= 4'h3e72;
         4'h95ea 	:	val_out <= 4'h3e72;
         4'h95eb 	:	val_out <= 4'h3e72;
         4'h95f0 	:	val_out <= 4'h3e5d;
         4'h95f1 	:	val_out <= 4'h3e5d;
         4'h95f2 	:	val_out <= 4'h3e5d;
         4'h95f3 	:	val_out <= 4'h3e5d;
         4'h95f8 	:	val_out <= 4'h3e47;
         4'h95f9 	:	val_out <= 4'h3e47;
         4'h95fa 	:	val_out <= 4'h3e47;
         4'h95fb 	:	val_out <= 4'h3e47;
         4'h9600 	:	val_out <= 4'h3e31;
         4'h9601 	:	val_out <= 4'h3e31;
         4'h9602 	:	val_out <= 4'h3e31;
         4'h9603 	:	val_out <= 4'h3e31;
         4'h9608 	:	val_out <= 4'h3e1c;
         4'h9609 	:	val_out <= 4'h3e1c;
         4'h960a 	:	val_out <= 4'h3e1c;
         4'h960b 	:	val_out <= 4'h3e1c;
         4'h9610 	:	val_out <= 4'h3e06;
         4'h9611 	:	val_out <= 4'h3e06;
         4'h9612 	:	val_out <= 4'h3e06;
         4'h9613 	:	val_out <= 4'h3e06;
         4'h9618 	:	val_out <= 4'h3df1;
         4'h9619 	:	val_out <= 4'h3df1;
         4'h961a 	:	val_out <= 4'h3df1;
         4'h961b 	:	val_out <= 4'h3df1;
         4'h9620 	:	val_out <= 4'h3ddb;
         4'h9621 	:	val_out <= 4'h3ddb;
         4'h9622 	:	val_out <= 4'h3ddb;
         4'h9623 	:	val_out <= 4'h3ddb;
         4'h9628 	:	val_out <= 4'h3dc6;
         4'h9629 	:	val_out <= 4'h3dc6;
         4'h962a 	:	val_out <= 4'h3dc6;
         4'h962b 	:	val_out <= 4'h3dc6;
         4'h9630 	:	val_out <= 4'h3db0;
         4'h9631 	:	val_out <= 4'h3db0;
         4'h9632 	:	val_out <= 4'h3db0;
         4'h9633 	:	val_out <= 4'h3db0;
         4'h9638 	:	val_out <= 4'h3d9b;
         4'h9639 	:	val_out <= 4'h3d9b;
         4'h963a 	:	val_out <= 4'h3d9b;
         4'h963b 	:	val_out <= 4'h3d9b;
         4'h9640 	:	val_out <= 4'h3d85;
         4'h9641 	:	val_out <= 4'h3d85;
         4'h9642 	:	val_out <= 4'h3d85;
         4'h9643 	:	val_out <= 4'h3d85;
         4'h9648 	:	val_out <= 4'h3d70;
         4'h9649 	:	val_out <= 4'h3d70;
         4'h964a 	:	val_out <= 4'h3d70;
         4'h964b 	:	val_out <= 4'h3d70;
         4'h9650 	:	val_out <= 4'h3d5a;
         4'h9651 	:	val_out <= 4'h3d5a;
         4'h9652 	:	val_out <= 4'h3d5a;
         4'h9653 	:	val_out <= 4'h3d5a;
         4'h9658 	:	val_out <= 4'h3d45;
         4'h9659 	:	val_out <= 4'h3d45;
         4'h965a 	:	val_out <= 4'h3d45;
         4'h965b 	:	val_out <= 4'h3d45;
         4'h9660 	:	val_out <= 4'h3d2f;
         4'h9661 	:	val_out <= 4'h3d2f;
         4'h9662 	:	val_out <= 4'h3d2f;
         4'h9663 	:	val_out <= 4'h3d2f;
         4'h9668 	:	val_out <= 4'h3d1a;
         4'h9669 	:	val_out <= 4'h3d1a;
         4'h966a 	:	val_out <= 4'h3d1a;
         4'h966b 	:	val_out <= 4'h3d1a;
         4'h9670 	:	val_out <= 4'h3d05;
         4'h9671 	:	val_out <= 4'h3d05;
         4'h9672 	:	val_out <= 4'h3d05;
         4'h9673 	:	val_out <= 4'h3d05;
         4'h9678 	:	val_out <= 4'h3cef;
         4'h9679 	:	val_out <= 4'h3cef;
         4'h967a 	:	val_out <= 4'h3cef;
         4'h967b 	:	val_out <= 4'h3cef;
         4'h9680 	:	val_out <= 4'h3cda;
         4'h9681 	:	val_out <= 4'h3cda;
         4'h9682 	:	val_out <= 4'h3cda;
         4'h9683 	:	val_out <= 4'h3cda;
         4'h9688 	:	val_out <= 4'h3cc4;
         4'h9689 	:	val_out <= 4'h3cc4;
         4'h968a 	:	val_out <= 4'h3cc4;
         4'h968b 	:	val_out <= 4'h3cc4;
         4'h9690 	:	val_out <= 4'h3caf;
         4'h9691 	:	val_out <= 4'h3caf;
         4'h9692 	:	val_out <= 4'h3caf;
         4'h9693 	:	val_out <= 4'h3caf;
         4'h9698 	:	val_out <= 4'h3c9a;
         4'h9699 	:	val_out <= 4'h3c9a;
         4'h969a 	:	val_out <= 4'h3c9a;
         4'h969b 	:	val_out <= 4'h3c9a;
         4'h96a0 	:	val_out <= 4'h3c84;
         4'h96a1 	:	val_out <= 4'h3c84;
         4'h96a2 	:	val_out <= 4'h3c84;
         4'h96a3 	:	val_out <= 4'h3c84;
         4'h96a8 	:	val_out <= 4'h3c6f;
         4'h96a9 	:	val_out <= 4'h3c6f;
         4'h96aa 	:	val_out <= 4'h3c6f;
         4'h96ab 	:	val_out <= 4'h3c6f;
         4'h96b0 	:	val_out <= 4'h3c5a;
         4'h96b1 	:	val_out <= 4'h3c5a;
         4'h96b2 	:	val_out <= 4'h3c5a;
         4'h96b3 	:	val_out <= 4'h3c5a;
         4'h96b8 	:	val_out <= 4'h3c44;
         4'h96b9 	:	val_out <= 4'h3c44;
         4'h96ba 	:	val_out <= 4'h3c44;
         4'h96bb 	:	val_out <= 4'h3c44;
         4'h96c0 	:	val_out <= 4'h3c2f;
         4'h96c1 	:	val_out <= 4'h3c2f;
         4'h96c2 	:	val_out <= 4'h3c2f;
         4'h96c3 	:	val_out <= 4'h3c2f;
         4'h96c8 	:	val_out <= 4'h3c1a;
         4'h96c9 	:	val_out <= 4'h3c1a;
         4'h96ca 	:	val_out <= 4'h3c1a;
         4'h96cb 	:	val_out <= 4'h3c1a;
         4'h96d0 	:	val_out <= 4'h3c04;
         4'h96d1 	:	val_out <= 4'h3c04;
         4'h96d2 	:	val_out <= 4'h3c04;
         4'h96d3 	:	val_out <= 4'h3c04;
         4'h96d8 	:	val_out <= 4'h3bef;
         4'h96d9 	:	val_out <= 4'h3bef;
         4'h96da 	:	val_out <= 4'h3bef;
         4'h96db 	:	val_out <= 4'h3bef;
         4'h96e0 	:	val_out <= 4'h3bda;
         4'h96e1 	:	val_out <= 4'h3bda;
         4'h96e2 	:	val_out <= 4'h3bda;
         4'h96e3 	:	val_out <= 4'h3bda;
         4'h96e8 	:	val_out <= 4'h3bc4;
         4'h96e9 	:	val_out <= 4'h3bc4;
         4'h96ea 	:	val_out <= 4'h3bc4;
         4'h96eb 	:	val_out <= 4'h3bc4;
         4'h96f0 	:	val_out <= 4'h3baf;
         4'h96f1 	:	val_out <= 4'h3baf;
         4'h96f2 	:	val_out <= 4'h3baf;
         4'h96f3 	:	val_out <= 4'h3baf;
         4'h96f8 	:	val_out <= 4'h3b9a;
         4'h96f9 	:	val_out <= 4'h3b9a;
         4'h96fa 	:	val_out <= 4'h3b9a;
         4'h96fb 	:	val_out <= 4'h3b9a;
         4'h9700 	:	val_out <= 4'h3b85;
         4'h9701 	:	val_out <= 4'h3b85;
         4'h9702 	:	val_out <= 4'h3b85;
         4'h9703 	:	val_out <= 4'h3b85;
         4'h9708 	:	val_out <= 4'h3b6f;
         4'h9709 	:	val_out <= 4'h3b6f;
         4'h970a 	:	val_out <= 4'h3b6f;
         4'h970b 	:	val_out <= 4'h3b6f;
         4'h9710 	:	val_out <= 4'h3b5a;
         4'h9711 	:	val_out <= 4'h3b5a;
         4'h9712 	:	val_out <= 4'h3b5a;
         4'h9713 	:	val_out <= 4'h3b5a;
         4'h9718 	:	val_out <= 4'h3b45;
         4'h9719 	:	val_out <= 4'h3b45;
         4'h971a 	:	val_out <= 4'h3b45;
         4'h971b 	:	val_out <= 4'h3b45;
         4'h9720 	:	val_out <= 4'h3b30;
         4'h9721 	:	val_out <= 4'h3b30;
         4'h9722 	:	val_out <= 4'h3b30;
         4'h9723 	:	val_out <= 4'h3b30;
         4'h9728 	:	val_out <= 4'h3b1b;
         4'h9729 	:	val_out <= 4'h3b1b;
         4'h972a 	:	val_out <= 4'h3b1b;
         4'h972b 	:	val_out <= 4'h3b1b;
         4'h9730 	:	val_out <= 4'h3b05;
         4'h9731 	:	val_out <= 4'h3b05;
         4'h9732 	:	val_out <= 4'h3b05;
         4'h9733 	:	val_out <= 4'h3b05;
         4'h9738 	:	val_out <= 4'h3af0;
         4'h9739 	:	val_out <= 4'h3af0;
         4'h973a 	:	val_out <= 4'h3af0;
         4'h973b 	:	val_out <= 4'h3af0;
         4'h9740 	:	val_out <= 4'h3adb;
         4'h9741 	:	val_out <= 4'h3adb;
         4'h9742 	:	val_out <= 4'h3adb;
         4'h9743 	:	val_out <= 4'h3adb;
         4'h9748 	:	val_out <= 4'h3ac6;
         4'h9749 	:	val_out <= 4'h3ac6;
         4'h974a 	:	val_out <= 4'h3ac6;
         4'h974b 	:	val_out <= 4'h3ac6;
         4'h9750 	:	val_out <= 4'h3ab1;
         4'h9751 	:	val_out <= 4'h3ab1;
         4'h9752 	:	val_out <= 4'h3ab1;
         4'h9753 	:	val_out <= 4'h3ab1;
         4'h9758 	:	val_out <= 4'h3a9c;
         4'h9759 	:	val_out <= 4'h3a9c;
         4'h975a 	:	val_out <= 4'h3a9c;
         4'h975b 	:	val_out <= 4'h3a9c;
         4'h9760 	:	val_out <= 4'h3a87;
         4'h9761 	:	val_out <= 4'h3a87;
         4'h9762 	:	val_out <= 4'h3a87;
         4'h9763 	:	val_out <= 4'h3a87;
         4'h9768 	:	val_out <= 4'h3a72;
         4'h9769 	:	val_out <= 4'h3a72;
         4'h976a 	:	val_out <= 4'h3a72;
         4'h976b 	:	val_out <= 4'h3a72;
         4'h9770 	:	val_out <= 4'h3a5c;
         4'h9771 	:	val_out <= 4'h3a5c;
         4'h9772 	:	val_out <= 4'h3a5c;
         4'h9773 	:	val_out <= 4'h3a5c;
         4'h9778 	:	val_out <= 4'h3a47;
         4'h9779 	:	val_out <= 4'h3a47;
         4'h977a 	:	val_out <= 4'h3a47;
         4'h977b 	:	val_out <= 4'h3a47;
         4'h9780 	:	val_out <= 4'h3a32;
         4'h9781 	:	val_out <= 4'h3a32;
         4'h9782 	:	val_out <= 4'h3a32;
         4'h9783 	:	val_out <= 4'h3a32;
         4'h9788 	:	val_out <= 4'h3a1d;
         4'h9789 	:	val_out <= 4'h3a1d;
         4'h978a 	:	val_out <= 4'h3a1d;
         4'h978b 	:	val_out <= 4'h3a1d;
         4'h9790 	:	val_out <= 4'h3a08;
         4'h9791 	:	val_out <= 4'h3a08;
         4'h9792 	:	val_out <= 4'h3a08;
         4'h9793 	:	val_out <= 4'h3a08;
         4'h9798 	:	val_out <= 4'h39f3;
         4'h9799 	:	val_out <= 4'h39f3;
         4'h979a 	:	val_out <= 4'h39f3;
         4'h979b 	:	val_out <= 4'h39f3;
         4'h97a0 	:	val_out <= 4'h39de;
         4'h97a1 	:	val_out <= 4'h39de;
         4'h97a2 	:	val_out <= 4'h39de;
         4'h97a3 	:	val_out <= 4'h39de;
         4'h97a8 	:	val_out <= 4'h39c9;
         4'h97a9 	:	val_out <= 4'h39c9;
         4'h97aa 	:	val_out <= 4'h39c9;
         4'h97ab 	:	val_out <= 4'h39c9;
         4'h97b0 	:	val_out <= 4'h39b4;
         4'h97b1 	:	val_out <= 4'h39b4;
         4'h97b2 	:	val_out <= 4'h39b4;
         4'h97b3 	:	val_out <= 4'h39b4;
         4'h97b8 	:	val_out <= 4'h399f;
         4'h97b9 	:	val_out <= 4'h399f;
         4'h97ba 	:	val_out <= 4'h399f;
         4'h97bb 	:	val_out <= 4'h399f;
         4'h97c0 	:	val_out <= 4'h398a;
         4'h97c1 	:	val_out <= 4'h398a;
         4'h97c2 	:	val_out <= 4'h398a;
         4'h97c3 	:	val_out <= 4'h398a;
         4'h97c8 	:	val_out <= 4'h3975;
         4'h97c9 	:	val_out <= 4'h3975;
         4'h97ca 	:	val_out <= 4'h3975;
         4'h97cb 	:	val_out <= 4'h3975;
         4'h97d0 	:	val_out <= 4'h3960;
         4'h97d1 	:	val_out <= 4'h3960;
         4'h97d2 	:	val_out <= 4'h3960;
         4'h97d3 	:	val_out <= 4'h3960;
         4'h97d8 	:	val_out <= 4'h394b;
         4'h97d9 	:	val_out <= 4'h394b;
         4'h97da 	:	val_out <= 4'h394b;
         4'h97db 	:	val_out <= 4'h394b;
         4'h97e0 	:	val_out <= 4'h3936;
         4'h97e1 	:	val_out <= 4'h3936;
         4'h97e2 	:	val_out <= 4'h3936;
         4'h97e3 	:	val_out <= 4'h3936;
         4'h97e8 	:	val_out <= 4'h3921;
         4'h97e9 	:	val_out <= 4'h3921;
         4'h97ea 	:	val_out <= 4'h3921;
         4'h97eb 	:	val_out <= 4'h3921;
         4'h97f0 	:	val_out <= 4'h390c;
         4'h97f1 	:	val_out <= 4'h390c;
         4'h97f2 	:	val_out <= 4'h390c;
         4'h97f3 	:	val_out <= 4'h390c;
         4'h97f8 	:	val_out <= 4'h38f7;
         4'h97f9 	:	val_out <= 4'h38f7;
         4'h97fa 	:	val_out <= 4'h38f7;
         4'h97fb 	:	val_out <= 4'h38f7;
         4'h9800 	:	val_out <= 4'h38e3;
         4'h9801 	:	val_out <= 4'h38e3;
         4'h9802 	:	val_out <= 4'h38e3;
         4'h9803 	:	val_out <= 4'h38e3;
         4'h9808 	:	val_out <= 4'h38ce;
         4'h9809 	:	val_out <= 4'h38ce;
         4'h980a 	:	val_out <= 4'h38ce;
         4'h980b 	:	val_out <= 4'h38ce;
         4'h9810 	:	val_out <= 4'h38b9;
         4'h9811 	:	val_out <= 4'h38b9;
         4'h9812 	:	val_out <= 4'h38b9;
         4'h9813 	:	val_out <= 4'h38b9;
         4'h9818 	:	val_out <= 4'h38a4;
         4'h9819 	:	val_out <= 4'h38a4;
         4'h981a 	:	val_out <= 4'h38a4;
         4'h981b 	:	val_out <= 4'h38a4;
         4'h9820 	:	val_out <= 4'h388f;
         4'h9821 	:	val_out <= 4'h388f;
         4'h9822 	:	val_out <= 4'h388f;
         4'h9823 	:	val_out <= 4'h388f;
         4'h9828 	:	val_out <= 4'h387a;
         4'h9829 	:	val_out <= 4'h387a;
         4'h982a 	:	val_out <= 4'h387a;
         4'h982b 	:	val_out <= 4'h387a;
         4'h9830 	:	val_out <= 4'h3865;
         4'h9831 	:	val_out <= 4'h3865;
         4'h9832 	:	val_out <= 4'h3865;
         4'h9833 	:	val_out <= 4'h3865;
         4'h9838 	:	val_out <= 4'h3851;
         4'h9839 	:	val_out <= 4'h3851;
         4'h983a 	:	val_out <= 4'h3851;
         4'h983b 	:	val_out <= 4'h3851;
         4'h9840 	:	val_out <= 4'h383c;
         4'h9841 	:	val_out <= 4'h383c;
         4'h9842 	:	val_out <= 4'h383c;
         4'h9843 	:	val_out <= 4'h383c;
         4'h9848 	:	val_out <= 4'h3827;
         4'h9849 	:	val_out <= 4'h3827;
         4'h984a 	:	val_out <= 4'h3827;
         4'h984b 	:	val_out <= 4'h3827;
         4'h9850 	:	val_out <= 4'h3812;
         4'h9851 	:	val_out <= 4'h3812;
         4'h9852 	:	val_out <= 4'h3812;
         4'h9853 	:	val_out <= 4'h3812;
         4'h9858 	:	val_out <= 4'h37fd;
         4'h9859 	:	val_out <= 4'h37fd;
         4'h985a 	:	val_out <= 4'h37fd;
         4'h985b 	:	val_out <= 4'h37fd;
         4'h9860 	:	val_out <= 4'h37e9;
         4'h9861 	:	val_out <= 4'h37e9;
         4'h9862 	:	val_out <= 4'h37e9;
         4'h9863 	:	val_out <= 4'h37e9;
         4'h9868 	:	val_out <= 4'h37d4;
         4'h9869 	:	val_out <= 4'h37d4;
         4'h986a 	:	val_out <= 4'h37d4;
         4'h986b 	:	val_out <= 4'h37d4;
         4'h9870 	:	val_out <= 4'h37bf;
         4'h9871 	:	val_out <= 4'h37bf;
         4'h9872 	:	val_out <= 4'h37bf;
         4'h9873 	:	val_out <= 4'h37bf;
         4'h9878 	:	val_out <= 4'h37aa;
         4'h9879 	:	val_out <= 4'h37aa;
         4'h987a 	:	val_out <= 4'h37aa;
         4'h987b 	:	val_out <= 4'h37aa;
         4'h9880 	:	val_out <= 4'h3796;
         4'h9881 	:	val_out <= 4'h3796;
         4'h9882 	:	val_out <= 4'h3796;
         4'h9883 	:	val_out <= 4'h3796;
         4'h9888 	:	val_out <= 4'h3781;
         4'h9889 	:	val_out <= 4'h3781;
         4'h988a 	:	val_out <= 4'h3781;
         4'h988b 	:	val_out <= 4'h3781;
         4'h9890 	:	val_out <= 4'h376c;
         4'h9891 	:	val_out <= 4'h376c;
         4'h9892 	:	val_out <= 4'h376c;
         4'h9893 	:	val_out <= 4'h376c;
         4'h9898 	:	val_out <= 4'h3757;
         4'h9899 	:	val_out <= 4'h3757;
         4'h989a 	:	val_out <= 4'h3757;
         4'h989b 	:	val_out <= 4'h3757;
         4'h98a0 	:	val_out <= 4'h3743;
         4'h98a1 	:	val_out <= 4'h3743;
         4'h98a2 	:	val_out <= 4'h3743;
         4'h98a3 	:	val_out <= 4'h3743;
         4'h98a8 	:	val_out <= 4'h372e;
         4'h98a9 	:	val_out <= 4'h372e;
         4'h98aa 	:	val_out <= 4'h372e;
         4'h98ab 	:	val_out <= 4'h372e;
         4'h98b0 	:	val_out <= 4'h3719;
         4'h98b1 	:	val_out <= 4'h3719;
         4'h98b2 	:	val_out <= 4'h3719;
         4'h98b3 	:	val_out <= 4'h3719;
         4'h98b8 	:	val_out <= 4'h3705;
         4'h98b9 	:	val_out <= 4'h3705;
         4'h98ba 	:	val_out <= 4'h3705;
         4'h98bb 	:	val_out <= 4'h3705;
         4'h98c0 	:	val_out <= 4'h36f0;
         4'h98c1 	:	val_out <= 4'h36f0;
         4'h98c2 	:	val_out <= 4'h36f0;
         4'h98c3 	:	val_out <= 4'h36f0;
         4'h98c8 	:	val_out <= 4'h36dc;
         4'h98c9 	:	val_out <= 4'h36dc;
         4'h98ca 	:	val_out <= 4'h36dc;
         4'h98cb 	:	val_out <= 4'h36dc;
         4'h98d0 	:	val_out <= 4'h36c7;
         4'h98d1 	:	val_out <= 4'h36c7;
         4'h98d2 	:	val_out <= 4'h36c7;
         4'h98d3 	:	val_out <= 4'h36c7;
         4'h98d8 	:	val_out <= 4'h36b2;
         4'h98d9 	:	val_out <= 4'h36b2;
         4'h98da 	:	val_out <= 4'h36b2;
         4'h98db 	:	val_out <= 4'h36b2;
         4'h98e0 	:	val_out <= 4'h369e;
         4'h98e1 	:	val_out <= 4'h369e;
         4'h98e2 	:	val_out <= 4'h369e;
         4'h98e3 	:	val_out <= 4'h369e;
         4'h98e8 	:	val_out <= 4'h3689;
         4'h98e9 	:	val_out <= 4'h3689;
         4'h98ea 	:	val_out <= 4'h3689;
         4'h98eb 	:	val_out <= 4'h3689;
         4'h98f0 	:	val_out <= 4'h3675;
         4'h98f1 	:	val_out <= 4'h3675;
         4'h98f2 	:	val_out <= 4'h3675;
         4'h98f3 	:	val_out <= 4'h3675;
         4'h98f8 	:	val_out <= 4'h3660;
         4'h98f9 	:	val_out <= 4'h3660;
         4'h98fa 	:	val_out <= 4'h3660;
         4'h98fb 	:	val_out <= 4'h3660;
         4'h9900 	:	val_out <= 4'h364b;
         4'h9901 	:	val_out <= 4'h364b;
         4'h9902 	:	val_out <= 4'h364b;
         4'h9903 	:	val_out <= 4'h364b;
         4'h9908 	:	val_out <= 4'h3637;
         4'h9909 	:	val_out <= 4'h3637;
         4'h990a 	:	val_out <= 4'h3637;
         4'h990b 	:	val_out <= 4'h3637;
         4'h9910 	:	val_out <= 4'h3622;
         4'h9911 	:	val_out <= 4'h3622;
         4'h9912 	:	val_out <= 4'h3622;
         4'h9913 	:	val_out <= 4'h3622;
         4'h9918 	:	val_out <= 4'h360e;
         4'h9919 	:	val_out <= 4'h360e;
         4'h991a 	:	val_out <= 4'h360e;
         4'h991b 	:	val_out <= 4'h360e;
         4'h9920 	:	val_out <= 4'h35f9;
         4'h9921 	:	val_out <= 4'h35f9;
         4'h9922 	:	val_out <= 4'h35f9;
         4'h9923 	:	val_out <= 4'h35f9;
         4'h9928 	:	val_out <= 4'h35e5;
         4'h9929 	:	val_out <= 4'h35e5;
         4'h992a 	:	val_out <= 4'h35e5;
         4'h992b 	:	val_out <= 4'h35e5;
         4'h9930 	:	val_out <= 4'h35d0;
         4'h9931 	:	val_out <= 4'h35d0;
         4'h9932 	:	val_out <= 4'h35d0;
         4'h9933 	:	val_out <= 4'h35d0;
         4'h9938 	:	val_out <= 4'h35bc;
         4'h9939 	:	val_out <= 4'h35bc;
         4'h993a 	:	val_out <= 4'h35bc;
         4'h993b 	:	val_out <= 4'h35bc;
         4'h9940 	:	val_out <= 4'h35a7;
         4'h9941 	:	val_out <= 4'h35a7;
         4'h9942 	:	val_out <= 4'h35a7;
         4'h9943 	:	val_out <= 4'h35a7;
         4'h9948 	:	val_out <= 4'h3593;
         4'h9949 	:	val_out <= 4'h3593;
         4'h994a 	:	val_out <= 4'h3593;
         4'h994b 	:	val_out <= 4'h3593;
         4'h9950 	:	val_out <= 4'h357e;
         4'h9951 	:	val_out <= 4'h357e;
         4'h9952 	:	val_out <= 4'h357e;
         4'h9953 	:	val_out <= 4'h357e;
         4'h9958 	:	val_out <= 4'h356a;
         4'h9959 	:	val_out <= 4'h356a;
         4'h995a 	:	val_out <= 4'h356a;
         4'h995b 	:	val_out <= 4'h356a;
         4'h9960 	:	val_out <= 4'h3556;
         4'h9961 	:	val_out <= 4'h3556;
         4'h9962 	:	val_out <= 4'h3556;
         4'h9963 	:	val_out <= 4'h3556;
         4'h9968 	:	val_out <= 4'h3541;
         4'h9969 	:	val_out <= 4'h3541;
         4'h996a 	:	val_out <= 4'h3541;
         4'h996b 	:	val_out <= 4'h3541;
         4'h9970 	:	val_out <= 4'h352d;
         4'h9971 	:	val_out <= 4'h352d;
         4'h9972 	:	val_out <= 4'h352d;
         4'h9973 	:	val_out <= 4'h352d;
         4'h9978 	:	val_out <= 4'h3518;
         4'h9979 	:	val_out <= 4'h3518;
         4'h997a 	:	val_out <= 4'h3518;
         4'h997b 	:	val_out <= 4'h3518;
         4'h9980 	:	val_out <= 4'h3504;
         4'h9981 	:	val_out <= 4'h3504;
         4'h9982 	:	val_out <= 4'h3504;
         4'h9983 	:	val_out <= 4'h3504;
         4'h9988 	:	val_out <= 4'h34f0;
         4'h9989 	:	val_out <= 4'h34f0;
         4'h998a 	:	val_out <= 4'h34f0;
         4'h998b 	:	val_out <= 4'h34f0;
         4'h9990 	:	val_out <= 4'h34db;
         4'h9991 	:	val_out <= 4'h34db;
         4'h9992 	:	val_out <= 4'h34db;
         4'h9993 	:	val_out <= 4'h34db;
         4'h9998 	:	val_out <= 4'h34c7;
         4'h9999 	:	val_out <= 4'h34c7;
         4'h999a 	:	val_out <= 4'h34c7;
         4'h999b 	:	val_out <= 4'h34c7;
         4'h99a0 	:	val_out <= 4'h34b3;
         4'h99a1 	:	val_out <= 4'h34b3;
         4'h99a2 	:	val_out <= 4'h34b3;
         4'h99a3 	:	val_out <= 4'h34b3;
         4'h99a8 	:	val_out <= 4'h349e;
         4'h99a9 	:	val_out <= 4'h349e;
         4'h99aa 	:	val_out <= 4'h349e;
         4'h99ab 	:	val_out <= 4'h349e;
         4'h99b0 	:	val_out <= 4'h348a;
         4'h99b1 	:	val_out <= 4'h348a;
         4'h99b2 	:	val_out <= 4'h348a;
         4'h99b3 	:	val_out <= 4'h348a;
         4'h99b8 	:	val_out <= 4'h3476;
         4'h99b9 	:	val_out <= 4'h3476;
         4'h99ba 	:	val_out <= 4'h3476;
         4'h99bb 	:	val_out <= 4'h3476;
         4'h99c0 	:	val_out <= 4'h3461;
         4'h99c1 	:	val_out <= 4'h3461;
         4'h99c2 	:	val_out <= 4'h3461;
         4'h99c3 	:	val_out <= 4'h3461;
         4'h99c8 	:	val_out <= 4'h344d;
         4'h99c9 	:	val_out <= 4'h344d;
         4'h99ca 	:	val_out <= 4'h344d;
         4'h99cb 	:	val_out <= 4'h344d;
         4'h99d0 	:	val_out <= 4'h3439;
         4'h99d1 	:	val_out <= 4'h3439;
         4'h99d2 	:	val_out <= 4'h3439;
         4'h99d3 	:	val_out <= 4'h3439;
         4'h99d8 	:	val_out <= 4'h3425;
         4'h99d9 	:	val_out <= 4'h3425;
         4'h99da 	:	val_out <= 4'h3425;
         4'h99db 	:	val_out <= 4'h3425;
         4'h99e0 	:	val_out <= 4'h3410;
         4'h99e1 	:	val_out <= 4'h3410;
         4'h99e2 	:	val_out <= 4'h3410;
         4'h99e3 	:	val_out <= 4'h3410;
         4'h99e8 	:	val_out <= 4'h33fc;
         4'h99e9 	:	val_out <= 4'h33fc;
         4'h99ea 	:	val_out <= 4'h33fc;
         4'h99eb 	:	val_out <= 4'h33fc;
         4'h99f0 	:	val_out <= 4'h33e8;
         4'h99f1 	:	val_out <= 4'h33e8;
         4'h99f2 	:	val_out <= 4'h33e8;
         4'h99f3 	:	val_out <= 4'h33e8;
         4'h99f8 	:	val_out <= 4'h33d4;
         4'h99f9 	:	val_out <= 4'h33d4;
         4'h99fa 	:	val_out <= 4'h33d4;
         4'h99fb 	:	val_out <= 4'h33d4;
         4'h9a00 	:	val_out <= 4'h33c0;
         4'h9a01 	:	val_out <= 4'h33c0;
         4'h9a02 	:	val_out <= 4'h33c0;
         4'h9a03 	:	val_out <= 4'h33c0;
         4'h9a08 	:	val_out <= 4'h33ab;
         4'h9a09 	:	val_out <= 4'h33ab;
         4'h9a0a 	:	val_out <= 4'h33ab;
         4'h9a0b 	:	val_out <= 4'h33ab;
         4'h9a10 	:	val_out <= 4'h3397;
         4'h9a11 	:	val_out <= 4'h3397;
         4'h9a12 	:	val_out <= 4'h3397;
         4'h9a13 	:	val_out <= 4'h3397;
         4'h9a18 	:	val_out <= 4'h3383;
         4'h9a19 	:	val_out <= 4'h3383;
         4'h9a1a 	:	val_out <= 4'h3383;
         4'h9a1b 	:	val_out <= 4'h3383;
         4'h9a20 	:	val_out <= 4'h336f;
         4'h9a21 	:	val_out <= 4'h336f;
         4'h9a22 	:	val_out <= 4'h336f;
         4'h9a23 	:	val_out <= 4'h336f;
         4'h9a28 	:	val_out <= 4'h335b;
         4'h9a29 	:	val_out <= 4'h335b;
         4'h9a2a 	:	val_out <= 4'h335b;
         4'h9a2b 	:	val_out <= 4'h335b;
         4'h9a30 	:	val_out <= 4'h3347;
         4'h9a31 	:	val_out <= 4'h3347;
         4'h9a32 	:	val_out <= 4'h3347;
         4'h9a33 	:	val_out <= 4'h3347;
         4'h9a38 	:	val_out <= 4'h3333;
         4'h9a39 	:	val_out <= 4'h3333;
         4'h9a3a 	:	val_out <= 4'h3333;
         4'h9a3b 	:	val_out <= 4'h3333;
         4'h9a40 	:	val_out <= 4'h331e;
         4'h9a41 	:	val_out <= 4'h331e;
         4'h9a42 	:	val_out <= 4'h331e;
         4'h9a43 	:	val_out <= 4'h331e;
         4'h9a48 	:	val_out <= 4'h330a;
         4'h9a49 	:	val_out <= 4'h330a;
         4'h9a4a 	:	val_out <= 4'h330a;
         4'h9a4b 	:	val_out <= 4'h330a;
         4'h9a50 	:	val_out <= 4'h32f6;
         4'h9a51 	:	val_out <= 4'h32f6;
         4'h9a52 	:	val_out <= 4'h32f6;
         4'h9a53 	:	val_out <= 4'h32f6;
         4'h9a58 	:	val_out <= 4'h32e2;
         4'h9a59 	:	val_out <= 4'h32e2;
         4'h9a5a 	:	val_out <= 4'h32e2;
         4'h9a5b 	:	val_out <= 4'h32e2;
         4'h9a60 	:	val_out <= 4'h32ce;
         4'h9a61 	:	val_out <= 4'h32ce;
         4'h9a62 	:	val_out <= 4'h32ce;
         4'h9a63 	:	val_out <= 4'h32ce;
         4'h9a68 	:	val_out <= 4'h32ba;
         4'h9a69 	:	val_out <= 4'h32ba;
         4'h9a6a 	:	val_out <= 4'h32ba;
         4'h9a6b 	:	val_out <= 4'h32ba;
         4'h9a70 	:	val_out <= 4'h32a6;
         4'h9a71 	:	val_out <= 4'h32a6;
         4'h9a72 	:	val_out <= 4'h32a6;
         4'h9a73 	:	val_out <= 4'h32a6;
         4'h9a78 	:	val_out <= 4'h3292;
         4'h9a79 	:	val_out <= 4'h3292;
         4'h9a7a 	:	val_out <= 4'h3292;
         4'h9a7b 	:	val_out <= 4'h3292;
         4'h9a80 	:	val_out <= 4'h327e;
         4'h9a81 	:	val_out <= 4'h327e;
         4'h9a82 	:	val_out <= 4'h327e;
         4'h9a83 	:	val_out <= 4'h327e;
         4'h9a88 	:	val_out <= 4'h326a;
         4'h9a89 	:	val_out <= 4'h326a;
         4'h9a8a 	:	val_out <= 4'h326a;
         4'h9a8b 	:	val_out <= 4'h326a;
         4'h9a90 	:	val_out <= 4'h3256;
         4'h9a91 	:	val_out <= 4'h3256;
         4'h9a92 	:	val_out <= 4'h3256;
         4'h9a93 	:	val_out <= 4'h3256;
         4'h9a98 	:	val_out <= 4'h3242;
         4'h9a99 	:	val_out <= 4'h3242;
         4'h9a9a 	:	val_out <= 4'h3242;
         4'h9a9b 	:	val_out <= 4'h3242;
         4'h9aa0 	:	val_out <= 4'h322e;
         4'h9aa1 	:	val_out <= 4'h322e;
         4'h9aa2 	:	val_out <= 4'h322e;
         4'h9aa3 	:	val_out <= 4'h322e;
         4'h9aa8 	:	val_out <= 4'h321a;
         4'h9aa9 	:	val_out <= 4'h321a;
         4'h9aaa 	:	val_out <= 4'h321a;
         4'h9aab 	:	val_out <= 4'h321a;
         4'h9ab0 	:	val_out <= 4'h3206;
         4'h9ab1 	:	val_out <= 4'h3206;
         4'h9ab2 	:	val_out <= 4'h3206;
         4'h9ab3 	:	val_out <= 4'h3206;
         4'h9ab8 	:	val_out <= 4'h31f2;
         4'h9ab9 	:	val_out <= 4'h31f2;
         4'h9aba 	:	val_out <= 4'h31f2;
         4'h9abb 	:	val_out <= 4'h31f2;
         4'h9ac0 	:	val_out <= 4'h31de;
         4'h9ac1 	:	val_out <= 4'h31de;
         4'h9ac2 	:	val_out <= 4'h31de;
         4'h9ac3 	:	val_out <= 4'h31de;
         4'h9ac8 	:	val_out <= 4'h31cb;
         4'h9ac9 	:	val_out <= 4'h31cb;
         4'h9aca 	:	val_out <= 4'h31cb;
         4'h9acb 	:	val_out <= 4'h31cb;
         4'h9ad0 	:	val_out <= 4'h31b7;
         4'h9ad1 	:	val_out <= 4'h31b7;
         4'h9ad2 	:	val_out <= 4'h31b7;
         4'h9ad3 	:	val_out <= 4'h31b7;
         4'h9ad8 	:	val_out <= 4'h31a3;
         4'h9ad9 	:	val_out <= 4'h31a3;
         4'h9ada 	:	val_out <= 4'h31a3;
         4'h9adb 	:	val_out <= 4'h31a3;
         4'h9ae0 	:	val_out <= 4'h318f;
         4'h9ae1 	:	val_out <= 4'h318f;
         4'h9ae2 	:	val_out <= 4'h318f;
         4'h9ae3 	:	val_out <= 4'h318f;
         4'h9ae8 	:	val_out <= 4'h317b;
         4'h9ae9 	:	val_out <= 4'h317b;
         4'h9aea 	:	val_out <= 4'h317b;
         4'h9aeb 	:	val_out <= 4'h317b;
         4'h9af0 	:	val_out <= 4'h3167;
         4'h9af1 	:	val_out <= 4'h3167;
         4'h9af2 	:	val_out <= 4'h3167;
         4'h9af3 	:	val_out <= 4'h3167;
         4'h9af8 	:	val_out <= 4'h3153;
         4'h9af9 	:	val_out <= 4'h3153;
         4'h9afa 	:	val_out <= 4'h3153;
         4'h9afb 	:	val_out <= 4'h3153;
         4'h9b00 	:	val_out <= 4'h3140;
         4'h9b01 	:	val_out <= 4'h3140;
         4'h9b02 	:	val_out <= 4'h3140;
         4'h9b03 	:	val_out <= 4'h3140;
         4'h9b08 	:	val_out <= 4'h312c;
         4'h9b09 	:	val_out <= 4'h312c;
         4'h9b0a 	:	val_out <= 4'h312c;
         4'h9b0b 	:	val_out <= 4'h312c;
         4'h9b10 	:	val_out <= 4'h3118;
         4'h9b11 	:	val_out <= 4'h3118;
         4'h9b12 	:	val_out <= 4'h3118;
         4'h9b13 	:	val_out <= 4'h3118;
         4'h9b18 	:	val_out <= 4'h3104;
         4'h9b19 	:	val_out <= 4'h3104;
         4'h9b1a 	:	val_out <= 4'h3104;
         4'h9b1b 	:	val_out <= 4'h3104;
         4'h9b20 	:	val_out <= 4'h30f0;
         4'h9b21 	:	val_out <= 4'h30f0;
         4'h9b22 	:	val_out <= 4'h30f0;
         4'h9b23 	:	val_out <= 4'h30f0;
         4'h9b28 	:	val_out <= 4'h30dd;
         4'h9b29 	:	val_out <= 4'h30dd;
         4'h9b2a 	:	val_out <= 4'h30dd;
         4'h9b2b 	:	val_out <= 4'h30dd;
         4'h9b30 	:	val_out <= 4'h30c9;
         4'h9b31 	:	val_out <= 4'h30c9;
         4'h9b32 	:	val_out <= 4'h30c9;
         4'h9b33 	:	val_out <= 4'h30c9;
         4'h9b38 	:	val_out <= 4'h30b5;
         4'h9b39 	:	val_out <= 4'h30b5;
         4'h9b3a 	:	val_out <= 4'h30b5;
         4'h9b3b 	:	val_out <= 4'h30b5;
         4'h9b40 	:	val_out <= 4'h30a1;
         4'h9b41 	:	val_out <= 4'h30a1;
         4'h9b42 	:	val_out <= 4'h30a1;
         4'h9b43 	:	val_out <= 4'h30a1;
         4'h9b48 	:	val_out <= 4'h308e;
         4'h9b49 	:	val_out <= 4'h308e;
         4'h9b4a 	:	val_out <= 4'h308e;
         4'h9b4b 	:	val_out <= 4'h308e;
         4'h9b50 	:	val_out <= 4'h307a;
         4'h9b51 	:	val_out <= 4'h307a;
         4'h9b52 	:	val_out <= 4'h307a;
         4'h9b53 	:	val_out <= 4'h307a;
         4'h9b58 	:	val_out <= 4'h3066;
         4'h9b59 	:	val_out <= 4'h3066;
         4'h9b5a 	:	val_out <= 4'h3066;
         4'h9b5b 	:	val_out <= 4'h3066;
         4'h9b60 	:	val_out <= 4'h3053;
         4'h9b61 	:	val_out <= 4'h3053;
         4'h9b62 	:	val_out <= 4'h3053;
         4'h9b63 	:	val_out <= 4'h3053;
         4'h9b68 	:	val_out <= 4'h303f;
         4'h9b69 	:	val_out <= 4'h303f;
         4'h9b6a 	:	val_out <= 4'h303f;
         4'h9b6b 	:	val_out <= 4'h303f;
         4'h9b70 	:	val_out <= 4'h302b;
         4'h9b71 	:	val_out <= 4'h302b;
         4'h9b72 	:	val_out <= 4'h302b;
         4'h9b73 	:	val_out <= 4'h302b;
         4'h9b78 	:	val_out <= 4'h3018;
         4'h9b79 	:	val_out <= 4'h3018;
         4'h9b7a 	:	val_out <= 4'h3018;
         4'h9b7b 	:	val_out <= 4'h3018;
         4'h9b80 	:	val_out <= 4'h3004;
         4'h9b81 	:	val_out <= 4'h3004;
         4'h9b82 	:	val_out <= 4'h3004;
         4'h9b83 	:	val_out <= 4'h3004;
         4'h9b88 	:	val_out <= 4'h2ff0;
         4'h9b89 	:	val_out <= 4'h2ff0;
         4'h9b8a 	:	val_out <= 4'h2ff0;
         4'h9b8b 	:	val_out <= 4'h2ff0;
         4'h9b90 	:	val_out <= 4'h2fdd;
         4'h9b91 	:	val_out <= 4'h2fdd;
         4'h9b92 	:	val_out <= 4'h2fdd;
         4'h9b93 	:	val_out <= 4'h2fdd;
         4'h9b98 	:	val_out <= 4'h2fc9;
         4'h9b99 	:	val_out <= 4'h2fc9;
         4'h9b9a 	:	val_out <= 4'h2fc9;
         4'h9b9b 	:	val_out <= 4'h2fc9;
         4'h9ba0 	:	val_out <= 4'h2fb6;
         4'h9ba1 	:	val_out <= 4'h2fb6;
         4'h9ba2 	:	val_out <= 4'h2fb6;
         4'h9ba3 	:	val_out <= 4'h2fb6;
         4'h9ba8 	:	val_out <= 4'h2fa2;
         4'h9ba9 	:	val_out <= 4'h2fa2;
         4'h9baa 	:	val_out <= 4'h2fa2;
         4'h9bab 	:	val_out <= 4'h2fa2;
         4'h9bb0 	:	val_out <= 4'h2f8f;
         4'h9bb1 	:	val_out <= 4'h2f8f;
         4'h9bb2 	:	val_out <= 4'h2f8f;
         4'h9bb3 	:	val_out <= 4'h2f8f;
         4'h9bb8 	:	val_out <= 4'h2f7b;
         4'h9bb9 	:	val_out <= 4'h2f7b;
         4'h9bba 	:	val_out <= 4'h2f7b;
         4'h9bbb 	:	val_out <= 4'h2f7b;
         4'h9bc0 	:	val_out <= 4'h2f68;
         4'h9bc1 	:	val_out <= 4'h2f68;
         4'h9bc2 	:	val_out <= 4'h2f68;
         4'h9bc3 	:	val_out <= 4'h2f68;
         4'h9bc8 	:	val_out <= 4'h2f54;
         4'h9bc9 	:	val_out <= 4'h2f54;
         4'h9bca 	:	val_out <= 4'h2f54;
         4'h9bcb 	:	val_out <= 4'h2f54;
         4'h9bd0 	:	val_out <= 4'h2f40;
         4'h9bd1 	:	val_out <= 4'h2f40;
         4'h9bd2 	:	val_out <= 4'h2f40;
         4'h9bd3 	:	val_out <= 4'h2f40;
         4'h9bd8 	:	val_out <= 4'h2f2d;
         4'h9bd9 	:	val_out <= 4'h2f2d;
         4'h9bda 	:	val_out <= 4'h2f2d;
         4'h9bdb 	:	val_out <= 4'h2f2d;
         4'h9be0 	:	val_out <= 4'h2f1a;
         4'h9be1 	:	val_out <= 4'h2f1a;
         4'h9be2 	:	val_out <= 4'h2f1a;
         4'h9be3 	:	val_out <= 4'h2f1a;
         4'h9be8 	:	val_out <= 4'h2f06;
         4'h9be9 	:	val_out <= 4'h2f06;
         4'h9bea 	:	val_out <= 4'h2f06;
         4'h9beb 	:	val_out <= 4'h2f06;
         4'h9bf0 	:	val_out <= 4'h2ef3;
         4'h9bf1 	:	val_out <= 4'h2ef3;
         4'h9bf2 	:	val_out <= 4'h2ef3;
         4'h9bf3 	:	val_out <= 4'h2ef3;
         4'h9bf8 	:	val_out <= 4'h2edf;
         4'h9bf9 	:	val_out <= 4'h2edf;
         4'h9bfa 	:	val_out <= 4'h2edf;
         4'h9bfb 	:	val_out <= 4'h2edf;
         4'h9c00 	:	val_out <= 4'h2ecc;
         4'h9c01 	:	val_out <= 4'h2ecc;
         4'h9c02 	:	val_out <= 4'h2ecc;
         4'h9c03 	:	val_out <= 4'h2ecc;
         4'h9c08 	:	val_out <= 4'h2eb8;
         4'h9c09 	:	val_out <= 4'h2eb8;
         4'h9c0a 	:	val_out <= 4'h2eb8;
         4'h9c0b 	:	val_out <= 4'h2eb8;
         4'h9c10 	:	val_out <= 4'h2ea5;
         4'h9c11 	:	val_out <= 4'h2ea5;
         4'h9c12 	:	val_out <= 4'h2ea5;
         4'h9c13 	:	val_out <= 4'h2ea5;
         4'h9c18 	:	val_out <= 4'h2e91;
         4'h9c19 	:	val_out <= 4'h2e91;
         4'h9c1a 	:	val_out <= 4'h2e91;
         4'h9c1b 	:	val_out <= 4'h2e91;
         4'h9c20 	:	val_out <= 4'h2e7e;
         4'h9c21 	:	val_out <= 4'h2e7e;
         4'h9c22 	:	val_out <= 4'h2e7e;
         4'h9c23 	:	val_out <= 4'h2e7e;
         4'h9c28 	:	val_out <= 4'h2e6b;
         4'h9c29 	:	val_out <= 4'h2e6b;
         4'h9c2a 	:	val_out <= 4'h2e6b;
         4'h9c2b 	:	val_out <= 4'h2e6b;
         4'h9c30 	:	val_out <= 4'h2e57;
         4'h9c31 	:	val_out <= 4'h2e57;
         4'h9c32 	:	val_out <= 4'h2e57;
         4'h9c33 	:	val_out <= 4'h2e57;
         4'h9c38 	:	val_out <= 4'h2e44;
         4'h9c39 	:	val_out <= 4'h2e44;
         4'h9c3a 	:	val_out <= 4'h2e44;
         4'h9c3b 	:	val_out <= 4'h2e44;
         4'h9c40 	:	val_out <= 4'h2e31;
         4'h9c41 	:	val_out <= 4'h2e31;
         4'h9c42 	:	val_out <= 4'h2e31;
         4'h9c43 	:	val_out <= 4'h2e31;
         4'h9c48 	:	val_out <= 4'h2e1d;
         4'h9c49 	:	val_out <= 4'h2e1d;
         4'h9c4a 	:	val_out <= 4'h2e1d;
         4'h9c4b 	:	val_out <= 4'h2e1d;
         4'h9c50 	:	val_out <= 4'h2e0a;
         4'h9c51 	:	val_out <= 4'h2e0a;
         4'h9c52 	:	val_out <= 4'h2e0a;
         4'h9c53 	:	val_out <= 4'h2e0a;
         4'h9c58 	:	val_out <= 4'h2df7;
         4'h9c59 	:	val_out <= 4'h2df7;
         4'h9c5a 	:	val_out <= 4'h2df7;
         4'h9c5b 	:	val_out <= 4'h2df7;
         4'h9c60 	:	val_out <= 4'h2de3;
         4'h9c61 	:	val_out <= 4'h2de3;
         4'h9c62 	:	val_out <= 4'h2de3;
         4'h9c63 	:	val_out <= 4'h2de3;
         4'h9c68 	:	val_out <= 4'h2dd0;
         4'h9c69 	:	val_out <= 4'h2dd0;
         4'h9c6a 	:	val_out <= 4'h2dd0;
         4'h9c6b 	:	val_out <= 4'h2dd0;
         4'h9c70 	:	val_out <= 4'h2dbd;
         4'h9c71 	:	val_out <= 4'h2dbd;
         4'h9c72 	:	val_out <= 4'h2dbd;
         4'h9c73 	:	val_out <= 4'h2dbd;
         4'h9c78 	:	val_out <= 4'h2daa;
         4'h9c79 	:	val_out <= 4'h2daa;
         4'h9c7a 	:	val_out <= 4'h2daa;
         4'h9c7b 	:	val_out <= 4'h2daa;
         4'h9c80 	:	val_out <= 4'h2d96;
         4'h9c81 	:	val_out <= 4'h2d96;
         4'h9c82 	:	val_out <= 4'h2d96;
         4'h9c83 	:	val_out <= 4'h2d96;
         4'h9c88 	:	val_out <= 4'h2d83;
         4'h9c89 	:	val_out <= 4'h2d83;
         4'h9c8a 	:	val_out <= 4'h2d83;
         4'h9c8b 	:	val_out <= 4'h2d83;
         4'h9c90 	:	val_out <= 4'h2d70;
         4'h9c91 	:	val_out <= 4'h2d70;
         4'h9c92 	:	val_out <= 4'h2d70;
         4'h9c93 	:	val_out <= 4'h2d70;
         4'h9c98 	:	val_out <= 4'h2d5d;
         4'h9c99 	:	val_out <= 4'h2d5d;
         4'h9c9a 	:	val_out <= 4'h2d5d;
         4'h9c9b 	:	val_out <= 4'h2d5d;
         4'h9ca0 	:	val_out <= 4'h2d4a;
         4'h9ca1 	:	val_out <= 4'h2d4a;
         4'h9ca2 	:	val_out <= 4'h2d4a;
         4'h9ca3 	:	val_out <= 4'h2d4a;
         4'h9ca8 	:	val_out <= 4'h2d36;
         4'h9ca9 	:	val_out <= 4'h2d36;
         4'h9caa 	:	val_out <= 4'h2d36;
         4'h9cab 	:	val_out <= 4'h2d36;
         4'h9cb0 	:	val_out <= 4'h2d23;
         4'h9cb1 	:	val_out <= 4'h2d23;
         4'h9cb2 	:	val_out <= 4'h2d23;
         4'h9cb3 	:	val_out <= 4'h2d23;
         4'h9cb8 	:	val_out <= 4'h2d10;
         4'h9cb9 	:	val_out <= 4'h2d10;
         4'h9cba 	:	val_out <= 4'h2d10;
         4'h9cbb 	:	val_out <= 4'h2d10;
         4'h9cc0 	:	val_out <= 4'h2cfd;
         4'h9cc1 	:	val_out <= 4'h2cfd;
         4'h9cc2 	:	val_out <= 4'h2cfd;
         4'h9cc3 	:	val_out <= 4'h2cfd;
         4'h9cc8 	:	val_out <= 4'h2cea;
         4'h9cc9 	:	val_out <= 4'h2cea;
         4'h9cca 	:	val_out <= 4'h2cea;
         4'h9ccb 	:	val_out <= 4'h2cea;
         4'h9cd0 	:	val_out <= 4'h2cd7;
         4'h9cd1 	:	val_out <= 4'h2cd7;
         4'h9cd2 	:	val_out <= 4'h2cd7;
         4'h9cd3 	:	val_out <= 4'h2cd7;
         4'h9cd8 	:	val_out <= 4'h2cc4;
         4'h9cd9 	:	val_out <= 4'h2cc4;
         4'h9cda 	:	val_out <= 4'h2cc4;
         4'h9cdb 	:	val_out <= 4'h2cc4;
         4'h9ce0 	:	val_out <= 4'h2cb1;
         4'h9ce1 	:	val_out <= 4'h2cb1;
         4'h9ce2 	:	val_out <= 4'h2cb1;
         4'h9ce3 	:	val_out <= 4'h2cb1;
         4'h9ce8 	:	val_out <= 4'h2c9d;
         4'h9ce9 	:	val_out <= 4'h2c9d;
         4'h9cea 	:	val_out <= 4'h2c9d;
         4'h9ceb 	:	val_out <= 4'h2c9d;
         4'h9cf0 	:	val_out <= 4'h2c8a;
         4'h9cf1 	:	val_out <= 4'h2c8a;
         4'h9cf2 	:	val_out <= 4'h2c8a;
         4'h9cf3 	:	val_out <= 4'h2c8a;
         4'h9cf8 	:	val_out <= 4'h2c77;
         4'h9cf9 	:	val_out <= 4'h2c77;
         4'h9cfa 	:	val_out <= 4'h2c77;
         4'h9cfb 	:	val_out <= 4'h2c77;
         4'h9d00 	:	val_out <= 4'h2c64;
         4'h9d01 	:	val_out <= 4'h2c64;
         4'h9d02 	:	val_out <= 4'h2c64;
         4'h9d03 	:	val_out <= 4'h2c64;
         4'h9d08 	:	val_out <= 4'h2c51;
         4'h9d09 	:	val_out <= 4'h2c51;
         4'h9d0a 	:	val_out <= 4'h2c51;
         4'h9d0b 	:	val_out <= 4'h2c51;
         4'h9d10 	:	val_out <= 4'h2c3e;
         4'h9d11 	:	val_out <= 4'h2c3e;
         4'h9d12 	:	val_out <= 4'h2c3e;
         4'h9d13 	:	val_out <= 4'h2c3e;
         4'h9d18 	:	val_out <= 4'h2c2b;
         4'h9d19 	:	val_out <= 4'h2c2b;
         4'h9d1a 	:	val_out <= 4'h2c2b;
         4'h9d1b 	:	val_out <= 4'h2c2b;
         4'h9d20 	:	val_out <= 4'h2c18;
         4'h9d21 	:	val_out <= 4'h2c18;
         4'h9d22 	:	val_out <= 4'h2c18;
         4'h9d23 	:	val_out <= 4'h2c18;
         4'h9d28 	:	val_out <= 4'h2c05;
         4'h9d29 	:	val_out <= 4'h2c05;
         4'h9d2a 	:	val_out <= 4'h2c05;
         4'h9d2b 	:	val_out <= 4'h2c05;
         4'h9d30 	:	val_out <= 4'h2bf2;
         4'h9d31 	:	val_out <= 4'h2bf2;
         4'h9d32 	:	val_out <= 4'h2bf2;
         4'h9d33 	:	val_out <= 4'h2bf2;
         4'h9d38 	:	val_out <= 4'h2bdf;
         4'h9d39 	:	val_out <= 4'h2bdf;
         4'h9d3a 	:	val_out <= 4'h2bdf;
         4'h9d3b 	:	val_out <= 4'h2bdf;
         4'h9d40 	:	val_out <= 4'h2bcc;
         4'h9d41 	:	val_out <= 4'h2bcc;
         4'h9d42 	:	val_out <= 4'h2bcc;
         4'h9d43 	:	val_out <= 4'h2bcc;
         4'h9d48 	:	val_out <= 4'h2bba;
         4'h9d49 	:	val_out <= 4'h2bba;
         4'h9d4a 	:	val_out <= 4'h2bba;
         4'h9d4b 	:	val_out <= 4'h2bba;
         4'h9d50 	:	val_out <= 4'h2ba7;
         4'h9d51 	:	val_out <= 4'h2ba7;
         4'h9d52 	:	val_out <= 4'h2ba7;
         4'h9d53 	:	val_out <= 4'h2ba7;
         4'h9d58 	:	val_out <= 4'h2b94;
         4'h9d59 	:	val_out <= 4'h2b94;
         4'h9d5a 	:	val_out <= 4'h2b94;
         4'h9d5b 	:	val_out <= 4'h2b94;
         4'h9d60 	:	val_out <= 4'h2b81;
         4'h9d61 	:	val_out <= 4'h2b81;
         4'h9d62 	:	val_out <= 4'h2b81;
         4'h9d63 	:	val_out <= 4'h2b81;
         4'h9d68 	:	val_out <= 4'h2b6e;
         4'h9d69 	:	val_out <= 4'h2b6e;
         4'h9d6a 	:	val_out <= 4'h2b6e;
         4'h9d6b 	:	val_out <= 4'h2b6e;
         4'h9d70 	:	val_out <= 4'h2b5b;
         4'h9d71 	:	val_out <= 4'h2b5b;
         4'h9d72 	:	val_out <= 4'h2b5b;
         4'h9d73 	:	val_out <= 4'h2b5b;
         4'h9d78 	:	val_out <= 4'h2b48;
         4'h9d79 	:	val_out <= 4'h2b48;
         4'h9d7a 	:	val_out <= 4'h2b48;
         4'h9d7b 	:	val_out <= 4'h2b48;
         4'h9d80 	:	val_out <= 4'h2b35;
         4'h9d81 	:	val_out <= 4'h2b35;
         4'h9d82 	:	val_out <= 4'h2b35;
         4'h9d83 	:	val_out <= 4'h2b35;
         4'h9d88 	:	val_out <= 4'h2b23;
         4'h9d89 	:	val_out <= 4'h2b23;
         4'h9d8a 	:	val_out <= 4'h2b23;
         4'h9d8b 	:	val_out <= 4'h2b23;
         4'h9d90 	:	val_out <= 4'h2b10;
         4'h9d91 	:	val_out <= 4'h2b10;
         4'h9d92 	:	val_out <= 4'h2b10;
         4'h9d93 	:	val_out <= 4'h2b10;
         4'h9d98 	:	val_out <= 4'h2afd;
         4'h9d99 	:	val_out <= 4'h2afd;
         4'h9d9a 	:	val_out <= 4'h2afd;
         4'h9d9b 	:	val_out <= 4'h2afd;
         4'h9da0 	:	val_out <= 4'h2aea;
         4'h9da1 	:	val_out <= 4'h2aea;
         4'h9da2 	:	val_out <= 4'h2aea;
         4'h9da3 	:	val_out <= 4'h2aea;
         4'h9da8 	:	val_out <= 4'h2ad7;
         4'h9da9 	:	val_out <= 4'h2ad7;
         4'h9daa 	:	val_out <= 4'h2ad7;
         4'h9dab 	:	val_out <= 4'h2ad7;
         4'h9db0 	:	val_out <= 4'h2ac5;
         4'h9db1 	:	val_out <= 4'h2ac5;
         4'h9db2 	:	val_out <= 4'h2ac5;
         4'h9db3 	:	val_out <= 4'h2ac5;
         4'h9db8 	:	val_out <= 4'h2ab2;
         4'h9db9 	:	val_out <= 4'h2ab2;
         4'h9dba 	:	val_out <= 4'h2ab2;
         4'h9dbb 	:	val_out <= 4'h2ab2;
         4'h9dc0 	:	val_out <= 4'h2a9f;
         4'h9dc1 	:	val_out <= 4'h2a9f;
         4'h9dc2 	:	val_out <= 4'h2a9f;
         4'h9dc3 	:	val_out <= 4'h2a9f;
         4'h9dc8 	:	val_out <= 4'h2a8d;
         4'h9dc9 	:	val_out <= 4'h2a8d;
         4'h9dca 	:	val_out <= 4'h2a8d;
         4'h9dcb 	:	val_out <= 4'h2a8d;
         4'h9dd0 	:	val_out <= 4'h2a7a;
         4'h9dd1 	:	val_out <= 4'h2a7a;
         4'h9dd2 	:	val_out <= 4'h2a7a;
         4'h9dd3 	:	val_out <= 4'h2a7a;
         4'h9dd8 	:	val_out <= 4'h2a67;
         4'h9dd9 	:	val_out <= 4'h2a67;
         4'h9dda 	:	val_out <= 4'h2a67;
         4'h9ddb 	:	val_out <= 4'h2a67;
         4'h9de0 	:	val_out <= 4'h2a54;
         4'h9de1 	:	val_out <= 4'h2a54;
         4'h9de2 	:	val_out <= 4'h2a54;
         4'h9de3 	:	val_out <= 4'h2a54;
         4'h9de8 	:	val_out <= 4'h2a42;
         4'h9de9 	:	val_out <= 4'h2a42;
         4'h9dea 	:	val_out <= 4'h2a42;
         4'h9deb 	:	val_out <= 4'h2a42;
         4'h9df0 	:	val_out <= 4'h2a2f;
         4'h9df1 	:	val_out <= 4'h2a2f;
         4'h9df2 	:	val_out <= 4'h2a2f;
         4'h9df3 	:	val_out <= 4'h2a2f;
         4'h9df8 	:	val_out <= 4'h2a1c;
         4'h9df9 	:	val_out <= 4'h2a1c;
         4'h9dfa 	:	val_out <= 4'h2a1c;
         4'h9dfb 	:	val_out <= 4'h2a1c;
         4'h9e00 	:	val_out <= 4'h2a0a;
         4'h9e01 	:	val_out <= 4'h2a0a;
         4'h9e02 	:	val_out <= 4'h2a0a;
         4'h9e03 	:	val_out <= 4'h2a0a;
         4'h9e08 	:	val_out <= 4'h29f7;
         4'h9e09 	:	val_out <= 4'h29f7;
         4'h9e0a 	:	val_out <= 4'h29f7;
         4'h9e0b 	:	val_out <= 4'h29f7;
         4'h9e10 	:	val_out <= 4'h29e5;
         4'h9e11 	:	val_out <= 4'h29e5;
         4'h9e12 	:	val_out <= 4'h29e5;
         4'h9e13 	:	val_out <= 4'h29e5;
         4'h9e18 	:	val_out <= 4'h29d2;
         4'h9e19 	:	val_out <= 4'h29d2;
         4'h9e1a 	:	val_out <= 4'h29d2;
         4'h9e1b 	:	val_out <= 4'h29d2;
         4'h9e20 	:	val_out <= 4'h29bf;
         4'h9e21 	:	val_out <= 4'h29bf;
         4'h9e22 	:	val_out <= 4'h29bf;
         4'h9e23 	:	val_out <= 4'h29bf;
         4'h9e28 	:	val_out <= 4'h29ad;
         4'h9e29 	:	val_out <= 4'h29ad;
         4'h9e2a 	:	val_out <= 4'h29ad;
         4'h9e2b 	:	val_out <= 4'h29ad;
         4'h9e30 	:	val_out <= 4'h299a;
         4'h9e31 	:	val_out <= 4'h299a;
         4'h9e32 	:	val_out <= 4'h299a;
         4'h9e33 	:	val_out <= 4'h299a;
         4'h9e38 	:	val_out <= 4'h2988;
         4'h9e39 	:	val_out <= 4'h2988;
         4'h9e3a 	:	val_out <= 4'h2988;
         4'h9e3b 	:	val_out <= 4'h2988;
         4'h9e40 	:	val_out <= 4'h2975;
         4'h9e41 	:	val_out <= 4'h2975;
         4'h9e42 	:	val_out <= 4'h2975;
         4'h9e43 	:	val_out <= 4'h2975;
         4'h9e48 	:	val_out <= 4'h2963;
         4'h9e49 	:	val_out <= 4'h2963;
         4'h9e4a 	:	val_out <= 4'h2963;
         4'h9e4b 	:	val_out <= 4'h2963;
         4'h9e50 	:	val_out <= 4'h2950;
         4'h9e51 	:	val_out <= 4'h2950;
         4'h9e52 	:	val_out <= 4'h2950;
         4'h9e53 	:	val_out <= 4'h2950;
         4'h9e58 	:	val_out <= 4'h293e;
         4'h9e59 	:	val_out <= 4'h293e;
         4'h9e5a 	:	val_out <= 4'h293e;
         4'h9e5b 	:	val_out <= 4'h293e;
         4'h9e60 	:	val_out <= 4'h292b;
         4'h9e61 	:	val_out <= 4'h292b;
         4'h9e62 	:	val_out <= 4'h292b;
         4'h9e63 	:	val_out <= 4'h292b;
         4'h9e68 	:	val_out <= 4'h2919;
         4'h9e69 	:	val_out <= 4'h2919;
         4'h9e6a 	:	val_out <= 4'h2919;
         4'h9e6b 	:	val_out <= 4'h2919;
         4'h9e70 	:	val_out <= 4'h2906;
         4'h9e71 	:	val_out <= 4'h2906;
         4'h9e72 	:	val_out <= 4'h2906;
         4'h9e73 	:	val_out <= 4'h2906;
         4'h9e78 	:	val_out <= 4'h28f4;
         4'h9e79 	:	val_out <= 4'h28f4;
         4'h9e7a 	:	val_out <= 4'h28f4;
         4'h9e7b 	:	val_out <= 4'h28f4;
         4'h9e80 	:	val_out <= 4'h28e2;
         4'h9e81 	:	val_out <= 4'h28e2;
         4'h9e82 	:	val_out <= 4'h28e2;
         4'h9e83 	:	val_out <= 4'h28e2;
         4'h9e88 	:	val_out <= 4'h28cf;
         4'h9e89 	:	val_out <= 4'h28cf;
         4'h9e8a 	:	val_out <= 4'h28cf;
         4'h9e8b 	:	val_out <= 4'h28cf;
         4'h9e90 	:	val_out <= 4'h28bd;
         4'h9e91 	:	val_out <= 4'h28bd;
         4'h9e92 	:	val_out <= 4'h28bd;
         4'h9e93 	:	val_out <= 4'h28bd;
         4'h9e98 	:	val_out <= 4'h28aa;
         4'h9e99 	:	val_out <= 4'h28aa;
         4'h9e9a 	:	val_out <= 4'h28aa;
         4'h9e9b 	:	val_out <= 4'h28aa;
         4'h9ea0 	:	val_out <= 4'h2898;
         4'h9ea1 	:	val_out <= 4'h2898;
         4'h9ea2 	:	val_out <= 4'h2898;
         4'h9ea3 	:	val_out <= 4'h2898;
         4'h9ea8 	:	val_out <= 4'h2886;
         4'h9ea9 	:	val_out <= 4'h2886;
         4'h9eaa 	:	val_out <= 4'h2886;
         4'h9eab 	:	val_out <= 4'h2886;
         4'h9eb0 	:	val_out <= 4'h2873;
         4'h9eb1 	:	val_out <= 4'h2873;
         4'h9eb2 	:	val_out <= 4'h2873;
         4'h9eb3 	:	val_out <= 4'h2873;
         4'h9eb8 	:	val_out <= 4'h2861;
         4'h9eb9 	:	val_out <= 4'h2861;
         4'h9eba 	:	val_out <= 4'h2861;
         4'h9ebb 	:	val_out <= 4'h2861;
         4'h9ec0 	:	val_out <= 4'h284f;
         4'h9ec1 	:	val_out <= 4'h284f;
         4'h9ec2 	:	val_out <= 4'h284f;
         4'h9ec3 	:	val_out <= 4'h284f;
         4'h9ec8 	:	val_out <= 4'h283c;
         4'h9ec9 	:	val_out <= 4'h283c;
         4'h9eca 	:	val_out <= 4'h283c;
         4'h9ecb 	:	val_out <= 4'h283c;
         4'h9ed0 	:	val_out <= 4'h282a;
         4'h9ed1 	:	val_out <= 4'h282a;
         4'h9ed2 	:	val_out <= 4'h282a;
         4'h9ed3 	:	val_out <= 4'h282a;
         4'h9ed8 	:	val_out <= 4'h2818;
         4'h9ed9 	:	val_out <= 4'h2818;
         4'h9eda 	:	val_out <= 4'h2818;
         4'h9edb 	:	val_out <= 4'h2818;
         4'h9ee0 	:	val_out <= 4'h2806;
         4'h9ee1 	:	val_out <= 4'h2806;
         4'h9ee2 	:	val_out <= 4'h2806;
         4'h9ee3 	:	val_out <= 4'h2806;
         4'h9ee8 	:	val_out <= 4'h27f3;
         4'h9ee9 	:	val_out <= 4'h27f3;
         4'h9eea 	:	val_out <= 4'h27f3;
         4'h9eeb 	:	val_out <= 4'h27f3;
         4'h9ef0 	:	val_out <= 4'h27e1;
         4'h9ef1 	:	val_out <= 4'h27e1;
         4'h9ef2 	:	val_out <= 4'h27e1;
         4'h9ef3 	:	val_out <= 4'h27e1;
         4'h9ef8 	:	val_out <= 4'h27cf;
         4'h9ef9 	:	val_out <= 4'h27cf;
         4'h9efa 	:	val_out <= 4'h27cf;
         4'h9efb 	:	val_out <= 4'h27cf;
         4'h9f00 	:	val_out <= 4'h27bd;
         4'h9f01 	:	val_out <= 4'h27bd;
         4'h9f02 	:	val_out <= 4'h27bd;
         4'h9f03 	:	val_out <= 4'h27bd;
         4'h9f08 	:	val_out <= 4'h27aa;
         4'h9f09 	:	val_out <= 4'h27aa;
         4'h9f0a 	:	val_out <= 4'h27aa;
         4'h9f0b 	:	val_out <= 4'h27aa;
         4'h9f10 	:	val_out <= 4'h2798;
         4'h9f11 	:	val_out <= 4'h2798;
         4'h9f12 	:	val_out <= 4'h2798;
         4'h9f13 	:	val_out <= 4'h2798;
         4'h9f18 	:	val_out <= 4'h2786;
         4'h9f19 	:	val_out <= 4'h2786;
         4'h9f1a 	:	val_out <= 4'h2786;
         4'h9f1b 	:	val_out <= 4'h2786;
         4'h9f20 	:	val_out <= 4'h2774;
         4'h9f21 	:	val_out <= 4'h2774;
         4'h9f22 	:	val_out <= 4'h2774;
         4'h9f23 	:	val_out <= 4'h2774;
         4'h9f28 	:	val_out <= 4'h2762;
         4'h9f29 	:	val_out <= 4'h2762;
         4'h9f2a 	:	val_out <= 4'h2762;
         4'h9f2b 	:	val_out <= 4'h2762;
         4'h9f30 	:	val_out <= 4'h2750;
         4'h9f31 	:	val_out <= 4'h2750;
         4'h9f32 	:	val_out <= 4'h2750;
         4'h9f33 	:	val_out <= 4'h2750;
         4'h9f38 	:	val_out <= 4'h273e;
         4'h9f39 	:	val_out <= 4'h273e;
         4'h9f3a 	:	val_out <= 4'h273e;
         4'h9f3b 	:	val_out <= 4'h273e;
         4'h9f40 	:	val_out <= 4'h272b;
         4'h9f41 	:	val_out <= 4'h272b;
         4'h9f42 	:	val_out <= 4'h272b;
         4'h9f43 	:	val_out <= 4'h272b;
         4'h9f48 	:	val_out <= 4'h2719;
         4'h9f49 	:	val_out <= 4'h2719;
         4'h9f4a 	:	val_out <= 4'h2719;
         4'h9f4b 	:	val_out <= 4'h2719;
         4'h9f50 	:	val_out <= 4'h2707;
         4'h9f51 	:	val_out <= 4'h2707;
         4'h9f52 	:	val_out <= 4'h2707;
         4'h9f53 	:	val_out <= 4'h2707;
         4'h9f58 	:	val_out <= 4'h26f5;
         4'h9f59 	:	val_out <= 4'h26f5;
         4'h9f5a 	:	val_out <= 4'h26f5;
         4'h9f5b 	:	val_out <= 4'h26f5;
         4'h9f60 	:	val_out <= 4'h26e3;
         4'h9f61 	:	val_out <= 4'h26e3;
         4'h9f62 	:	val_out <= 4'h26e3;
         4'h9f63 	:	val_out <= 4'h26e3;
         4'h9f68 	:	val_out <= 4'h26d1;
         4'h9f69 	:	val_out <= 4'h26d1;
         4'h9f6a 	:	val_out <= 4'h26d1;
         4'h9f6b 	:	val_out <= 4'h26d1;
         4'h9f70 	:	val_out <= 4'h26bf;
         4'h9f71 	:	val_out <= 4'h26bf;
         4'h9f72 	:	val_out <= 4'h26bf;
         4'h9f73 	:	val_out <= 4'h26bf;
         4'h9f78 	:	val_out <= 4'h26ad;
         4'h9f79 	:	val_out <= 4'h26ad;
         4'h9f7a 	:	val_out <= 4'h26ad;
         4'h9f7b 	:	val_out <= 4'h26ad;
         4'h9f80 	:	val_out <= 4'h269b;
         4'h9f81 	:	val_out <= 4'h269b;
         4'h9f82 	:	val_out <= 4'h269b;
         4'h9f83 	:	val_out <= 4'h269b;
         4'h9f88 	:	val_out <= 4'h2689;
         4'h9f89 	:	val_out <= 4'h2689;
         4'h9f8a 	:	val_out <= 4'h2689;
         4'h9f8b 	:	val_out <= 4'h2689;
         4'h9f90 	:	val_out <= 4'h2677;
         4'h9f91 	:	val_out <= 4'h2677;
         4'h9f92 	:	val_out <= 4'h2677;
         4'h9f93 	:	val_out <= 4'h2677;
         4'h9f98 	:	val_out <= 4'h2665;
         4'h9f99 	:	val_out <= 4'h2665;
         4'h9f9a 	:	val_out <= 4'h2665;
         4'h9f9b 	:	val_out <= 4'h2665;
         4'h9fa0 	:	val_out <= 4'h2653;
         4'h9fa1 	:	val_out <= 4'h2653;
         4'h9fa2 	:	val_out <= 4'h2653;
         4'h9fa3 	:	val_out <= 4'h2653;
         4'h9fa8 	:	val_out <= 4'h2641;
         4'h9fa9 	:	val_out <= 4'h2641;
         4'h9faa 	:	val_out <= 4'h2641;
         4'h9fab 	:	val_out <= 4'h2641;
         4'h9fb0 	:	val_out <= 4'h262f;
         4'h9fb1 	:	val_out <= 4'h262f;
         4'h9fb2 	:	val_out <= 4'h262f;
         4'h9fb3 	:	val_out <= 4'h262f;
         4'h9fb8 	:	val_out <= 4'h261e;
         4'h9fb9 	:	val_out <= 4'h261e;
         4'h9fba 	:	val_out <= 4'h261e;
         4'h9fbb 	:	val_out <= 4'h261e;
         4'h9fc0 	:	val_out <= 4'h260c;
         4'h9fc1 	:	val_out <= 4'h260c;
         4'h9fc2 	:	val_out <= 4'h260c;
         4'h9fc3 	:	val_out <= 4'h260c;
         4'h9fc8 	:	val_out <= 4'h25fa;
         4'h9fc9 	:	val_out <= 4'h25fa;
         4'h9fca 	:	val_out <= 4'h25fa;
         4'h9fcb 	:	val_out <= 4'h25fa;
         4'h9fd0 	:	val_out <= 4'h25e8;
         4'h9fd1 	:	val_out <= 4'h25e8;
         4'h9fd2 	:	val_out <= 4'h25e8;
         4'h9fd3 	:	val_out <= 4'h25e8;
         4'h9fd8 	:	val_out <= 4'h25d6;
         4'h9fd9 	:	val_out <= 4'h25d6;
         4'h9fda 	:	val_out <= 4'h25d6;
         4'h9fdb 	:	val_out <= 4'h25d6;
         4'h9fe0 	:	val_out <= 4'h25c4;
         4'h9fe1 	:	val_out <= 4'h25c4;
         4'h9fe2 	:	val_out <= 4'h25c4;
         4'h9fe3 	:	val_out <= 4'h25c4;
         4'h9fe8 	:	val_out <= 4'h25b2;
         4'h9fe9 	:	val_out <= 4'h25b2;
         4'h9fea 	:	val_out <= 4'h25b2;
         4'h9feb 	:	val_out <= 4'h25b2;
         4'h9ff0 	:	val_out <= 4'h25a1;
         4'h9ff1 	:	val_out <= 4'h25a1;
         4'h9ff2 	:	val_out <= 4'h25a1;
         4'h9ff3 	:	val_out <= 4'h25a1;
         4'h9ff8 	:	val_out <= 4'h258f;
         4'h9ff9 	:	val_out <= 4'h258f;
         4'h9ffa 	:	val_out <= 4'h258f;
         4'h9ffb 	:	val_out <= 4'h258f;
         4'ha000 	:	val_out <= 4'h257d;
         4'ha001 	:	val_out <= 4'h257d;
         4'ha002 	:	val_out <= 4'h257d;
         4'ha003 	:	val_out <= 4'h257d;
         4'ha008 	:	val_out <= 4'h256b;
         4'ha009 	:	val_out <= 4'h256b;
         4'ha00a 	:	val_out <= 4'h256b;
         4'ha00b 	:	val_out <= 4'h256b;
         4'ha010 	:	val_out <= 4'h255a;
         4'ha011 	:	val_out <= 4'h255a;
         4'ha012 	:	val_out <= 4'h255a;
         4'ha013 	:	val_out <= 4'h255a;
         4'ha018 	:	val_out <= 4'h2548;
         4'ha019 	:	val_out <= 4'h2548;
         4'ha01a 	:	val_out <= 4'h2548;
         4'ha01b 	:	val_out <= 4'h2548;
         4'ha020 	:	val_out <= 4'h2536;
         4'ha021 	:	val_out <= 4'h2536;
         4'ha022 	:	val_out <= 4'h2536;
         4'ha023 	:	val_out <= 4'h2536;
         4'ha028 	:	val_out <= 4'h2524;
         4'ha029 	:	val_out <= 4'h2524;
         4'ha02a 	:	val_out <= 4'h2524;
         4'ha02b 	:	val_out <= 4'h2524;
         4'ha030 	:	val_out <= 4'h2513;
         4'ha031 	:	val_out <= 4'h2513;
         4'ha032 	:	val_out <= 4'h2513;
         4'ha033 	:	val_out <= 4'h2513;
         4'ha038 	:	val_out <= 4'h2501;
         4'ha039 	:	val_out <= 4'h2501;
         4'ha03a 	:	val_out <= 4'h2501;
         4'ha03b 	:	val_out <= 4'h2501;
         4'ha040 	:	val_out <= 4'h24ef;
         4'ha041 	:	val_out <= 4'h24ef;
         4'ha042 	:	val_out <= 4'h24ef;
         4'ha043 	:	val_out <= 4'h24ef;
         4'ha048 	:	val_out <= 4'h24de;
         4'ha049 	:	val_out <= 4'h24de;
         4'ha04a 	:	val_out <= 4'h24de;
         4'ha04b 	:	val_out <= 4'h24de;
         4'ha050 	:	val_out <= 4'h24cc;
         4'ha051 	:	val_out <= 4'h24cc;
         4'ha052 	:	val_out <= 4'h24cc;
         4'ha053 	:	val_out <= 4'h24cc;
         4'ha058 	:	val_out <= 4'h24ba;
         4'ha059 	:	val_out <= 4'h24ba;
         4'ha05a 	:	val_out <= 4'h24ba;
         4'ha05b 	:	val_out <= 4'h24ba;
         4'ha060 	:	val_out <= 4'h24a9;
         4'ha061 	:	val_out <= 4'h24a9;
         4'ha062 	:	val_out <= 4'h24a9;
         4'ha063 	:	val_out <= 4'h24a9;
         4'ha068 	:	val_out <= 4'h2497;
         4'ha069 	:	val_out <= 4'h2497;
         4'ha06a 	:	val_out <= 4'h2497;
         4'ha06b 	:	val_out <= 4'h2497;
         4'ha070 	:	val_out <= 4'h2486;
         4'ha071 	:	val_out <= 4'h2486;
         4'ha072 	:	val_out <= 4'h2486;
         4'ha073 	:	val_out <= 4'h2486;
         4'ha078 	:	val_out <= 4'h2474;
         4'ha079 	:	val_out <= 4'h2474;
         4'ha07a 	:	val_out <= 4'h2474;
         4'ha07b 	:	val_out <= 4'h2474;
         4'ha080 	:	val_out <= 4'h2462;
         4'ha081 	:	val_out <= 4'h2462;
         4'ha082 	:	val_out <= 4'h2462;
         4'ha083 	:	val_out <= 4'h2462;
         4'ha088 	:	val_out <= 4'h2451;
         4'ha089 	:	val_out <= 4'h2451;
         4'ha08a 	:	val_out <= 4'h2451;
         4'ha08b 	:	val_out <= 4'h2451;
         4'ha090 	:	val_out <= 4'h243f;
         4'ha091 	:	val_out <= 4'h243f;
         4'ha092 	:	val_out <= 4'h243f;
         4'ha093 	:	val_out <= 4'h243f;
         4'ha098 	:	val_out <= 4'h242e;
         4'ha099 	:	val_out <= 4'h242e;
         4'ha09a 	:	val_out <= 4'h242e;
         4'ha09b 	:	val_out <= 4'h242e;
         4'ha0a0 	:	val_out <= 4'h241c;
         4'ha0a1 	:	val_out <= 4'h241c;
         4'ha0a2 	:	val_out <= 4'h241c;
         4'ha0a3 	:	val_out <= 4'h241c;
         4'ha0a8 	:	val_out <= 4'h240b;
         4'ha0a9 	:	val_out <= 4'h240b;
         4'ha0aa 	:	val_out <= 4'h240b;
         4'ha0ab 	:	val_out <= 4'h240b;
         4'ha0b0 	:	val_out <= 4'h23f9;
         4'ha0b1 	:	val_out <= 4'h23f9;
         4'ha0b2 	:	val_out <= 4'h23f9;
         4'ha0b3 	:	val_out <= 4'h23f9;
         4'ha0b8 	:	val_out <= 4'h23e8;
         4'ha0b9 	:	val_out <= 4'h23e8;
         4'ha0ba 	:	val_out <= 4'h23e8;
         4'ha0bb 	:	val_out <= 4'h23e8;
         4'ha0c0 	:	val_out <= 4'h23d6;
         4'ha0c1 	:	val_out <= 4'h23d6;
         4'ha0c2 	:	val_out <= 4'h23d6;
         4'ha0c3 	:	val_out <= 4'h23d6;
         4'ha0c8 	:	val_out <= 4'h23c5;
         4'ha0c9 	:	val_out <= 4'h23c5;
         4'ha0ca 	:	val_out <= 4'h23c5;
         4'ha0cb 	:	val_out <= 4'h23c5;
         4'ha0d0 	:	val_out <= 4'h23b4;
         4'ha0d1 	:	val_out <= 4'h23b4;
         4'ha0d2 	:	val_out <= 4'h23b4;
         4'ha0d3 	:	val_out <= 4'h23b4;
         4'ha0d8 	:	val_out <= 4'h23a2;
         4'ha0d9 	:	val_out <= 4'h23a2;
         4'ha0da 	:	val_out <= 4'h23a2;
         4'ha0db 	:	val_out <= 4'h23a2;
         4'ha0e0 	:	val_out <= 4'h2391;
         4'ha0e1 	:	val_out <= 4'h2391;
         4'ha0e2 	:	val_out <= 4'h2391;
         4'ha0e3 	:	val_out <= 4'h2391;
         4'ha0e8 	:	val_out <= 4'h237f;
         4'ha0e9 	:	val_out <= 4'h237f;
         4'ha0ea 	:	val_out <= 4'h237f;
         4'ha0eb 	:	val_out <= 4'h237f;
         4'ha0f0 	:	val_out <= 4'h236e;
         4'ha0f1 	:	val_out <= 4'h236e;
         4'ha0f2 	:	val_out <= 4'h236e;
         4'ha0f3 	:	val_out <= 4'h236e;
         4'ha0f8 	:	val_out <= 4'h235d;
         4'ha0f9 	:	val_out <= 4'h235d;
         4'ha0fa 	:	val_out <= 4'h235d;
         4'ha0fb 	:	val_out <= 4'h235d;
         4'ha100 	:	val_out <= 4'h234b;
         4'ha101 	:	val_out <= 4'h234b;
         4'ha102 	:	val_out <= 4'h234b;
         4'ha103 	:	val_out <= 4'h234b;
         4'ha108 	:	val_out <= 4'h233a;
         4'ha109 	:	val_out <= 4'h233a;
         4'ha10a 	:	val_out <= 4'h233a;
         4'ha10b 	:	val_out <= 4'h233a;
         4'ha110 	:	val_out <= 4'h2329;
         4'ha111 	:	val_out <= 4'h2329;
         4'ha112 	:	val_out <= 4'h2329;
         4'ha113 	:	val_out <= 4'h2329;
         4'ha118 	:	val_out <= 4'h2317;
         4'ha119 	:	val_out <= 4'h2317;
         4'ha11a 	:	val_out <= 4'h2317;
         4'ha11b 	:	val_out <= 4'h2317;
         4'ha120 	:	val_out <= 4'h2306;
         4'ha121 	:	val_out <= 4'h2306;
         4'ha122 	:	val_out <= 4'h2306;
         4'ha123 	:	val_out <= 4'h2306;
         4'ha128 	:	val_out <= 4'h22f5;
         4'ha129 	:	val_out <= 4'h22f5;
         4'ha12a 	:	val_out <= 4'h22f5;
         4'ha12b 	:	val_out <= 4'h22f5;
         4'ha130 	:	val_out <= 4'h22e4;
         4'ha131 	:	val_out <= 4'h22e4;
         4'ha132 	:	val_out <= 4'h22e4;
         4'ha133 	:	val_out <= 4'h22e4;
         4'ha138 	:	val_out <= 4'h22d2;
         4'ha139 	:	val_out <= 4'h22d2;
         4'ha13a 	:	val_out <= 4'h22d2;
         4'ha13b 	:	val_out <= 4'h22d2;
         4'ha140 	:	val_out <= 4'h22c1;
         4'ha141 	:	val_out <= 4'h22c1;
         4'ha142 	:	val_out <= 4'h22c1;
         4'ha143 	:	val_out <= 4'h22c1;
         4'ha148 	:	val_out <= 4'h22b0;
         4'ha149 	:	val_out <= 4'h22b0;
         4'ha14a 	:	val_out <= 4'h22b0;
         4'ha14b 	:	val_out <= 4'h22b0;
         4'ha150 	:	val_out <= 4'h229f;
         4'ha151 	:	val_out <= 4'h229f;
         4'ha152 	:	val_out <= 4'h229f;
         4'ha153 	:	val_out <= 4'h229f;
         4'ha158 	:	val_out <= 4'h228e;
         4'ha159 	:	val_out <= 4'h228e;
         4'ha15a 	:	val_out <= 4'h228e;
         4'ha15b 	:	val_out <= 4'h228e;
         4'ha160 	:	val_out <= 4'h227c;
         4'ha161 	:	val_out <= 4'h227c;
         4'ha162 	:	val_out <= 4'h227c;
         4'ha163 	:	val_out <= 4'h227c;
         4'ha168 	:	val_out <= 4'h226b;
         4'ha169 	:	val_out <= 4'h226b;
         4'ha16a 	:	val_out <= 4'h226b;
         4'ha16b 	:	val_out <= 4'h226b;
         4'ha170 	:	val_out <= 4'h225a;
         4'ha171 	:	val_out <= 4'h225a;
         4'ha172 	:	val_out <= 4'h225a;
         4'ha173 	:	val_out <= 4'h225a;
         4'ha178 	:	val_out <= 4'h2249;
         4'ha179 	:	val_out <= 4'h2249;
         4'ha17a 	:	val_out <= 4'h2249;
         4'ha17b 	:	val_out <= 4'h2249;
         4'ha180 	:	val_out <= 4'h2238;
         4'ha181 	:	val_out <= 4'h2238;
         4'ha182 	:	val_out <= 4'h2238;
         4'ha183 	:	val_out <= 4'h2238;
         4'ha188 	:	val_out <= 4'h2227;
         4'ha189 	:	val_out <= 4'h2227;
         4'ha18a 	:	val_out <= 4'h2227;
         4'ha18b 	:	val_out <= 4'h2227;
         4'ha190 	:	val_out <= 4'h2216;
         4'ha191 	:	val_out <= 4'h2216;
         4'ha192 	:	val_out <= 4'h2216;
         4'ha193 	:	val_out <= 4'h2216;
         4'ha198 	:	val_out <= 4'h2205;
         4'ha199 	:	val_out <= 4'h2205;
         4'ha19a 	:	val_out <= 4'h2205;
         4'ha19b 	:	val_out <= 4'h2205;
         4'ha1a0 	:	val_out <= 4'h21f4;
         4'ha1a1 	:	val_out <= 4'h21f4;
         4'ha1a2 	:	val_out <= 4'h21f4;
         4'ha1a3 	:	val_out <= 4'h21f4;
         4'ha1a8 	:	val_out <= 4'h21e3;
         4'ha1a9 	:	val_out <= 4'h21e3;
         4'ha1aa 	:	val_out <= 4'h21e3;
         4'ha1ab 	:	val_out <= 4'h21e3;
         4'ha1b0 	:	val_out <= 4'h21d2;
         4'ha1b1 	:	val_out <= 4'h21d2;
         4'ha1b2 	:	val_out <= 4'h21d2;
         4'ha1b3 	:	val_out <= 4'h21d2;
         4'ha1b8 	:	val_out <= 4'h21c0;
         4'ha1b9 	:	val_out <= 4'h21c0;
         4'ha1ba 	:	val_out <= 4'h21c0;
         4'ha1bb 	:	val_out <= 4'h21c0;
         4'ha1c0 	:	val_out <= 4'h21af;
         4'ha1c1 	:	val_out <= 4'h21af;
         4'ha1c2 	:	val_out <= 4'h21af;
         4'ha1c3 	:	val_out <= 4'h21af;
         4'ha1c8 	:	val_out <= 4'h219f;
         4'ha1c9 	:	val_out <= 4'h219f;
         4'ha1ca 	:	val_out <= 4'h219f;
         4'ha1cb 	:	val_out <= 4'h219f;
         4'ha1d0 	:	val_out <= 4'h218e;
         4'ha1d1 	:	val_out <= 4'h218e;
         4'ha1d2 	:	val_out <= 4'h218e;
         4'ha1d3 	:	val_out <= 4'h218e;
         4'ha1d8 	:	val_out <= 4'h217d;
         4'ha1d9 	:	val_out <= 4'h217d;
         4'ha1da 	:	val_out <= 4'h217d;
         4'ha1db 	:	val_out <= 4'h217d;
         4'ha1e0 	:	val_out <= 4'h216c;
         4'ha1e1 	:	val_out <= 4'h216c;
         4'ha1e2 	:	val_out <= 4'h216c;
         4'ha1e3 	:	val_out <= 4'h216c;
         4'ha1e8 	:	val_out <= 4'h215b;
         4'ha1e9 	:	val_out <= 4'h215b;
         4'ha1ea 	:	val_out <= 4'h215b;
         4'ha1eb 	:	val_out <= 4'h215b;
         4'ha1f0 	:	val_out <= 4'h214a;
         4'ha1f1 	:	val_out <= 4'h214a;
         4'ha1f2 	:	val_out <= 4'h214a;
         4'ha1f3 	:	val_out <= 4'h214a;
         4'ha1f8 	:	val_out <= 4'h2139;
         4'ha1f9 	:	val_out <= 4'h2139;
         4'ha1fa 	:	val_out <= 4'h2139;
         4'ha1fb 	:	val_out <= 4'h2139;
         4'ha200 	:	val_out <= 4'h2128;
         4'ha201 	:	val_out <= 4'h2128;
         4'ha202 	:	val_out <= 4'h2128;
         4'ha203 	:	val_out <= 4'h2128;
         4'ha208 	:	val_out <= 4'h2117;
         4'ha209 	:	val_out <= 4'h2117;
         4'ha20a 	:	val_out <= 4'h2117;
         4'ha20b 	:	val_out <= 4'h2117;
         4'ha210 	:	val_out <= 4'h2106;
         4'ha211 	:	val_out <= 4'h2106;
         4'ha212 	:	val_out <= 4'h2106;
         4'ha213 	:	val_out <= 4'h2106;
         4'ha218 	:	val_out <= 4'h20f5;
         4'ha219 	:	val_out <= 4'h20f5;
         4'ha21a 	:	val_out <= 4'h20f5;
         4'ha21b 	:	val_out <= 4'h20f5;
         4'ha220 	:	val_out <= 4'h20e5;
         4'ha221 	:	val_out <= 4'h20e5;
         4'ha222 	:	val_out <= 4'h20e5;
         4'ha223 	:	val_out <= 4'h20e5;
         4'ha228 	:	val_out <= 4'h20d4;
         4'ha229 	:	val_out <= 4'h20d4;
         4'ha22a 	:	val_out <= 4'h20d4;
         4'ha22b 	:	val_out <= 4'h20d4;
         4'ha230 	:	val_out <= 4'h20c3;
         4'ha231 	:	val_out <= 4'h20c3;
         4'ha232 	:	val_out <= 4'h20c3;
         4'ha233 	:	val_out <= 4'h20c3;
         4'ha238 	:	val_out <= 4'h20b2;
         4'ha239 	:	val_out <= 4'h20b2;
         4'ha23a 	:	val_out <= 4'h20b2;
         4'ha23b 	:	val_out <= 4'h20b2;
         4'ha240 	:	val_out <= 4'h20a1;
         4'ha241 	:	val_out <= 4'h20a1;
         4'ha242 	:	val_out <= 4'h20a1;
         4'ha243 	:	val_out <= 4'h20a1;
         4'ha248 	:	val_out <= 4'h2091;
         4'ha249 	:	val_out <= 4'h2091;
         4'ha24a 	:	val_out <= 4'h2091;
         4'ha24b 	:	val_out <= 4'h2091;
         4'ha250 	:	val_out <= 4'h2080;
         4'ha251 	:	val_out <= 4'h2080;
         4'ha252 	:	val_out <= 4'h2080;
         4'ha253 	:	val_out <= 4'h2080;
         4'ha258 	:	val_out <= 4'h206f;
         4'ha259 	:	val_out <= 4'h206f;
         4'ha25a 	:	val_out <= 4'h206f;
         4'ha25b 	:	val_out <= 4'h206f;
         4'ha260 	:	val_out <= 4'h205f;
         4'ha261 	:	val_out <= 4'h205f;
         4'ha262 	:	val_out <= 4'h205f;
         4'ha263 	:	val_out <= 4'h205f;
         4'ha268 	:	val_out <= 4'h204e;
         4'ha269 	:	val_out <= 4'h204e;
         4'ha26a 	:	val_out <= 4'h204e;
         4'ha26b 	:	val_out <= 4'h204e;
         4'ha270 	:	val_out <= 4'h203d;
         4'ha271 	:	val_out <= 4'h203d;
         4'ha272 	:	val_out <= 4'h203d;
         4'ha273 	:	val_out <= 4'h203d;
         4'ha278 	:	val_out <= 4'h202c;
         4'ha279 	:	val_out <= 4'h202c;
         4'ha27a 	:	val_out <= 4'h202c;
         4'ha27b 	:	val_out <= 4'h202c;
         4'ha280 	:	val_out <= 4'h201c;
         4'ha281 	:	val_out <= 4'h201c;
         4'ha282 	:	val_out <= 4'h201c;
         4'ha283 	:	val_out <= 4'h201c;
         4'ha288 	:	val_out <= 4'h200b;
         4'ha289 	:	val_out <= 4'h200b;
         4'ha28a 	:	val_out <= 4'h200b;
         4'ha28b 	:	val_out <= 4'h200b;
         4'ha290 	:	val_out <= 4'h1ffb;
         4'ha291 	:	val_out <= 4'h1ffb;
         4'ha292 	:	val_out <= 4'h1ffb;
         4'ha293 	:	val_out <= 4'h1ffb;
         4'ha298 	:	val_out <= 4'h1fea;
         4'ha299 	:	val_out <= 4'h1fea;
         4'ha29a 	:	val_out <= 4'h1fea;
         4'ha29b 	:	val_out <= 4'h1fea;
         4'ha2a0 	:	val_out <= 4'h1fd9;
         4'ha2a1 	:	val_out <= 4'h1fd9;
         4'ha2a2 	:	val_out <= 4'h1fd9;
         4'ha2a3 	:	val_out <= 4'h1fd9;
         4'ha2a8 	:	val_out <= 4'h1fc9;
         4'ha2a9 	:	val_out <= 4'h1fc9;
         4'ha2aa 	:	val_out <= 4'h1fc9;
         4'ha2ab 	:	val_out <= 4'h1fc9;
         4'ha2b0 	:	val_out <= 4'h1fb8;
         4'ha2b1 	:	val_out <= 4'h1fb8;
         4'ha2b2 	:	val_out <= 4'h1fb8;
         4'ha2b3 	:	val_out <= 4'h1fb8;
         4'ha2b8 	:	val_out <= 4'h1fa8;
         4'ha2b9 	:	val_out <= 4'h1fa8;
         4'ha2ba 	:	val_out <= 4'h1fa8;
         4'ha2bb 	:	val_out <= 4'h1fa8;
         4'ha2c0 	:	val_out <= 4'h1f97;
         4'ha2c1 	:	val_out <= 4'h1f97;
         4'ha2c2 	:	val_out <= 4'h1f97;
         4'ha2c3 	:	val_out <= 4'h1f97;
         4'ha2c8 	:	val_out <= 4'h1f87;
         4'ha2c9 	:	val_out <= 4'h1f87;
         4'ha2ca 	:	val_out <= 4'h1f87;
         4'ha2cb 	:	val_out <= 4'h1f87;
         4'ha2d0 	:	val_out <= 4'h1f76;
         4'ha2d1 	:	val_out <= 4'h1f76;
         4'ha2d2 	:	val_out <= 4'h1f76;
         4'ha2d3 	:	val_out <= 4'h1f76;
         4'ha2d8 	:	val_out <= 4'h1f66;
         4'ha2d9 	:	val_out <= 4'h1f66;
         4'ha2da 	:	val_out <= 4'h1f66;
         4'ha2db 	:	val_out <= 4'h1f66;
         4'ha2e0 	:	val_out <= 4'h1f55;
         4'ha2e1 	:	val_out <= 4'h1f55;
         4'ha2e2 	:	val_out <= 4'h1f55;
         4'ha2e3 	:	val_out <= 4'h1f55;
         4'ha2e8 	:	val_out <= 4'h1f45;
         4'ha2e9 	:	val_out <= 4'h1f45;
         4'ha2ea 	:	val_out <= 4'h1f45;
         4'ha2eb 	:	val_out <= 4'h1f45;
         4'ha2f0 	:	val_out <= 4'h1f34;
         4'ha2f1 	:	val_out <= 4'h1f34;
         4'ha2f2 	:	val_out <= 4'h1f34;
         4'ha2f3 	:	val_out <= 4'h1f34;
         4'ha2f8 	:	val_out <= 4'h1f24;
         4'ha2f9 	:	val_out <= 4'h1f24;
         4'ha2fa 	:	val_out <= 4'h1f24;
         4'ha2fb 	:	val_out <= 4'h1f24;
         4'ha300 	:	val_out <= 4'h1f13;
         4'ha301 	:	val_out <= 4'h1f13;
         4'ha302 	:	val_out <= 4'h1f13;
         4'ha303 	:	val_out <= 4'h1f13;
         4'ha308 	:	val_out <= 4'h1f03;
         4'ha309 	:	val_out <= 4'h1f03;
         4'ha30a 	:	val_out <= 4'h1f03;
         4'ha30b 	:	val_out <= 4'h1f03;
         4'ha310 	:	val_out <= 4'h1ef2;
         4'ha311 	:	val_out <= 4'h1ef2;
         4'ha312 	:	val_out <= 4'h1ef2;
         4'ha313 	:	val_out <= 4'h1ef2;
         4'ha318 	:	val_out <= 4'h1ee2;
         4'ha319 	:	val_out <= 4'h1ee2;
         4'ha31a 	:	val_out <= 4'h1ee2;
         4'ha31b 	:	val_out <= 4'h1ee2;
         4'ha320 	:	val_out <= 4'h1ed2;
         4'ha321 	:	val_out <= 4'h1ed2;
         4'ha322 	:	val_out <= 4'h1ed2;
         4'ha323 	:	val_out <= 4'h1ed2;
         4'ha328 	:	val_out <= 4'h1ec1;
         4'ha329 	:	val_out <= 4'h1ec1;
         4'ha32a 	:	val_out <= 4'h1ec1;
         4'ha32b 	:	val_out <= 4'h1ec1;
         4'ha330 	:	val_out <= 4'h1eb1;
         4'ha331 	:	val_out <= 4'h1eb1;
         4'ha332 	:	val_out <= 4'h1eb1;
         4'ha333 	:	val_out <= 4'h1eb1;
         4'ha338 	:	val_out <= 4'h1ea1;
         4'ha339 	:	val_out <= 4'h1ea1;
         4'ha33a 	:	val_out <= 4'h1ea1;
         4'ha33b 	:	val_out <= 4'h1ea1;
         4'ha340 	:	val_out <= 4'h1e90;
         4'ha341 	:	val_out <= 4'h1e90;
         4'ha342 	:	val_out <= 4'h1e90;
         4'ha343 	:	val_out <= 4'h1e90;
         4'ha348 	:	val_out <= 4'h1e80;
         4'ha349 	:	val_out <= 4'h1e80;
         4'ha34a 	:	val_out <= 4'h1e80;
         4'ha34b 	:	val_out <= 4'h1e80;
         4'ha350 	:	val_out <= 4'h1e70;
         4'ha351 	:	val_out <= 4'h1e70;
         4'ha352 	:	val_out <= 4'h1e70;
         4'ha353 	:	val_out <= 4'h1e70;
         4'ha358 	:	val_out <= 4'h1e60;
         4'ha359 	:	val_out <= 4'h1e60;
         4'ha35a 	:	val_out <= 4'h1e60;
         4'ha35b 	:	val_out <= 4'h1e60;
         4'ha360 	:	val_out <= 4'h1e4f;
         4'ha361 	:	val_out <= 4'h1e4f;
         4'ha362 	:	val_out <= 4'h1e4f;
         4'ha363 	:	val_out <= 4'h1e4f;
         4'ha368 	:	val_out <= 4'h1e3f;
         4'ha369 	:	val_out <= 4'h1e3f;
         4'ha36a 	:	val_out <= 4'h1e3f;
         4'ha36b 	:	val_out <= 4'h1e3f;
         4'ha370 	:	val_out <= 4'h1e2f;
         4'ha371 	:	val_out <= 4'h1e2f;
         4'ha372 	:	val_out <= 4'h1e2f;
         4'ha373 	:	val_out <= 4'h1e2f;
         4'ha378 	:	val_out <= 4'h1e1f;
         4'ha379 	:	val_out <= 4'h1e1f;
         4'ha37a 	:	val_out <= 4'h1e1f;
         4'ha37b 	:	val_out <= 4'h1e1f;
         4'ha380 	:	val_out <= 4'h1e0e;
         4'ha381 	:	val_out <= 4'h1e0e;
         4'ha382 	:	val_out <= 4'h1e0e;
         4'ha383 	:	val_out <= 4'h1e0e;
         4'ha388 	:	val_out <= 4'h1dfe;
         4'ha389 	:	val_out <= 4'h1dfe;
         4'ha38a 	:	val_out <= 4'h1dfe;
         4'ha38b 	:	val_out <= 4'h1dfe;
         4'ha390 	:	val_out <= 4'h1dee;
         4'ha391 	:	val_out <= 4'h1dee;
         4'ha392 	:	val_out <= 4'h1dee;
         4'ha393 	:	val_out <= 4'h1dee;
         4'ha398 	:	val_out <= 4'h1dde;
         4'ha399 	:	val_out <= 4'h1dde;
         4'ha39a 	:	val_out <= 4'h1dde;
         4'ha39b 	:	val_out <= 4'h1dde;
         4'ha3a0 	:	val_out <= 4'h1dce;
         4'ha3a1 	:	val_out <= 4'h1dce;
         4'ha3a2 	:	val_out <= 4'h1dce;
         4'ha3a3 	:	val_out <= 4'h1dce;
         4'ha3a8 	:	val_out <= 4'h1dbe;
         4'ha3a9 	:	val_out <= 4'h1dbe;
         4'ha3aa 	:	val_out <= 4'h1dbe;
         4'ha3ab 	:	val_out <= 4'h1dbe;
         4'ha3b0 	:	val_out <= 4'h1dae;
         4'ha3b1 	:	val_out <= 4'h1dae;
         4'ha3b2 	:	val_out <= 4'h1dae;
         4'ha3b3 	:	val_out <= 4'h1dae;
         4'ha3b8 	:	val_out <= 4'h1d9e;
         4'ha3b9 	:	val_out <= 4'h1d9e;
         4'ha3ba 	:	val_out <= 4'h1d9e;
         4'ha3bb 	:	val_out <= 4'h1d9e;
         4'ha3c0 	:	val_out <= 4'h1d8e;
         4'ha3c1 	:	val_out <= 4'h1d8e;
         4'ha3c2 	:	val_out <= 4'h1d8e;
         4'ha3c3 	:	val_out <= 4'h1d8e;
         4'ha3c8 	:	val_out <= 4'h1d7d;
         4'ha3c9 	:	val_out <= 4'h1d7d;
         4'ha3ca 	:	val_out <= 4'h1d7d;
         4'ha3cb 	:	val_out <= 4'h1d7d;
         4'ha3d0 	:	val_out <= 4'h1d6d;
         4'ha3d1 	:	val_out <= 4'h1d6d;
         4'ha3d2 	:	val_out <= 4'h1d6d;
         4'ha3d3 	:	val_out <= 4'h1d6d;
         4'ha3d8 	:	val_out <= 4'h1d5d;
         4'ha3d9 	:	val_out <= 4'h1d5d;
         4'ha3da 	:	val_out <= 4'h1d5d;
         4'ha3db 	:	val_out <= 4'h1d5d;
         4'ha3e0 	:	val_out <= 4'h1d4d;
         4'ha3e1 	:	val_out <= 4'h1d4d;
         4'ha3e2 	:	val_out <= 4'h1d4d;
         4'ha3e3 	:	val_out <= 4'h1d4d;
         4'ha3e8 	:	val_out <= 4'h1d3d;
         4'ha3e9 	:	val_out <= 4'h1d3d;
         4'ha3ea 	:	val_out <= 4'h1d3d;
         4'ha3eb 	:	val_out <= 4'h1d3d;
         4'ha3f0 	:	val_out <= 4'h1d2d;
         4'ha3f1 	:	val_out <= 4'h1d2d;
         4'ha3f2 	:	val_out <= 4'h1d2d;
         4'ha3f3 	:	val_out <= 4'h1d2d;
         4'ha3f8 	:	val_out <= 4'h1d1d;
         4'ha3f9 	:	val_out <= 4'h1d1d;
         4'ha3fa 	:	val_out <= 4'h1d1d;
         4'ha3fb 	:	val_out <= 4'h1d1d;
         4'ha400 	:	val_out <= 4'h1d0d;
         4'ha401 	:	val_out <= 4'h1d0d;
         4'ha402 	:	val_out <= 4'h1d0d;
         4'ha403 	:	val_out <= 4'h1d0d;
         4'ha408 	:	val_out <= 4'h1cfe;
         4'ha409 	:	val_out <= 4'h1cfe;
         4'ha40a 	:	val_out <= 4'h1cfe;
         4'ha40b 	:	val_out <= 4'h1cfe;
         4'ha410 	:	val_out <= 4'h1cee;
         4'ha411 	:	val_out <= 4'h1cee;
         4'ha412 	:	val_out <= 4'h1cee;
         4'ha413 	:	val_out <= 4'h1cee;
         4'ha418 	:	val_out <= 4'h1cde;
         4'ha419 	:	val_out <= 4'h1cde;
         4'ha41a 	:	val_out <= 4'h1cde;
         4'ha41b 	:	val_out <= 4'h1cde;
         4'ha420 	:	val_out <= 4'h1cce;
         4'ha421 	:	val_out <= 4'h1cce;
         4'ha422 	:	val_out <= 4'h1cce;
         4'ha423 	:	val_out <= 4'h1cce;
         4'ha428 	:	val_out <= 4'h1cbe;
         4'ha429 	:	val_out <= 4'h1cbe;
         4'ha42a 	:	val_out <= 4'h1cbe;
         4'ha42b 	:	val_out <= 4'h1cbe;
         4'ha430 	:	val_out <= 4'h1cae;
         4'ha431 	:	val_out <= 4'h1cae;
         4'ha432 	:	val_out <= 4'h1cae;
         4'ha433 	:	val_out <= 4'h1cae;
         4'ha438 	:	val_out <= 4'h1c9e;
         4'ha439 	:	val_out <= 4'h1c9e;
         4'ha43a 	:	val_out <= 4'h1c9e;
         4'ha43b 	:	val_out <= 4'h1c9e;
         4'ha440 	:	val_out <= 4'h1c8e;
         4'ha441 	:	val_out <= 4'h1c8e;
         4'ha442 	:	val_out <= 4'h1c8e;
         4'ha443 	:	val_out <= 4'h1c8e;
         4'ha448 	:	val_out <= 4'h1c7f;
         4'ha449 	:	val_out <= 4'h1c7f;
         4'ha44a 	:	val_out <= 4'h1c7f;
         4'ha44b 	:	val_out <= 4'h1c7f;
         4'ha450 	:	val_out <= 4'h1c6f;
         4'ha451 	:	val_out <= 4'h1c6f;
         4'ha452 	:	val_out <= 4'h1c6f;
         4'ha453 	:	val_out <= 4'h1c6f;
         4'ha458 	:	val_out <= 4'h1c5f;
         4'ha459 	:	val_out <= 4'h1c5f;
         4'ha45a 	:	val_out <= 4'h1c5f;
         4'ha45b 	:	val_out <= 4'h1c5f;
         4'ha460 	:	val_out <= 4'h1c4f;
         4'ha461 	:	val_out <= 4'h1c4f;
         4'ha462 	:	val_out <= 4'h1c4f;
         4'ha463 	:	val_out <= 4'h1c4f;
         4'ha468 	:	val_out <= 4'h1c3f;
         4'ha469 	:	val_out <= 4'h1c3f;
         4'ha46a 	:	val_out <= 4'h1c3f;
         4'ha46b 	:	val_out <= 4'h1c3f;
         4'ha470 	:	val_out <= 4'h1c30;
         4'ha471 	:	val_out <= 4'h1c30;
         4'ha472 	:	val_out <= 4'h1c30;
         4'ha473 	:	val_out <= 4'h1c30;
         4'ha478 	:	val_out <= 4'h1c20;
         4'ha479 	:	val_out <= 4'h1c20;
         4'ha47a 	:	val_out <= 4'h1c20;
         4'ha47b 	:	val_out <= 4'h1c20;
         4'ha480 	:	val_out <= 4'h1c10;
         4'ha481 	:	val_out <= 4'h1c10;
         4'ha482 	:	val_out <= 4'h1c10;
         4'ha483 	:	val_out <= 4'h1c10;
         4'ha488 	:	val_out <= 4'h1c01;
         4'ha489 	:	val_out <= 4'h1c01;
         4'ha48a 	:	val_out <= 4'h1c01;
         4'ha48b 	:	val_out <= 4'h1c01;
         4'ha490 	:	val_out <= 4'h1bf1;
         4'ha491 	:	val_out <= 4'h1bf1;
         4'ha492 	:	val_out <= 4'h1bf1;
         4'ha493 	:	val_out <= 4'h1bf1;
         4'ha498 	:	val_out <= 4'h1be1;
         4'ha499 	:	val_out <= 4'h1be1;
         4'ha49a 	:	val_out <= 4'h1be1;
         4'ha49b 	:	val_out <= 4'h1be1;
         4'ha4a0 	:	val_out <= 4'h1bd2;
         4'ha4a1 	:	val_out <= 4'h1bd2;
         4'ha4a2 	:	val_out <= 4'h1bd2;
         4'ha4a3 	:	val_out <= 4'h1bd2;
         4'ha4a8 	:	val_out <= 4'h1bc2;
         4'ha4a9 	:	val_out <= 4'h1bc2;
         4'ha4aa 	:	val_out <= 4'h1bc2;
         4'ha4ab 	:	val_out <= 4'h1bc2;
         4'ha4b0 	:	val_out <= 4'h1bb2;
         4'ha4b1 	:	val_out <= 4'h1bb2;
         4'ha4b2 	:	val_out <= 4'h1bb2;
         4'ha4b3 	:	val_out <= 4'h1bb2;
         4'ha4b8 	:	val_out <= 4'h1ba3;
         4'ha4b9 	:	val_out <= 4'h1ba3;
         4'ha4ba 	:	val_out <= 4'h1ba3;
         4'ha4bb 	:	val_out <= 4'h1ba3;
         4'ha4c0 	:	val_out <= 4'h1b93;
         4'ha4c1 	:	val_out <= 4'h1b93;
         4'ha4c2 	:	val_out <= 4'h1b93;
         4'ha4c3 	:	val_out <= 4'h1b93;
         4'ha4c8 	:	val_out <= 4'h1b84;
         4'ha4c9 	:	val_out <= 4'h1b84;
         4'ha4ca 	:	val_out <= 4'h1b84;
         4'ha4cb 	:	val_out <= 4'h1b84;
         4'ha4d0 	:	val_out <= 4'h1b74;
         4'ha4d1 	:	val_out <= 4'h1b74;
         4'ha4d2 	:	val_out <= 4'h1b74;
         4'ha4d3 	:	val_out <= 4'h1b74;
         4'ha4d8 	:	val_out <= 4'h1b64;
         4'ha4d9 	:	val_out <= 4'h1b64;
         4'ha4da 	:	val_out <= 4'h1b64;
         4'ha4db 	:	val_out <= 4'h1b64;
         4'ha4e0 	:	val_out <= 4'h1b55;
         4'ha4e1 	:	val_out <= 4'h1b55;
         4'ha4e2 	:	val_out <= 4'h1b55;
         4'ha4e3 	:	val_out <= 4'h1b55;
         4'ha4e8 	:	val_out <= 4'h1b45;
         4'ha4e9 	:	val_out <= 4'h1b45;
         4'ha4ea 	:	val_out <= 4'h1b45;
         4'ha4eb 	:	val_out <= 4'h1b45;
         4'ha4f0 	:	val_out <= 4'h1b36;
         4'ha4f1 	:	val_out <= 4'h1b36;
         4'ha4f2 	:	val_out <= 4'h1b36;
         4'ha4f3 	:	val_out <= 4'h1b36;
         4'ha4f8 	:	val_out <= 4'h1b26;
         4'ha4f9 	:	val_out <= 4'h1b26;
         4'ha4fa 	:	val_out <= 4'h1b26;
         4'ha4fb 	:	val_out <= 4'h1b26;
         4'ha500 	:	val_out <= 4'h1b17;
         4'ha501 	:	val_out <= 4'h1b17;
         4'ha502 	:	val_out <= 4'h1b17;
         4'ha503 	:	val_out <= 4'h1b17;
         4'ha508 	:	val_out <= 4'h1b08;
         4'ha509 	:	val_out <= 4'h1b08;
         4'ha50a 	:	val_out <= 4'h1b08;
         4'ha50b 	:	val_out <= 4'h1b08;
         4'ha510 	:	val_out <= 4'h1af8;
         4'ha511 	:	val_out <= 4'h1af8;
         4'ha512 	:	val_out <= 4'h1af8;
         4'ha513 	:	val_out <= 4'h1af8;
         4'ha518 	:	val_out <= 4'h1ae9;
         4'ha519 	:	val_out <= 4'h1ae9;
         4'ha51a 	:	val_out <= 4'h1ae9;
         4'ha51b 	:	val_out <= 4'h1ae9;
         4'ha520 	:	val_out <= 4'h1ad9;
         4'ha521 	:	val_out <= 4'h1ad9;
         4'ha522 	:	val_out <= 4'h1ad9;
         4'ha523 	:	val_out <= 4'h1ad9;
         4'ha528 	:	val_out <= 4'h1aca;
         4'ha529 	:	val_out <= 4'h1aca;
         4'ha52a 	:	val_out <= 4'h1aca;
         4'ha52b 	:	val_out <= 4'h1aca;
         4'ha530 	:	val_out <= 4'h1aba;
         4'ha531 	:	val_out <= 4'h1aba;
         4'ha532 	:	val_out <= 4'h1aba;
         4'ha533 	:	val_out <= 4'h1aba;
         4'ha538 	:	val_out <= 4'h1aab;
         4'ha539 	:	val_out <= 4'h1aab;
         4'ha53a 	:	val_out <= 4'h1aab;
         4'ha53b 	:	val_out <= 4'h1aab;
         4'ha540 	:	val_out <= 4'h1a9c;
         4'ha541 	:	val_out <= 4'h1a9c;
         4'ha542 	:	val_out <= 4'h1a9c;
         4'ha543 	:	val_out <= 4'h1a9c;
         4'ha548 	:	val_out <= 4'h1a8c;
         4'ha549 	:	val_out <= 4'h1a8c;
         4'ha54a 	:	val_out <= 4'h1a8c;
         4'ha54b 	:	val_out <= 4'h1a8c;
         4'ha550 	:	val_out <= 4'h1a7d;
         4'ha551 	:	val_out <= 4'h1a7d;
         4'ha552 	:	val_out <= 4'h1a7d;
         4'ha553 	:	val_out <= 4'h1a7d;
         4'ha558 	:	val_out <= 4'h1a6e;
         4'ha559 	:	val_out <= 4'h1a6e;
         4'ha55a 	:	val_out <= 4'h1a6e;
         4'ha55b 	:	val_out <= 4'h1a6e;
         4'ha560 	:	val_out <= 4'h1a5f;
         4'ha561 	:	val_out <= 4'h1a5f;
         4'ha562 	:	val_out <= 4'h1a5f;
         4'ha563 	:	val_out <= 4'h1a5f;
         4'ha568 	:	val_out <= 4'h1a4f;
         4'ha569 	:	val_out <= 4'h1a4f;
         4'ha56a 	:	val_out <= 4'h1a4f;
         4'ha56b 	:	val_out <= 4'h1a4f;
         4'ha570 	:	val_out <= 4'h1a40;
         4'ha571 	:	val_out <= 4'h1a40;
         4'ha572 	:	val_out <= 4'h1a40;
         4'ha573 	:	val_out <= 4'h1a40;
         4'ha578 	:	val_out <= 4'h1a31;
         4'ha579 	:	val_out <= 4'h1a31;
         4'ha57a 	:	val_out <= 4'h1a31;
         4'ha57b 	:	val_out <= 4'h1a31;
         4'ha580 	:	val_out <= 4'h1a22;
         4'ha581 	:	val_out <= 4'h1a22;
         4'ha582 	:	val_out <= 4'h1a22;
         4'ha583 	:	val_out <= 4'h1a22;
         4'ha588 	:	val_out <= 4'h1a12;
         4'ha589 	:	val_out <= 4'h1a12;
         4'ha58a 	:	val_out <= 4'h1a12;
         4'ha58b 	:	val_out <= 4'h1a12;
         4'ha590 	:	val_out <= 4'h1a03;
         4'ha591 	:	val_out <= 4'h1a03;
         4'ha592 	:	val_out <= 4'h1a03;
         4'ha593 	:	val_out <= 4'h1a03;
         4'ha598 	:	val_out <= 4'h19f4;
         4'ha599 	:	val_out <= 4'h19f4;
         4'ha59a 	:	val_out <= 4'h19f4;
         4'ha59b 	:	val_out <= 4'h19f4;
         4'ha5a0 	:	val_out <= 4'h19e5;
         4'ha5a1 	:	val_out <= 4'h19e5;
         4'ha5a2 	:	val_out <= 4'h19e5;
         4'ha5a3 	:	val_out <= 4'h19e5;
         4'ha5a8 	:	val_out <= 4'h19d6;
         4'ha5a9 	:	val_out <= 4'h19d6;
         4'ha5aa 	:	val_out <= 4'h19d6;
         4'ha5ab 	:	val_out <= 4'h19d6;
         4'ha5b0 	:	val_out <= 4'h19c6;
         4'ha5b1 	:	val_out <= 4'h19c6;
         4'ha5b2 	:	val_out <= 4'h19c6;
         4'ha5b3 	:	val_out <= 4'h19c6;
         4'ha5b8 	:	val_out <= 4'h19b7;
         4'ha5b9 	:	val_out <= 4'h19b7;
         4'ha5ba 	:	val_out <= 4'h19b7;
         4'ha5bb 	:	val_out <= 4'h19b7;
         4'ha5c0 	:	val_out <= 4'h19a8;
         4'ha5c1 	:	val_out <= 4'h19a8;
         4'ha5c2 	:	val_out <= 4'h19a8;
         4'ha5c3 	:	val_out <= 4'h19a8;
         4'ha5c8 	:	val_out <= 4'h1999;
         4'ha5c9 	:	val_out <= 4'h1999;
         4'ha5ca 	:	val_out <= 4'h1999;
         4'ha5cb 	:	val_out <= 4'h1999;
         4'ha5d0 	:	val_out <= 4'h198a;
         4'ha5d1 	:	val_out <= 4'h198a;
         4'ha5d2 	:	val_out <= 4'h198a;
         4'ha5d3 	:	val_out <= 4'h198a;
         4'ha5d8 	:	val_out <= 4'h197b;
         4'ha5d9 	:	val_out <= 4'h197b;
         4'ha5da 	:	val_out <= 4'h197b;
         4'ha5db 	:	val_out <= 4'h197b;
         4'ha5e0 	:	val_out <= 4'h196c;
         4'ha5e1 	:	val_out <= 4'h196c;
         4'ha5e2 	:	val_out <= 4'h196c;
         4'ha5e3 	:	val_out <= 4'h196c;
         4'ha5e8 	:	val_out <= 4'h195d;
         4'ha5e9 	:	val_out <= 4'h195d;
         4'ha5ea 	:	val_out <= 4'h195d;
         4'ha5eb 	:	val_out <= 4'h195d;
         4'ha5f0 	:	val_out <= 4'h194e;
         4'ha5f1 	:	val_out <= 4'h194e;
         4'ha5f2 	:	val_out <= 4'h194e;
         4'ha5f3 	:	val_out <= 4'h194e;
         4'ha5f8 	:	val_out <= 4'h193f;
         4'ha5f9 	:	val_out <= 4'h193f;
         4'ha5fa 	:	val_out <= 4'h193f;
         4'ha5fb 	:	val_out <= 4'h193f;
         4'ha600 	:	val_out <= 4'h1930;
         4'ha601 	:	val_out <= 4'h1930;
         4'ha602 	:	val_out <= 4'h1930;
         4'ha603 	:	val_out <= 4'h1930;
         4'ha608 	:	val_out <= 4'h1921;
         4'ha609 	:	val_out <= 4'h1921;
         4'ha60a 	:	val_out <= 4'h1921;
         4'ha60b 	:	val_out <= 4'h1921;
         4'ha610 	:	val_out <= 4'h1912;
         4'ha611 	:	val_out <= 4'h1912;
         4'ha612 	:	val_out <= 4'h1912;
         4'ha613 	:	val_out <= 4'h1912;
         4'ha618 	:	val_out <= 4'h1903;
         4'ha619 	:	val_out <= 4'h1903;
         4'ha61a 	:	val_out <= 4'h1903;
         4'ha61b 	:	val_out <= 4'h1903;
         4'ha620 	:	val_out <= 4'h18f4;
         4'ha621 	:	val_out <= 4'h18f4;
         4'ha622 	:	val_out <= 4'h18f4;
         4'ha623 	:	val_out <= 4'h18f4;
         4'ha628 	:	val_out <= 4'h18e5;
         4'ha629 	:	val_out <= 4'h18e5;
         4'ha62a 	:	val_out <= 4'h18e5;
         4'ha62b 	:	val_out <= 4'h18e5;
         4'ha630 	:	val_out <= 4'h18d6;
         4'ha631 	:	val_out <= 4'h18d6;
         4'ha632 	:	val_out <= 4'h18d6;
         4'ha633 	:	val_out <= 4'h18d6;
         4'ha638 	:	val_out <= 4'h18c8;
         4'ha639 	:	val_out <= 4'h18c8;
         4'ha63a 	:	val_out <= 4'h18c8;
         4'ha63b 	:	val_out <= 4'h18c8;
         4'ha640 	:	val_out <= 4'h18b9;
         4'ha641 	:	val_out <= 4'h18b9;
         4'ha642 	:	val_out <= 4'h18b9;
         4'ha643 	:	val_out <= 4'h18b9;
         4'ha648 	:	val_out <= 4'h18aa;
         4'ha649 	:	val_out <= 4'h18aa;
         4'ha64a 	:	val_out <= 4'h18aa;
         4'ha64b 	:	val_out <= 4'h18aa;
         4'ha650 	:	val_out <= 4'h189b;
         4'ha651 	:	val_out <= 4'h189b;
         4'ha652 	:	val_out <= 4'h189b;
         4'ha653 	:	val_out <= 4'h189b;
         4'ha658 	:	val_out <= 4'h188c;
         4'ha659 	:	val_out <= 4'h188c;
         4'ha65a 	:	val_out <= 4'h188c;
         4'ha65b 	:	val_out <= 4'h188c;
         4'ha660 	:	val_out <= 4'h187d;
         4'ha661 	:	val_out <= 4'h187d;
         4'ha662 	:	val_out <= 4'h187d;
         4'ha663 	:	val_out <= 4'h187d;
         4'ha668 	:	val_out <= 4'h186f;
         4'ha669 	:	val_out <= 4'h186f;
         4'ha66a 	:	val_out <= 4'h186f;
         4'ha66b 	:	val_out <= 4'h186f;
         4'ha670 	:	val_out <= 4'h1860;
         4'ha671 	:	val_out <= 4'h1860;
         4'ha672 	:	val_out <= 4'h1860;
         4'ha673 	:	val_out <= 4'h1860;
         4'ha678 	:	val_out <= 4'h1851;
         4'ha679 	:	val_out <= 4'h1851;
         4'ha67a 	:	val_out <= 4'h1851;
         4'ha67b 	:	val_out <= 4'h1851;
         4'ha680 	:	val_out <= 4'h1842;
         4'ha681 	:	val_out <= 4'h1842;
         4'ha682 	:	val_out <= 4'h1842;
         4'ha683 	:	val_out <= 4'h1842;
         4'ha688 	:	val_out <= 4'h1834;
         4'ha689 	:	val_out <= 4'h1834;
         4'ha68a 	:	val_out <= 4'h1834;
         4'ha68b 	:	val_out <= 4'h1834;
         4'ha690 	:	val_out <= 4'h1825;
         4'ha691 	:	val_out <= 4'h1825;
         4'ha692 	:	val_out <= 4'h1825;
         4'ha693 	:	val_out <= 4'h1825;
         4'ha698 	:	val_out <= 4'h1816;
         4'ha699 	:	val_out <= 4'h1816;
         4'ha69a 	:	val_out <= 4'h1816;
         4'ha69b 	:	val_out <= 4'h1816;
         4'ha6a0 	:	val_out <= 4'h1808;
         4'ha6a1 	:	val_out <= 4'h1808;
         4'ha6a2 	:	val_out <= 4'h1808;
         4'ha6a3 	:	val_out <= 4'h1808;
         4'ha6a8 	:	val_out <= 4'h17f9;
         4'ha6a9 	:	val_out <= 4'h17f9;
         4'ha6aa 	:	val_out <= 4'h17f9;
         4'ha6ab 	:	val_out <= 4'h17f9;
         4'ha6b0 	:	val_out <= 4'h17ea;
         4'ha6b1 	:	val_out <= 4'h17ea;
         4'ha6b2 	:	val_out <= 4'h17ea;
         4'ha6b3 	:	val_out <= 4'h17ea;
         4'ha6b8 	:	val_out <= 4'h17dc;
         4'ha6b9 	:	val_out <= 4'h17dc;
         4'ha6ba 	:	val_out <= 4'h17dc;
         4'ha6bb 	:	val_out <= 4'h17dc;
         4'ha6c0 	:	val_out <= 4'h17cd;
         4'ha6c1 	:	val_out <= 4'h17cd;
         4'ha6c2 	:	val_out <= 4'h17cd;
         4'ha6c3 	:	val_out <= 4'h17cd;
         4'ha6c8 	:	val_out <= 4'h17bf;
         4'ha6c9 	:	val_out <= 4'h17bf;
         4'ha6ca 	:	val_out <= 4'h17bf;
         4'ha6cb 	:	val_out <= 4'h17bf;
         4'ha6d0 	:	val_out <= 4'h17b0;
         4'ha6d1 	:	val_out <= 4'h17b0;
         4'ha6d2 	:	val_out <= 4'h17b0;
         4'ha6d3 	:	val_out <= 4'h17b0;
         4'ha6d8 	:	val_out <= 4'h17a1;
         4'ha6d9 	:	val_out <= 4'h17a1;
         4'ha6da 	:	val_out <= 4'h17a1;
         4'ha6db 	:	val_out <= 4'h17a1;
         4'ha6e0 	:	val_out <= 4'h1793;
         4'ha6e1 	:	val_out <= 4'h1793;
         4'ha6e2 	:	val_out <= 4'h1793;
         4'ha6e3 	:	val_out <= 4'h1793;
         4'ha6e8 	:	val_out <= 4'h1784;
         4'ha6e9 	:	val_out <= 4'h1784;
         4'ha6ea 	:	val_out <= 4'h1784;
         4'ha6eb 	:	val_out <= 4'h1784;
         4'ha6f0 	:	val_out <= 4'h1776;
         4'ha6f1 	:	val_out <= 4'h1776;
         4'ha6f2 	:	val_out <= 4'h1776;
         4'ha6f3 	:	val_out <= 4'h1776;
         4'ha6f8 	:	val_out <= 4'h1767;
         4'ha6f9 	:	val_out <= 4'h1767;
         4'ha6fa 	:	val_out <= 4'h1767;
         4'ha6fb 	:	val_out <= 4'h1767;
         4'ha700 	:	val_out <= 4'h1759;
         4'ha701 	:	val_out <= 4'h1759;
         4'ha702 	:	val_out <= 4'h1759;
         4'ha703 	:	val_out <= 4'h1759;
         4'ha708 	:	val_out <= 4'h174a;
         4'ha709 	:	val_out <= 4'h174a;
         4'ha70a 	:	val_out <= 4'h174a;
         4'ha70b 	:	val_out <= 4'h174a;
         4'ha710 	:	val_out <= 4'h173c;
         4'ha711 	:	val_out <= 4'h173c;
         4'ha712 	:	val_out <= 4'h173c;
         4'ha713 	:	val_out <= 4'h173c;
         4'ha718 	:	val_out <= 4'h172e;
         4'ha719 	:	val_out <= 4'h172e;
         4'ha71a 	:	val_out <= 4'h172e;
         4'ha71b 	:	val_out <= 4'h172e;
         4'ha720 	:	val_out <= 4'h171f;
         4'ha721 	:	val_out <= 4'h171f;
         4'ha722 	:	val_out <= 4'h171f;
         4'ha723 	:	val_out <= 4'h171f;
         4'ha728 	:	val_out <= 4'h1711;
         4'ha729 	:	val_out <= 4'h1711;
         4'ha72a 	:	val_out <= 4'h1711;
         4'ha72b 	:	val_out <= 4'h1711;
         4'ha730 	:	val_out <= 4'h1702;
         4'ha731 	:	val_out <= 4'h1702;
         4'ha732 	:	val_out <= 4'h1702;
         4'ha733 	:	val_out <= 4'h1702;
         4'ha738 	:	val_out <= 4'h16f4;
         4'ha739 	:	val_out <= 4'h16f4;
         4'ha73a 	:	val_out <= 4'h16f4;
         4'ha73b 	:	val_out <= 4'h16f4;
         4'ha740 	:	val_out <= 4'h16e6;
         4'ha741 	:	val_out <= 4'h16e6;
         4'ha742 	:	val_out <= 4'h16e6;
         4'ha743 	:	val_out <= 4'h16e6;
         4'ha748 	:	val_out <= 4'h16d7;
         4'ha749 	:	val_out <= 4'h16d7;
         4'ha74a 	:	val_out <= 4'h16d7;
         4'ha74b 	:	val_out <= 4'h16d7;
         4'ha750 	:	val_out <= 4'h16c9;
         4'ha751 	:	val_out <= 4'h16c9;
         4'ha752 	:	val_out <= 4'h16c9;
         4'ha753 	:	val_out <= 4'h16c9;
         4'ha758 	:	val_out <= 4'h16bb;
         4'ha759 	:	val_out <= 4'h16bb;
         4'ha75a 	:	val_out <= 4'h16bb;
         4'ha75b 	:	val_out <= 4'h16bb;
         4'ha760 	:	val_out <= 4'h16ac;
         4'ha761 	:	val_out <= 4'h16ac;
         4'ha762 	:	val_out <= 4'h16ac;
         4'ha763 	:	val_out <= 4'h16ac;
         4'ha768 	:	val_out <= 4'h169e;
         4'ha769 	:	val_out <= 4'h169e;
         4'ha76a 	:	val_out <= 4'h169e;
         4'ha76b 	:	val_out <= 4'h169e;
         4'ha770 	:	val_out <= 4'h1690;
         4'ha771 	:	val_out <= 4'h1690;
         4'ha772 	:	val_out <= 4'h1690;
         4'ha773 	:	val_out <= 4'h1690;
         4'ha778 	:	val_out <= 4'h1682;
         4'ha779 	:	val_out <= 4'h1682;
         4'ha77a 	:	val_out <= 4'h1682;
         4'ha77b 	:	val_out <= 4'h1682;
         4'ha780 	:	val_out <= 4'h1673;
         4'ha781 	:	val_out <= 4'h1673;
         4'ha782 	:	val_out <= 4'h1673;
         4'ha783 	:	val_out <= 4'h1673;
         4'ha788 	:	val_out <= 4'h1665;
         4'ha789 	:	val_out <= 4'h1665;
         4'ha78a 	:	val_out <= 4'h1665;
         4'ha78b 	:	val_out <= 4'h1665;
         4'ha790 	:	val_out <= 4'h1657;
         4'ha791 	:	val_out <= 4'h1657;
         4'ha792 	:	val_out <= 4'h1657;
         4'ha793 	:	val_out <= 4'h1657;
         4'ha798 	:	val_out <= 4'h1649;
         4'ha799 	:	val_out <= 4'h1649;
         4'ha79a 	:	val_out <= 4'h1649;
         4'ha79b 	:	val_out <= 4'h1649;
         4'ha7a0 	:	val_out <= 4'h163b;
         4'ha7a1 	:	val_out <= 4'h163b;
         4'ha7a2 	:	val_out <= 4'h163b;
         4'ha7a3 	:	val_out <= 4'h163b;
         4'ha7a8 	:	val_out <= 4'h162c;
         4'ha7a9 	:	val_out <= 4'h162c;
         4'ha7aa 	:	val_out <= 4'h162c;
         4'ha7ab 	:	val_out <= 4'h162c;
         4'ha7b0 	:	val_out <= 4'h161e;
         4'ha7b1 	:	val_out <= 4'h161e;
         4'ha7b2 	:	val_out <= 4'h161e;
         4'ha7b3 	:	val_out <= 4'h161e;
         4'ha7b8 	:	val_out <= 4'h1610;
         4'ha7b9 	:	val_out <= 4'h1610;
         4'ha7ba 	:	val_out <= 4'h1610;
         4'ha7bb 	:	val_out <= 4'h1610;
         4'ha7c0 	:	val_out <= 4'h1602;
         4'ha7c1 	:	val_out <= 4'h1602;
         4'ha7c2 	:	val_out <= 4'h1602;
         4'ha7c3 	:	val_out <= 4'h1602;
         4'ha7c8 	:	val_out <= 4'h15f4;
         4'ha7c9 	:	val_out <= 4'h15f4;
         4'ha7ca 	:	val_out <= 4'h15f4;
         4'ha7cb 	:	val_out <= 4'h15f4;
         4'ha7d0 	:	val_out <= 4'h15e6;
         4'ha7d1 	:	val_out <= 4'h15e6;
         4'ha7d2 	:	val_out <= 4'h15e6;
         4'ha7d3 	:	val_out <= 4'h15e6;
         4'ha7d8 	:	val_out <= 4'h15d8;
         4'ha7d9 	:	val_out <= 4'h15d8;
         4'ha7da 	:	val_out <= 4'h15d8;
         4'ha7db 	:	val_out <= 4'h15d8;
         4'ha7e0 	:	val_out <= 4'h15ca;
         4'ha7e1 	:	val_out <= 4'h15ca;
         4'ha7e2 	:	val_out <= 4'h15ca;
         4'ha7e3 	:	val_out <= 4'h15ca;
         4'ha7e8 	:	val_out <= 4'h15bc;
         4'ha7e9 	:	val_out <= 4'h15bc;
         4'ha7ea 	:	val_out <= 4'h15bc;
         4'ha7eb 	:	val_out <= 4'h15bc;
         4'ha7f0 	:	val_out <= 4'h15ae;
         4'ha7f1 	:	val_out <= 4'h15ae;
         4'ha7f2 	:	val_out <= 4'h15ae;
         4'ha7f3 	:	val_out <= 4'h15ae;
         4'ha7f8 	:	val_out <= 4'h15a0;
         4'ha7f9 	:	val_out <= 4'h15a0;
         4'ha7fa 	:	val_out <= 4'h15a0;
         4'ha7fb 	:	val_out <= 4'h15a0;
         4'ha800 	:	val_out <= 4'h1592;
         4'ha801 	:	val_out <= 4'h1592;
         4'ha802 	:	val_out <= 4'h1592;
         4'ha803 	:	val_out <= 4'h1592;
         4'ha808 	:	val_out <= 4'h1584;
         4'ha809 	:	val_out <= 4'h1584;
         4'ha80a 	:	val_out <= 4'h1584;
         4'ha80b 	:	val_out <= 4'h1584;
         4'ha810 	:	val_out <= 4'h1576;
         4'ha811 	:	val_out <= 4'h1576;
         4'ha812 	:	val_out <= 4'h1576;
         4'ha813 	:	val_out <= 4'h1576;
         4'ha818 	:	val_out <= 4'h1568;
         4'ha819 	:	val_out <= 4'h1568;
         4'ha81a 	:	val_out <= 4'h1568;
         4'ha81b 	:	val_out <= 4'h1568;
         4'ha820 	:	val_out <= 4'h155a;
         4'ha821 	:	val_out <= 4'h155a;
         4'ha822 	:	val_out <= 4'h155a;
         4'ha823 	:	val_out <= 4'h155a;
         4'ha828 	:	val_out <= 4'h154c;
         4'ha829 	:	val_out <= 4'h154c;
         4'ha82a 	:	val_out <= 4'h154c;
         4'ha82b 	:	val_out <= 4'h154c;
         4'ha830 	:	val_out <= 4'h153e;
         4'ha831 	:	val_out <= 4'h153e;
         4'ha832 	:	val_out <= 4'h153e;
         4'ha833 	:	val_out <= 4'h153e;
         4'ha838 	:	val_out <= 4'h1531;
         4'ha839 	:	val_out <= 4'h1531;
         4'ha83a 	:	val_out <= 4'h1531;
         4'ha83b 	:	val_out <= 4'h1531;
         4'ha840 	:	val_out <= 4'h1523;
         4'ha841 	:	val_out <= 4'h1523;
         4'ha842 	:	val_out <= 4'h1523;
         4'ha843 	:	val_out <= 4'h1523;
         4'ha848 	:	val_out <= 4'h1515;
         4'ha849 	:	val_out <= 4'h1515;
         4'ha84a 	:	val_out <= 4'h1515;
         4'ha84b 	:	val_out <= 4'h1515;
         4'ha850 	:	val_out <= 4'h1507;
         4'ha851 	:	val_out <= 4'h1507;
         4'ha852 	:	val_out <= 4'h1507;
         4'ha853 	:	val_out <= 4'h1507;
         4'ha858 	:	val_out <= 4'h14f9;
         4'ha859 	:	val_out <= 4'h14f9;
         4'ha85a 	:	val_out <= 4'h14f9;
         4'ha85b 	:	val_out <= 4'h14f9;
         4'ha860 	:	val_out <= 4'h14ec;
         4'ha861 	:	val_out <= 4'h14ec;
         4'ha862 	:	val_out <= 4'h14ec;
         4'ha863 	:	val_out <= 4'h14ec;
         4'ha868 	:	val_out <= 4'h14de;
         4'ha869 	:	val_out <= 4'h14de;
         4'ha86a 	:	val_out <= 4'h14de;
         4'ha86b 	:	val_out <= 4'h14de;
         4'ha870 	:	val_out <= 4'h14d0;
         4'ha871 	:	val_out <= 4'h14d0;
         4'ha872 	:	val_out <= 4'h14d0;
         4'ha873 	:	val_out <= 4'h14d0;
         4'ha878 	:	val_out <= 4'h14c2;
         4'ha879 	:	val_out <= 4'h14c2;
         4'ha87a 	:	val_out <= 4'h14c2;
         4'ha87b 	:	val_out <= 4'h14c2;
         4'ha880 	:	val_out <= 4'h14b5;
         4'ha881 	:	val_out <= 4'h14b5;
         4'ha882 	:	val_out <= 4'h14b5;
         4'ha883 	:	val_out <= 4'h14b5;
         4'ha888 	:	val_out <= 4'h14a7;
         4'ha889 	:	val_out <= 4'h14a7;
         4'ha88a 	:	val_out <= 4'h14a7;
         4'ha88b 	:	val_out <= 4'h14a7;
         4'ha890 	:	val_out <= 4'h1499;
         4'ha891 	:	val_out <= 4'h1499;
         4'ha892 	:	val_out <= 4'h1499;
         4'ha893 	:	val_out <= 4'h1499;
         4'ha898 	:	val_out <= 4'h148c;
         4'ha899 	:	val_out <= 4'h148c;
         4'ha89a 	:	val_out <= 4'h148c;
         4'ha89b 	:	val_out <= 4'h148c;
         4'ha8a0 	:	val_out <= 4'h147e;
         4'ha8a1 	:	val_out <= 4'h147e;
         4'ha8a2 	:	val_out <= 4'h147e;
         4'ha8a3 	:	val_out <= 4'h147e;
         4'ha8a8 	:	val_out <= 4'h1470;
         4'ha8a9 	:	val_out <= 4'h1470;
         4'ha8aa 	:	val_out <= 4'h1470;
         4'ha8ab 	:	val_out <= 4'h1470;
         4'ha8b0 	:	val_out <= 4'h1463;
         4'ha8b1 	:	val_out <= 4'h1463;
         4'ha8b2 	:	val_out <= 4'h1463;
         4'ha8b3 	:	val_out <= 4'h1463;
         4'ha8b8 	:	val_out <= 4'h1455;
         4'ha8b9 	:	val_out <= 4'h1455;
         4'ha8ba 	:	val_out <= 4'h1455;
         4'ha8bb 	:	val_out <= 4'h1455;
         4'ha8c0 	:	val_out <= 4'h1447;
         4'ha8c1 	:	val_out <= 4'h1447;
         4'ha8c2 	:	val_out <= 4'h1447;
         4'ha8c3 	:	val_out <= 4'h1447;
         4'ha8c8 	:	val_out <= 4'h143a;
         4'ha8c9 	:	val_out <= 4'h143a;
         4'ha8ca 	:	val_out <= 4'h143a;
         4'ha8cb 	:	val_out <= 4'h143a;
         4'ha8d0 	:	val_out <= 4'h142c;
         4'ha8d1 	:	val_out <= 4'h142c;
         4'ha8d2 	:	val_out <= 4'h142c;
         4'ha8d3 	:	val_out <= 4'h142c;
         4'ha8d8 	:	val_out <= 4'h141f;
         4'ha8d9 	:	val_out <= 4'h141f;
         4'ha8da 	:	val_out <= 4'h141f;
         4'ha8db 	:	val_out <= 4'h141f;
         4'ha8e0 	:	val_out <= 4'h1411;
         4'ha8e1 	:	val_out <= 4'h1411;
         4'ha8e2 	:	val_out <= 4'h1411;
         4'ha8e3 	:	val_out <= 4'h1411;
         4'ha8e8 	:	val_out <= 4'h1404;
         4'ha8e9 	:	val_out <= 4'h1404;
         4'ha8ea 	:	val_out <= 4'h1404;
         4'ha8eb 	:	val_out <= 4'h1404;
         4'ha8f0 	:	val_out <= 4'h13f6;
         4'ha8f1 	:	val_out <= 4'h13f6;
         4'ha8f2 	:	val_out <= 4'h13f6;
         4'ha8f3 	:	val_out <= 4'h13f6;
         4'ha8f8 	:	val_out <= 4'h13e9;
         4'ha8f9 	:	val_out <= 4'h13e9;
         4'ha8fa 	:	val_out <= 4'h13e9;
         4'ha8fb 	:	val_out <= 4'h13e9;
         4'ha900 	:	val_out <= 4'h13db;
         4'ha901 	:	val_out <= 4'h13db;
         4'ha902 	:	val_out <= 4'h13db;
         4'ha903 	:	val_out <= 4'h13db;
         4'ha908 	:	val_out <= 4'h13ce;
         4'ha909 	:	val_out <= 4'h13ce;
         4'ha90a 	:	val_out <= 4'h13ce;
         4'ha90b 	:	val_out <= 4'h13ce;
         4'ha910 	:	val_out <= 4'h13c0;
         4'ha911 	:	val_out <= 4'h13c0;
         4'ha912 	:	val_out <= 4'h13c0;
         4'ha913 	:	val_out <= 4'h13c0;
         4'ha918 	:	val_out <= 4'h13b3;
         4'ha919 	:	val_out <= 4'h13b3;
         4'ha91a 	:	val_out <= 4'h13b3;
         4'ha91b 	:	val_out <= 4'h13b3;
         4'ha920 	:	val_out <= 4'h13a6;
         4'ha921 	:	val_out <= 4'h13a6;
         4'ha922 	:	val_out <= 4'h13a6;
         4'ha923 	:	val_out <= 4'h13a6;
         4'ha928 	:	val_out <= 4'h1398;
         4'ha929 	:	val_out <= 4'h1398;
         4'ha92a 	:	val_out <= 4'h1398;
         4'ha92b 	:	val_out <= 4'h1398;
         4'ha930 	:	val_out <= 4'h138b;
         4'ha931 	:	val_out <= 4'h138b;
         4'ha932 	:	val_out <= 4'h138b;
         4'ha933 	:	val_out <= 4'h138b;
         4'ha938 	:	val_out <= 4'h137e;
         4'ha939 	:	val_out <= 4'h137e;
         4'ha93a 	:	val_out <= 4'h137e;
         4'ha93b 	:	val_out <= 4'h137e;
         4'ha940 	:	val_out <= 4'h1370;
         4'ha941 	:	val_out <= 4'h1370;
         4'ha942 	:	val_out <= 4'h1370;
         4'ha943 	:	val_out <= 4'h1370;
         4'ha948 	:	val_out <= 4'h1363;
         4'ha949 	:	val_out <= 4'h1363;
         4'ha94a 	:	val_out <= 4'h1363;
         4'ha94b 	:	val_out <= 4'h1363;
         4'ha950 	:	val_out <= 4'h1356;
         4'ha951 	:	val_out <= 4'h1356;
         4'ha952 	:	val_out <= 4'h1356;
         4'ha953 	:	val_out <= 4'h1356;
         4'ha958 	:	val_out <= 4'h1348;
         4'ha959 	:	val_out <= 4'h1348;
         4'ha95a 	:	val_out <= 4'h1348;
         4'ha95b 	:	val_out <= 4'h1348;
         4'ha960 	:	val_out <= 4'h133b;
         4'ha961 	:	val_out <= 4'h133b;
         4'ha962 	:	val_out <= 4'h133b;
         4'ha963 	:	val_out <= 4'h133b;
         4'ha968 	:	val_out <= 4'h132e;
         4'ha969 	:	val_out <= 4'h132e;
         4'ha96a 	:	val_out <= 4'h132e;
         4'ha96b 	:	val_out <= 4'h132e;
         4'ha970 	:	val_out <= 4'h1321;
         4'ha971 	:	val_out <= 4'h1321;
         4'ha972 	:	val_out <= 4'h1321;
         4'ha973 	:	val_out <= 4'h1321;
         4'ha978 	:	val_out <= 4'h1313;
         4'ha979 	:	val_out <= 4'h1313;
         4'ha97a 	:	val_out <= 4'h1313;
         4'ha97b 	:	val_out <= 4'h1313;
         4'ha980 	:	val_out <= 4'h1306;
         4'ha981 	:	val_out <= 4'h1306;
         4'ha982 	:	val_out <= 4'h1306;
         4'ha983 	:	val_out <= 4'h1306;
         4'ha988 	:	val_out <= 4'h12f9;
         4'ha989 	:	val_out <= 4'h12f9;
         4'ha98a 	:	val_out <= 4'h12f9;
         4'ha98b 	:	val_out <= 4'h12f9;
         4'ha990 	:	val_out <= 4'h12ec;
         4'ha991 	:	val_out <= 4'h12ec;
         4'ha992 	:	val_out <= 4'h12ec;
         4'ha993 	:	val_out <= 4'h12ec;
         4'ha998 	:	val_out <= 4'h12df;
         4'ha999 	:	val_out <= 4'h12df;
         4'ha99a 	:	val_out <= 4'h12df;
         4'ha99b 	:	val_out <= 4'h12df;
         4'ha9a0 	:	val_out <= 4'h12d2;
         4'ha9a1 	:	val_out <= 4'h12d2;
         4'ha9a2 	:	val_out <= 4'h12d2;
         4'ha9a3 	:	val_out <= 4'h12d2;
         4'ha9a8 	:	val_out <= 4'h12c5;
         4'ha9a9 	:	val_out <= 4'h12c5;
         4'ha9aa 	:	val_out <= 4'h12c5;
         4'ha9ab 	:	val_out <= 4'h12c5;
         4'ha9b0 	:	val_out <= 4'h12b7;
         4'ha9b1 	:	val_out <= 4'h12b7;
         4'ha9b2 	:	val_out <= 4'h12b7;
         4'ha9b3 	:	val_out <= 4'h12b7;
         4'ha9b8 	:	val_out <= 4'h12aa;
         4'ha9b9 	:	val_out <= 4'h12aa;
         4'ha9ba 	:	val_out <= 4'h12aa;
         4'ha9bb 	:	val_out <= 4'h12aa;
         4'ha9c0 	:	val_out <= 4'h129d;
         4'ha9c1 	:	val_out <= 4'h129d;
         4'ha9c2 	:	val_out <= 4'h129d;
         4'ha9c3 	:	val_out <= 4'h129d;
         4'ha9c8 	:	val_out <= 4'h1290;
         4'ha9c9 	:	val_out <= 4'h1290;
         4'ha9ca 	:	val_out <= 4'h1290;
         4'ha9cb 	:	val_out <= 4'h1290;
         4'ha9d0 	:	val_out <= 4'h1283;
         4'ha9d1 	:	val_out <= 4'h1283;
         4'ha9d2 	:	val_out <= 4'h1283;
         4'ha9d3 	:	val_out <= 4'h1283;
         4'ha9d8 	:	val_out <= 4'h1276;
         4'ha9d9 	:	val_out <= 4'h1276;
         4'ha9da 	:	val_out <= 4'h1276;
         4'ha9db 	:	val_out <= 4'h1276;
         4'ha9e0 	:	val_out <= 4'h1269;
         4'ha9e1 	:	val_out <= 4'h1269;
         4'ha9e2 	:	val_out <= 4'h1269;
         4'ha9e3 	:	val_out <= 4'h1269;
         4'ha9e8 	:	val_out <= 4'h125c;
         4'ha9e9 	:	val_out <= 4'h125c;
         4'ha9ea 	:	val_out <= 4'h125c;
         4'ha9eb 	:	val_out <= 4'h125c;
         4'ha9f0 	:	val_out <= 4'h124f;
         4'ha9f1 	:	val_out <= 4'h124f;
         4'ha9f2 	:	val_out <= 4'h124f;
         4'ha9f3 	:	val_out <= 4'h124f;
         4'ha9f8 	:	val_out <= 4'h1242;
         4'ha9f9 	:	val_out <= 4'h1242;
         4'ha9fa 	:	val_out <= 4'h1242;
         4'ha9fb 	:	val_out <= 4'h1242;
         4'haa00 	:	val_out <= 4'h1235;
         4'haa01 	:	val_out <= 4'h1235;
         4'haa02 	:	val_out <= 4'h1235;
         4'haa03 	:	val_out <= 4'h1235;
         4'haa08 	:	val_out <= 4'h1229;
         4'haa09 	:	val_out <= 4'h1229;
         4'haa0a 	:	val_out <= 4'h1229;
         4'haa0b 	:	val_out <= 4'h1229;
         4'haa10 	:	val_out <= 4'h121c;
         4'haa11 	:	val_out <= 4'h121c;
         4'haa12 	:	val_out <= 4'h121c;
         4'haa13 	:	val_out <= 4'h121c;
         4'haa18 	:	val_out <= 4'h120f;
         4'haa19 	:	val_out <= 4'h120f;
         4'haa1a 	:	val_out <= 4'h120f;
         4'haa1b 	:	val_out <= 4'h120f;
         4'haa20 	:	val_out <= 4'h1202;
         4'haa21 	:	val_out <= 4'h1202;
         4'haa22 	:	val_out <= 4'h1202;
         4'haa23 	:	val_out <= 4'h1202;
         4'haa28 	:	val_out <= 4'h11f5;
         4'haa29 	:	val_out <= 4'h11f5;
         4'haa2a 	:	val_out <= 4'h11f5;
         4'haa2b 	:	val_out <= 4'h11f5;
         4'haa30 	:	val_out <= 4'h11e8;
         4'haa31 	:	val_out <= 4'h11e8;
         4'haa32 	:	val_out <= 4'h11e8;
         4'haa33 	:	val_out <= 4'h11e8;
         4'haa38 	:	val_out <= 4'h11db;
         4'haa39 	:	val_out <= 4'h11db;
         4'haa3a 	:	val_out <= 4'h11db;
         4'haa3b 	:	val_out <= 4'h11db;
         4'haa40 	:	val_out <= 4'h11cf;
         4'haa41 	:	val_out <= 4'h11cf;
         4'haa42 	:	val_out <= 4'h11cf;
         4'haa43 	:	val_out <= 4'h11cf;
         4'haa48 	:	val_out <= 4'h11c2;
         4'haa49 	:	val_out <= 4'h11c2;
         4'haa4a 	:	val_out <= 4'h11c2;
         4'haa4b 	:	val_out <= 4'h11c2;
         4'haa50 	:	val_out <= 4'h11b5;
         4'haa51 	:	val_out <= 4'h11b5;
         4'haa52 	:	val_out <= 4'h11b5;
         4'haa53 	:	val_out <= 4'h11b5;
         4'haa58 	:	val_out <= 4'h11a8;
         4'haa59 	:	val_out <= 4'h11a8;
         4'haa5a 	:	val_out <= 4'h11a8;
         4'haa5b 	:	val_out <= 4'h11a8;
         4'haa60 	:	val_out <= 4'h119c;
         4'haa61 	:	val_out <= 4'h119c;
         4'haa62 	:	val_out <= 4'h119c;
         4'haa63 	:	val_out <= 4'h119c;
         4'haa68 	:	val_out <= 4'h118f;
         4'haa69 	:	val_out <= 4'h118f;
         4'haa6a 	:	val_out <= 4'h118f;
         4'haa6b 	:	val_out <= 4'h118f;
         4'haa70 	:	val_out <= 4'h1182;
         4'haa71 	:	val_out <= 4'h1182;
         4'haa72 	:	val_out <= 4'h1182;
         4'haa73 	:	val_out <= 4'h1182;
         4'haa78 	:	val_out <= 4'h1176;
         4'haa79 	:	val_out <= 4'h1176;
         4'haa7a 	:	val_out <= 4'h1176;
         4'haa7b 	:	val_out <= 4'h1176;
         4'haa80 	:	val_out <= 4'h1169;
         4'haa81 	:	val_out <= 4'h1169;
         4'haa82 	:	val_out <= 4'h1169;
         4'haa83 	:	val_out <= 4'h1169;
         4'haa88 	:	val_out <= 4'h115c;
         4'haa89 	:	val_out <= 4'h115c;
         4'haa8a 	:	val_out <= 4'h115c;
         4'haa8b 	:	val_out <= 4'h115c;
         4'haa90 	:	val_out <= 4'h1150;
         4'haa91 	:	val_out <= 4'h1150;
         4'haa92 	:	val_out <= 4'h1150;
         4'haa93 	:	val_out <= 4'h1150;
         4'haa98 	:	val_out <= 4'h1143;
         4'haa99 	:	val_out <= 4'h1143;
         4'haa9a 	:	val_out <= 4'h1143;
         4'haa9b 	:	val_out <= 4'h1143;
         4'haaa0 	:	val_out <= 4'h1136;
         4'haaa1 	:	val_out <= 4'h1136;
         4'haaa2 	:	val_out <= 4'h1136;
         4'haaa3 	:	val_out <= 4'h1136;
         4'haaa8 	:	val_out <= 4'h112a;
         4'haaa9 	:	val_out <= 4'h112a;
         4'haaaa 	:	val_out <= 4'h112a;
         4'haaab 	:	val_out <= 4'h112a;
         4'haab0 	:	val_out <= 4'h111d;
         4'haab1 	:	val_out <= 4'h111d;
         4'haab2 	:	val_out <= 4'h111d;
         4'haab3 	:	val_out <= 4'h111d;
         4'haab8 	:	val_out <= 4'h1111;
         4'haab9 	:	val_out <= 4'h1111;
         4'haaba 	:	val_out <= 4'h1111;
         4'haabb 	:	val_out <= 4'h1111;
         4'haac0 	:	val_out <= 4'h1104;
         4'haac1 	:	val_out <= 4'h1104;
         4'haac2 	:	val_out <= 4'h1104;
         4'haac3 	:	val_out <= 4'h1104;
         4'haac8 	:	val_out <= 4'h10f8;
         4'haac9 	:	val_out <= 4'h10f8;
         4'haaca 	:	val_out <= 4'h10f8;
         4'haacb 	:	val_out <= 4'h10f8;
         4'haad0 	:	val_out <= 4'h10eb;
         4'haad1 	:	val_out <= 4'h10eb;
         4'haad2 	:	val_out <= 4'h10eb;
         4'haad3 	:	val_out <= 4'h10eb;
         4'haad8 	:	val_out <= 4'h10df;
         4'haad9 	:	val_out <= 4'h10df;
         4'haada 	:	val_out <= 4'h10df;
         4'haadb 	:	val_out <= 4'h10df;
         4'haae0 	:	val_out <= 4'h10d2;
         4'haae1 	:	val_out <= 4'h10d2;
         4'haae2 	:	val_out <= 4'h10d2;
         4'haae3 	:	val_out <= 4'h10d2;
         4'haae8 	:	val_out <= 4'h10c6;
         4'haae9 	:	val_out <= 4'h10c6;
         4'haaea 	:	val_out <= 4'h10c6;
         4'haaeb 	:	val_out <= 4'h10c6;
         4'haaf0 	:	val_out <= 4'h10b9;
         4'haaf1 	:	val_out <= 4'h10b9;
         4'haaf2 	:	val_out <= 4'h10b9;
         4'haaf3 	:	val_out <= 4'h10b9;
         4'haaf8 	:	val_out <= 4'h10ad;
         4'haaf9 	:	val_out <= 4'h10ad;
         4'haafa 	:	val_out <= 4'h10ad;
         4'haafb 	:	val_out <= 4'h10ad;
         4'hab00 	:	val_out <= 4'h10a0;
         4'hab01 	:	val_out <= 4'h10a0;
         4'hab02 	:	val_out <= 4'h10a0;
         4'hab03 	:	val_out <= 4'h10a0;
         4'hab08 	:	val_out <= 4'h1094;
         4'hab09 	:	val_out <= 4'h1094;
         4'hab0a 	:	val_out <= 4'h1094;
         4'hab0b 	:	val_out <= 4'h1094;
         4'hab10 	:	val_out <= 4'h1088;
         4'hab11 	:	val_out <= 4'h1088;
         4'hab12 	:	val_out <= 4'h1088;
         4'hab13 	:	val_out <= 4'h1088;
         4'hab18 	:	val_out <= 4'h107b;
         4'hab19 	:	val_out <= 4'h107b;
         4'hab1a 	:	val_out <= 4'h107b;
         4'hab1b 	:	val_out <= 4'h107b;
         4'hab20 	:	val_out <= 4'h106f;
         4'hab21 	:	val_out <= 4'h106f;
         4'hab22 	:	val_out <= 4'h106f;
         4'hab23 	:	val_out <= 4'h106f;
         4'hab28 	:	val_out <= 4'h1063;
         4'hab29 	:	val_out <= 4'h1063;
         4'hab2a 	:	val_out <= 4'h1063;
         4'hab2b 	:	val_out <= 4'h1063;
         4'hab30 	:	val_out <= 4'h1056;
         4'hab31 	:	val_out <= 4'h1056;
         4'hab32 	:	val_out <= 4'h1056;
         4'hab33 	:	val_out <= 4'h1056;
         4'hab38 	:	val_out <= 4'h104a;
         4'hab39 	:	val_out <= 4'h104a;
         4'hab3a 	:	val_out <= 4'h104a;
         4'hab3b 	:	val_out <= 4'h104a;
         4'hab40 	:	val_out <= 4'h103e;
         4'hab41 	:	val_out <= 4'h103e;
         4'hab42 	:	val_out <= 4'h103e;
         4'hab43 	:	val_out <= 4'h103e;
         4'hab48 	:	val_out <= 4'h1032;
         4'hab49 	:	val_out <= 4'h1032;
         4'hab4a 	:	val_out <= 4'h1032;
         4'hab4b 	:	val_out <= 4'h1032;
         4'hab50 	:	val_out <= 4'h1025;
         4'hab51 	:	val_out <= 4'h1025;
         4'hab52 	:	val_out <= 4'h1025;
         4'hab53 	:	val_out <= 4'h1025;
         4'hab58 	:	val_out <= 4'h1019;
         4'hab59 	:	val_out <= 4'h1019;
         4'hab5a 	:	val_out <= 4'h1019;
         4'hab5b 	:	val_out <= 4'h1019;
         4'hab60 	:	val_out <= 4'h100d;
         4'hab61 	:	val_out <= 4'h100d;
         4'hab62 	:	val_out <= 4'h100d;
         4'hab63 	:	val_out <= 4'h100d;
         4'hab68 	:	val_out <= 4'h1001;
         4'hab69 	:	val_out <= 4'h1001;
         4'hab6a 	:	val_out <= 4'h1001;
         4'hab6b 	:	val_out <= 4'h1001;
         4'hab70 	:	val_out <= 4'h0ff5;
         4'hab71 	:	val_out <= 4'h0ff5;
         4'hab72 	:	val_out <= 4'h0ff5;
         4'hab73 	:	val_out <= 4'h0ff5;
         4'hab78 	:	val_out <= 4'h0fe9;
         4'hab79 	:	val_out <= 4'h0fe9;
         4'hab7a 	:	val_out <= 4'h0fe9;
         4'hab7b 	:	val_out <= 4'h0fe9;
         4'hab80 	:	val_out <= 4'h0fdc;
         4'hab81 	:	val_out <= 4'h0fdc;
         4'hab82 	:	val_out <= 4'h0fdc;
         4'hab83 	:	val_out <= 4'h0fdc;
         4'hab88 	:	val_out <= 4'h0fd0;
         4'hab89 	:	val_out <= 4'h0fd0;
         4'hab8a 	:	val_out <= 4'h0fd0;
         4'hab8b 	:	val_out <= 4'h0fd0;
         4'hab90 	:	val_out <= 4'h0fc4;
         4'hab91 	:	val_out <= 4'h0fc4;
         4'hab92 	:	val_out <= 4'h0fc4;
         4'hab93 	:	val_out <= 4'h0fc4;
         4'hab98 	:	val_out <= 4'h0fb8;
         4'hab99 	:	val_out <= 4'h0fb8;
         4'hab9a 	:	val_out <= 4'h0fb8;
         4'hab9b 	:	val_out <= 4'h0fb8;
         4'haba0 	:	val_out <= 4'h0fac;
         4'haba1 	:	val_out <= 4'h0fac;
         4'haba2 	:	val_out <= 4'h0fac;
         4'haba3 	:	val_out <= 4'h0fac;
         4'haba8 	:	val_out <= 4'h0fa0;
         4'haba9 	:	val_out <= 4'h0fa0;
         4'habaa 	:	val_out <= 4'h0fa0;
         4'habab 	:	val_out <= 4'h0fa0;
         4'habb0 	:	val_out <= 4'h0f94;
         4'habb1 	:	val_out <= 4'h0f94;
         4'habb2 	:	val_out <= 4'h0f94;
         4'habb3 	:	val_out <= 4'h0f94;
         4'habb8 	:	val_out <= 4'h0f88;
         4'habb9 	:	val_out <= 4'h0f88;
         4'habba 	:	val_out <= 4'h0f88;
         4'habbb 	:	val_out <= 4'h0f88;
         4'habc0 	:	val_out <= 4'h0f7c;
         4'habc1 	:	val_out <= 4'h0f7c;
         4'habc2 	:	val_out <= 4'h0f7c;
         4'habc3 	:	val_out <= 4'h0f7c;
         4'habc8 	:	val_out <= 4'h0f70;
         4'habc9 	:	val_out <= 4'h0f70;
         4'habca 	:	val_out <= 4'h0f70;
         4'habcb 	:	val_out <= 4'h0f70;
         4'habd0 	:	val_out <= 4'h0f64;
         4'habd1 	:	val_out <= 4'h0f64;
         4'habd2 	:	val_out <= 4'h0f64;
         4'habd3 	:	val_out <= 4'h0f64;
         4'habd8 	:	val_out <= 4'h0f58;
         4'habd9 	:	val_out <= 4'h0f58;
         4'habda 	:	val_out <= 4'h0f58;
         4'habdb 	:	val_out <= 4'h0f58;
         4'habe0 	:	val_out <= 4'h0f4c;
         4'habe1 	:	val_out <= 4'h0f4c;
         4'habe2 	:	val_out <= 4'h0f4c;
         4'habe3 	:	val_out <= 4'h0f4c;
         4'habe8 	:	val_out <= 4'h0f40;
         4'habe9 	:	val_out <= 4'h0f40;
         4'habea 	:	val_out <= 4'h0f40;
         4'habeb 	:	val_out <= 4'h0f40;
         4'habf0 	:	val_out <= 4'h0f34;
         4'habf1 	:	val_out <= 4'h0f34;
         4'habf2 	:	val_out <= 4'h0f34;
         4'habf3 	:	val_out <= 4'h0f34;
         4'habf8 	:	val_out <= 4'h0f29;
         4'habf9 	:	val_out <= 4'h0f29;
         4'habfa 	:	val_out <= 4'h0f29;
         4'habfb 	:	val_out <= 4'h0f29;
         4'hac00 	:	val_out <= 4'h0f1d;
         4'hac01 	:	val_out <= 4'h0f1d;
         4'hac02 	:	val_out <= 4'h0f1d;
         4'hac03 	:	val_out <= 4'h0f1d;
         4'hac08 	:	val_out <= 4'h0f11;
         4'hac09 	:	val_out <= 4'h0f11;
         4'hac0a 	:	val_out <= 4'h0f11;
         4'hac0b 	:	val_out <= 4'h0f11;
         4'hac10 	:	val_out <= 4'h0f05;
         4'hac11 	:	val_out <= 4'h0f05;
         4'hac12 	:	val_out <= 4'h0f05;
         4'hac13 	:	val_out <= 4'h0f05;
         4'hac18 	:	val_out <= 4'h0ef9;
         4'hac19 	:	val_out <= 4'h0ef9;
         4'hac1a 	:	val_out <= 4'h0ef9;
         4'hac1b 	:	val_out <= 4'h0ef9;
         4'hac20 	:	val_out <= 4'h0eed;
         4'hac21 	:	val_out <= 4'h0eed;
         4'hac22 	:	val_out <= 4'h0eed;
         4'hac23 	:	val_out <= 4'h0eed;
         4'hac28 	:	val_out <= 4'h0ee2;
         4'hac29 	:	val_out <= 4'h0ee2;
         4'hac2a 	:	val_out <= 4'h0ee2;
         4'hac2b 	:	val_out <= 4'h0ee2;
         4'hac30 	:	val_out <= 4'h0ed6;
         4'hac31 	:	val_out <= 4'h0ed6;
         4'hac32 	:	val_out <= 4'h0ed6;
         4'hac33 	:	val_out <= 4'h0ed6;
         4'hac38 	:	val_out <= 4'h0eca;
         4'hac39 	:	val_out <= 4'h0eca;
         4'hac3a 	:	val_out <= 4'h0eca;
         4'hac3b 	:	val_out <= 4'h0eca;
         4'hac40 	:	val_out <= 4'h0ebe;
         4'hac41 	:	val_out <= 4'h0ebe;
         4'hac42 	:	val_out <= 4'h0ebe;
         4'hac43 	:	val_out <= 4'h0ebe;
         4'hac48 	:	val_out <= 4'h0eb3;
         4'hac49 	:	val_out <= 4'h0eb3;
         4'hac4a 	:	val_out <= 4'h0eb3;
         4'hac4b 	:	val_out <= 4'h0eb3;
         4'hac50 	:	val_out <= 4'h0ea7;
         4'hac51 	:	val_out <= 4'h0ea7;
         4'hac52 	:	val_out <= 4'h0ea7;
         4'hac53 	:	val_out <= 4'h0ea7;
         4'hac58 	:	val_out <= 4'h0e9b;
         4'hac59 	:	val_out <= 4'h0e9b;
         4'hac5a 	:	val_out <= 4'h0e9b;
         4'hac5b 	:	val_out <= 4'h0e9b;
         4'hac60 	:	val_out <= 4'h0e90;
         4'hac61 	:	val_out <= 4'h0e90;
         4'hac62 	:	val_out <= 4'h0e90;
         4'hac63 	:	val_out <= 4'h0e90;
         4'hac68 	:	val_out <= 4'h0e84;
         4'hac69 	:	val_out <= 4'h0e84;
         4'hac6a 	:	val_out <= 4'h0e84;
         4'hac6b 	:	val_out <= 4'h0e84;
         4'hac70 	:	val_out <= 4'h0e79;
         4'hac71 	:	val_out <= 4'h0e79;
         4'hac72 	:	val_out <= 4'h0e79;
         4'hac73 	:	val_out <= 4'h0e79;
         4'hac78 	:	val_out <= 4'h0e6d;
         4'hac79 	:	val_out <= 4'h0e6d;
         4'hac7a 	:	val_out <= 4'h0e6d;
         4'hac7b 	:	val_out <= 4'h0e6d;
         4'hac80 	:	val_out <= 4'h0e61;
         4'hac81 	:	val_out <= 4'h0e61;
         4'hac82 	:	val_out <= 4'h0e61;
         4'hac83 	:	val_out <= 4'h0e61;
         4'hac88 	:	val_out <= 4'h0e56;
         4'hac89 	:	val_out <= 4'h0e56;
         4'hac8a 	:	val_out <= 4'h0e56;
         4'hac8b 	:	val_out <= 4'h0e56;
         4'hac90 	:	val_out <= 4'h0e4a;
         4'hac91 	:	val_out <= 4'h0e4a;
         4'hac92 	:	val_out <= 4'h0e4a;
         4'hac93 	:	val_out <= 4'h0e4a;
         4'hac98 	:	val_out <= 4'h0e3f;
         4'hac99 	:	val_out <= 4'h0e3f;
         4'hac9a 	:	val_out <= 4'h0e3f;
         4'hac9b 	:	val_out <= 4'h0e3f;
         4'haca0 	:	val_out <= 4'h0e33;
         4'haca1 	:	val_out <= 4'h0e33;
         4'haca2 	:	val_out <= 4'h0e33;
         4'haca3 	:	val_out <= 4'h0e33;
         4'haca8 	:	val_out <= 4'h0e28;
         4'haca9 	:	val_out <= 4'h0e28;
         4'hacaa 	:	val_out <= 4'h0e28;
         4'hacab 	:	val_out <= 4'h0e28;
         4'hacb0 	:	val_out <= 4'h0e1c;
         4'hacb1 	:	val_out <= 4'h0e1c;
         4'hacb2 	:	val_out <= 4'h0e1c;
         4'hacb3 	:	val_out <= 4'h0e1c;
         4'hacb8 	:	val_out <= 4'h0e11;
         4'hacb9 	:	val_out <= 4'h0e11;
         4'hacba 	:	val_out <= 4'h0e11;
         4'hacbb 	:	val_out <= 4'h0e11;
         4'hacc0 	:	val_out <= 4'h0e05;
         4'hacc1 	:	val_out <= 4'h0e05;
         4'hacc2 	:	val_out <= 4'h0e05;
         4'hacc3 	:	val_out <= 4'h0e05;
         4'hacc8 	:	val_out <= 4'h0dfa;
         4'hacc9 	:	val_out <= 4'h0dfa;
         4'hacca 	:	val_out <= 4'h0dfa;
         4'haccb 	:	val_out <= 4'h0dfa;
         4'hacd0 	:	val_out <= 4'h0dee;
         4'hacd1 	:	val_out <= 4'h0dee;
         4'hacd2 	:	val_out <= 4'h0dee;
         4'hacd3 	:	val_out <= 4'h0dee;
         4'hacd8 	:	val_out <= 4'h0de3;
         4'hacd9 	:	val_out <= 4'h0de3;
         4'hacda 	:	val_out <= 4'h0de3;
         4'hacdb 	:	val_out <= 4'h0de3;
         4'hace0 	:	val_out <= 4'h0dd8;
         4'hace1 	:	val_out <= 4'h0dd8;
         4'hace2 	:	val_out <= 4'h0dd8;
         4'hace3 	:	val_out <= 4'h0dd8;
         4'hace8 	:	val_out <= 4'h0dcc;
         4'hace9 	:	val_out <= 4'h0dcc;
         4'hacea 	:	val_out <= 4'h0dcc;
         4'haceb 	:	val_out <= 4'h0dcc;
         4'hacf0 	:	val_out <= 4'h0dc1;
         4'hacf1 	:	val_out <= 4'h0dc1;
         4'hacf2 	:	val_out <= 4'h0dc1;
         4'hacf3 	:	val_out <= 4'h0dc1;
         4'hacf8 	:	val_out <= 4'h0db6;
         4'hacf9 	:	val_out <= 4'h0db6;
         4'hacfa 	:	val_out <= 4'h0db6;
         4'hacfb 	:	val_out <= 4'h0db6;
         4'had00 	:	val_out <= 4'h0daa;
         4'had01 	:	val_out <= 4'h0daa;
         4'had02 	:	val_out <= 4'h0daa;
         4'had03 	:	val_out <= 4'h0daa;
         4'had08 	:	val_out <= 4'h0d9f;
         4'had09 	:	val_out <= 4'h0d9f;
         4'had0a 	:	val_out <= 4'h0d9f;
         4'had0b 	:	val_out <= 4'h0d9f;
         4'had10 	:	val_out <= 4'h0d94;
         4'had11 	:	val_out <= 4'h0d94;
         4'had12 	:	val_out <= 4'h0d94;
         4'had13 	:	val_out <= 4'h0d94;
         4'had18 	:	val_out <= 4'h0d89;
         4'had19 	:	val_out <= 4'h0d89;
         4'had1a 	:	val_out <= 4'h0d89;
         4'had1b 	:	val_out <= 4'h0d89;
         4'had20 	:	val_out <= 4'h0d7d;
         4'had21 	:	val_out <= 4'h0d7d;
         4'had22 	:	val_out <= 4'h0d7d;
         4'had23 	:	val_out <= 4'h0d7d;
         4'had28 	:	val_out <= 4'h0d72;
         4'had29 	:	val_out <= 4'h0d72;
         4'had2a 	:	val_out <= 4'h0d72;
         4'had2b 	:	val_out <= 4'h0d72;
         4'had30 	:	val_out <= 4'h0d67;
         4'had31 	:	val_out <= 4'h0d67;
         4'had32 	:	val_out <= 4'h0d67;
         4'had33 	:	val_out <= 4'h0d67;
         4'had38 	:	val_out <= 4'h0d5c;
         4'had39 	:	val_out <= 4'h0d5c;
         4'had3a 	:	val_out <= 4'h0d5c;
         4'had3b 	:	val_out <= 4'h0d5c;
         4'had40 	:	val_out <= 4'h0d50;
         4'had41 	:	val_out <= 4'h0d50;
         4'had42 	:	val_out <= 4'h0d50;
         4'had43 	:	val_out <= 4'h0d50;
         4'had48 	:	val_out <= 4'h0d45;
         4'had49 	:	val_out <= 4'h0d45;
         4'had4a 	:	val_out <= 4'h0d45;
         4'had4b 	:	val_out <= 4'h0d45;
         4'had50 	:	val_out <= 4'h0d3a;
         4'had51 	:	val_out <= 4'h0d3a;
         4'had52 	:	val_out <= 4'h0d3a;
         4'had53 	:	val_out <= 4'h0d3a;
         4'had58 	:	val_out <= 4'h0d2f;
         4'had59 	:	val_out <= 4'h0d2f;
         4'had5a 	:	val_out <= 4'h0d2f;
         4'had5b 	:	val_out <= 4'h0d2f;
         4'had60 	:	val_out <= 4'h0d24;
         4'had61 	:	val_out <= 4'h0d24;
         4'had62 	:	val_out <= 4'h0d24;
         4'had63 	:	val_out <= 4'h0d24;
         4'had68 	:	val_out <= 4'h0d19;
         4'had69 	:	val_out <= 4'h0d19;
         4'had6a 	:	val_out <= 4'h0d19;
         4'had6b 	:	val_out <= 4'h0d19;
         4'had70 	:	val_out <= 4'h0d0e;
         4'had71 	:	val_out <= 4'h0d0e;
         4'had72 	:	val_out <= 4'h0d0e;
         4'had73 	:	val_out <= 4'h0d0e;
         4'had78 	:	val_out <= 4'h0d03;
         4'had79 	:	val_out <= 4'h0d03;
         4'had7a 	:	val_out <= 4'h0d03;
         4'had7b 	:	val_out <= 4'h0d03;
         4'had80 	:	val_out <= 4'h0cf8;
         4'had81 	:	val_out <= 4'h0cf8;
         4'had82 	:	val_out <= 4'h0cf8;
         4'had83 	:	val_out <= 4'h0cf8;
         4'had88 	:	val_out <= 4'h0ced;
         4'had89 	:	val_out <= 4'h0ced;
         4'had8a 	:	val_out <= 4'h0ced;
         4'had8b 	:	val_out <= 4'h0ced;
         4'had90 	:	val_out <= 4'h0ce2;
         4'had91 	:	val_out <= 4'h0ce2;
         4'had92 	:	val_out <= 4'h0ce2;
         4'had93 	:	val_out <= 4'h0ce2;
         4'had98 	:	val_out <= 4'h0cd7;
         4'had99 	:	val_out <= 4'h0cd7;
         4'had9a 	:	val_out <= 4'h0cd7;
         4'had9b 	:	val_out <= 4'h0cd7;
         4'hada0 	:	val_out <= 4'h0ccc;
         4'hada1 	:	val_out <= 4'h0ccc;
         4'hada2 	:	val_out <= 4'h0ccc;
         4'hada3 	:	val_out <= 4'h0ccc;
         4'hada8 	:	val_out <= 4'h0cc1;
         4'hada9 	:	val_out <= 4'h0cc1;
         4'hadaa 	:	val_out <= 4'h0cc1;
         4'hadab 	:	val_out <= 4'h0cc1;
         4'hadb0 	:	val_out <= 4'h0cb6;
         4'hadb1 	:	val_out <= 4'h0cb6;
         4'hadb2 	:	val_out <= 4'h0cb6;
         4'hadb3 	:	val_out <= 4'h0cb6;
         4'hadb8 	:	val_out <= 4'h0cab;
         4'hadb9 	:	val_out <= 4'h0cab;
         4'hadba 	:	val_out <= 4'h0cab;
         4'hadbb 	:	val_out <= 4'h0cab;
         4'hadc0 	:	val_out <= 4'h0ca0;
         4'hadc1 	:	val_out <= 4'h0ca0;
         4'hadc2 	:	val_out <= 4'h0ca0;
         4'hadc3 	:	val_out <= 4'h0ca0;
         4'hadc8 	:	val_out <= 4'h0c95;
         4'hadc9 	:	val_out <= 4'h0c95;
         4'hadca 	:	val_out <= 4'h0c95;
         4'hadcb 	:	val_out <= 4'h0c95;
         4'hadd0 	:	val_out <= 4'h0c8a;
         4'hadd1 	:	val_out <= 4'h0c8a;
         4'hadd2 	:	val_out <= 4'h0c8a;
         4'hadd3 	:	val_out <= 4'h0c8a;
         4'hadd8 	:	val_out <= 4'h0c80;
         4'hadd9 	:	val_out <= 4'h0c80;
         4'hadda 	:	val_out <= 4'h0c80;
         4'haddb 	:	val_out <= 4'h0c80;
         4'hade0 	:	val_out <= 4'h0c75;
         4'hade1 	:	val_out <= 4'h0c75;
         4'hade2 	:	val_out <= 4'h0c75;
         4'hade3 	:	val_out <= 4'h0c75;
         4'hade8 	:	val_out <= 4'h0c6a;
         4'hade9 	:	val_out <= 4'h0c6a;
         4'hadea 	:	val_out <= 4'h0c6a;
         4'hadeb 	:	val_out <= 4'h0c6a;
         4'hadf0 	:	val_out <= 4'h0c5f;
         4'hadf1 	:	val_out <= 4'h0c5f;
         4'hadf2 	:	val_out <= 4'h0c5f;
         4'hadf3 	:	val_out <= 4'h0c5f;
         4'hadf8 	:	val_out <= 4'h0c54;
         4'hadf9 	:	val_out <= 4'h0c54;
         4'hadfa 	:	val_out <= 4'h0c54;
         4'hadfb 	:	val_out <= 4'h0c54;
         4'hae00 	:	val_out <= 4'h0c4a;
         4'hae01 	:	val_out <= 4'h0c4a;
         4'hae02 	:	val_out <= 4'h0c4a;
         4'hae03 	:	val_out <= 4'h0c4a;
         4'hae08 	:	val_out <= 4'h0c3f;
         4'hae09 	:	val_out <= 4'h0c3f;
         4'hae0a 	:	val_out <= 4'h0c3f;
         4'hae0b 	:	val_out <= 4'h0c3f;
         4'hae10 	:	val_out <= 4'h0c34;
         4'hae11 	:	val_out <= 4'h0c34;
         4'hae12 	:	val_out <= 4'h0c34;
         4'hae13 	:	val_out <= 4'h0c34;
         4'hae18 	:	val_out <= 4'h0c29;
         4'hae19 	:	val_out <= 4'h0c29;
         4'hae1a 	:	val_out <= 4'h0c29;
         4'hae1b 	:	val_out <= 4'h0c29;
         4'hae20 	:	val_out <= 4'h0c1f;
         4'hae21 	:	val_out <= 4'h0c1f;
         4'hae22 	:	val_out <= 4'h0c1f;
         4'hae23 	:	val_out <= 4'h0c1f;
         4'hae28 	:	val_out <= 4'h0c14;
         4'hae29 	:	val_out <= 4'h0c14;
         4'hae2a 	:	val_out <= 4'h0c14;
         4'hae2b 	:	val_out <= 4'h0c14;
         4'hae30 	:	val_out <= 4'h0c09;
         4'hae31 	:	val_out <= 4'h0c09;
         4'hae32 	:	val_out <= 4'h0c09;
         4'hae33 	:	val_out <= 4'h0c09;
         4'hae38 	:	val_out <= 4'h0bff;
         4'hae39 	:	val_out <= 4'h0bff;
         4'hae3a 	:	val_out <= 4'h0bff;
         4'hae3b 	:	val_out <= 4'h0bff;
         4'hae40 	:	val_out <= 4'h0bf4;
         4'hae41 	:	val_out <= 4'h0bf4;
         4'hae42 	:	val_out <= 4'h0bf4;
         4'hae43 	:	val_out <= 4'h0bf4;
         4'hae48 	:	val_out <= 4'h0bea;
         4'hae49 	:	val_out <= 4'h0bea;
         4'hae4a 	:	val_out <= 4'h0bea;
         4'hae4b 	:	val_out <= 4'h0bea;
         4'hae50 	:	val_out <= 4'h0bdf;
         4'hae51 	:	val_out <= 4'h0bdf;
         4'hae52 	:	val_out <= 4'h0bdf;
         4'hae53 	:	val_out <= 4'h0bdf;
         4'hae58 	:	val_out <= 4'h0bd4;
         4'hae59 	:	val_out <= 4'h0bd4;
         4'hae5a 	:	val_out <= 4'h0bd4;
         4'hae5b 	:	val_out <= 4'h0bd4;
         4'hae60 	:	val_out <= 4'h0bca;
         4'hae61 	:	val_out <= 4'h0bca;
         4'hae62 	:	val_out <= 4'h0bca;
         4'hae63 	:	val_out <= 4'h0bca;
         4'hae68 	:	val_out <= 4'h0bbf;
         4'hae69 	:	val_out <= 4'h0bbf;
         4'hae6a 	:	val_out <= 4'h0bbf;
         4'hae6b 	:	val_out <= 4'h0bbf;
         4'hae70 	:	val_out <= 4'h0bb5;
         4'hae71 	:	val_out <= 4'h0bb5;
         4'hae72 	:	val_out <= 4'h0bb5;
         4'hae73 	:	val_out <= 4'h0bb5;
         4'hae78 	:	val_out <= 4'h0baa;
         4'hae79 	:	val_out <= 4'h0baa;
         4'hae7a 	:	val_out <= 4'h0baa;
         4'hae7b 	:	val_out <= 4'h0baa;
         4'hae80 	:	val_out <= 4'h0ba0;
         4'hae81 	:	val_out <= 4'h0ba0;
         4'hae82 	:	val_out <= 4'h0ba0;
         4'hae83 	:	val_out <= 4'h0ba0;
         4'hae88 	:	val_out <= 4'h0b95;
         4'hae89 	:	val_out <= 4'h0b95;
         4'hae8a 	:	val_out <= 4'h0b95;
         4'hae8b 	:	val_out <= 4'h0b95;
         4'hae90 	:	val_out <= 4'h0b8b;
         4'hae91 	:	val_out <= 4'h0b8b;
         4'hae92 	:	val_out <= 4'h0b8b;
         4'hae93 	:	val_out <= 4'h0b8b;
         4'hae98 	:	val_out <= 4'h0b81;
         4'hae99 	:	val_out <= 4'h0b81;
         4'hae9a 	:	val_out <= 4'h0b81;
         4'hae9b 	:	val_out <= 4'h0b81;
         4'haea0 	:	val_out <= 4'h0b76;
         4'haea1 	:	val_out <= 4'h0b76;
         4'haea2 	:	val_out <= 4'h0b76;
         4'haea3 	:	val_out <= 4'h0b76;
         4'haea8 	:	val_out <= 4'h0b6c;
         4'haea9 	:	val_out <= 4'h0b6c;
         4'haeaa 	:	val_out <= 4'h0b6c;
         4'haeab 	:	val_out <= 4'h0b6c;
         4'haeb0 	:	val_out <= 4'h0b61;
         4'haeb1 	:	val_out <= 4'h0b61;
         4'haeb2 	:	val_out <= 4'h0b61;
         4'haeb3 	:	val_out <= 4'h0b61;
         4'haeb8 	:	val_out <= 4'h0b57;
         4'haeb9 	:	val_out <= 4'h0b57;
         4'haeba 	:	val_out <= 4'h0b57;
         4'haebb 	:	val_out <= 4'h0b57;
         4'haec0 	:	val_out <= 4'h0b4d;
         4'haec1 	:	val_out <= 4'h0b4d;
         4'haec2 	:	val_out <= 4'h0b4d;
         4'haec3 	:	val_out <= 4'h0b4d;
         4'haec8 	:	val_out <= 4'h0b42;
         4'haec9 	:	val_out <= 4'h0b42;
         4'haeca 	:	val_out <= 4'h0b42;
         4'haecb 	:	val_out <= 4'h0b42;
         4'haed0 	:	val_out <= 4'h0b38;
         4'haed1 	:	val_out <= 4'h0b38;
         4'haed2 	:	val_out <= 4'h0b38;
         4'haed3 	:	val_out <= 4'h0b38;
         4'haed8 	:	val_out <= 4'h0b2e;
         4'haed9 	:	val_out <= 4'h0b2e;
         4'haeda 	:	val_out <= 4'h0b2e;
         4'haedb 	:	val_out <= 4'h0b2e;
         4'haee0 	:	val_out <= 4'h0b24;
         4'haee1 	:	val_out <= 4'h0b24;
         4'haee2 	:	val_out <= 4'h0b24;
         4'haee3 	:	val_out <= 4'h0b24;
         4'haee8 	:	val_out <= 4'h0b19;
         4'haee9 	:	val_out <= 4'h0b19;
         4'haeea 	:	val_out <= 4'h0b19;
         4'haeeb 	:	val_out <= 4'h0b19;
         4'haef0 	:	val_out <= 4'h0b0f;
         4'haef1 	:	val_out <= 4'h0b0f;
         4'haef2 	:	val_out <= 4'h0b0f;
         4'haef3 	:	val_out <= 4'h0b0f;
         4'haef8 	:	val_out <= 4'h0b05;
         4'haef9 	:	val_out <= 4'h0b05;
         4'haefa 	:	val_out <= 4'h0b05;
         4'haefb 	:	val_out <= 4'h0b05;
         4'haf00 	:	val_out <= 4'h0afb;
         4'haf01 	:	val_out <= 4'h0afb;
         4'haf02 	:	val_out <= 4'h0afb;
         4'haf03 	:	val_out <= 4'h0afb;
         4'haf08 	:	val_out <= 4'h0af0;
         4'haf09 	:	val_out <= 4'h0af0;
         4'haf0a 	:	val_out <= 4'h0af0;
         4'haf0b 	:	val_out <= 4'h0af0;
         4'haf10 	:	val_out <= 4'h0ae6;
         4'haf11 	:	val_out <= 4'h0ae6;
         4'haf12 	:	val_out <= 4'h0ae6;
         4'haf13 	:	val_out <= 4'h0ae6;
         4'haf18 	:	val_out <= 4'h0adc;
         4'haf19 	:	val_out <= 4'h0adc;
         4'haf1a 	:	val_out <= 4'h0adc;
         4'haf1b 	:	val_out <= 4'h0adc;
         4'haf20 	:	val_out <= 4'h0ad2;
         4'haf21 	:	val_out <= 4'h0ad2;
         4'haf22 	:	val_out <= 4'h0ad2;
         4'haf23 	:	val_out <= 4'h0ad2;
         4'haf28 	:	val_out <= 4'h0ac8;
         4'haf29 	:	val_out <= 4'h0ac8;
         4'haf2a 	:	val_out <= 4'h0ac8;
         4'haf2b 	:	val_out <= 4'h0ac8;
         4'haf30 	:	val_out <= 4'h0abe;
         4'haf31 	:	val_out <= 4'h0abe;
         4'haf32 	:	val_out <= 4'h0abe;
         4'haf33 	:	val_out <= 4'h0abe;
         4'haf38 	:	val_out <= 4'h0ab4;
         4'haf39 	:	val_out <= 4'h0ab4;
         4'haf3a 	:	val_out <= 4'h0ab4;
         4'haf3b 	:	val_out <= 4'h0ab4;
         4'haf40 	:	val_out <= 4'h0aaa;
         4'haf41 	:	val_out <= 4'h0aaa;
         4'haf42 	:	val_out <= 4'h0aaa;
         4'haf43 	:	val_out <= 4'h0aaa;
         4'haf48 	:	val_out <= 4'h0aa0;
         4'haf49 	:	val_out <= 4'h0aa0;
         4'haf4a 	:	val_out <= 4'h0aa0;
         4'haf4b 	:	val_out <= 4'h0aa0;
         4'haf50 	:	val_out <= 4'h0a96;
         4'haf51 	:	val_out <= 4'h0a96;
         4'haf52 	:	val_out <= 4'h0a96;
         4'haf53 	:	val_out <= 4'h0a96;
         4'haf58 	:	val_out <= 4'h0a8c;
         4'haf59 	:	val_out <= 4'h0a8c;
         4'haf5a 	:	val_out <= 4'h0a8c;
         4'haf5b 	:	val_out <= 4'h0a8c;
         4'haf60 	:	val_out <= 4'h0a82;
         4'haf61 	:	val_out <= 4'h0a82;
         4'haf62 	:	val_out <= 4'h0a82;
         4'haf63 	:	val_out <= 4'h0a82;
         4'haf68 	:	val_out <= 4'h0a78;
         4'haf69 	:	val_out <= 4'h0a78;
         4'haf6a 	:	val_out <= 4'h0a78;
         4'haf6b 	:	val_out <= 4'h0a78;
         4'haf70 	:	val_out <= 4'h0a6e;
         4'haf71 	:	val_out <= 4'h0a6e;
         4'haf72 	:	val_out <= 4'h0a6e;
         4'haf73 	:	val_out <= 4'h0a6e;
         4'haf78 	:	val_out <= 4'h0a64;
         4'haf79 	:	val_out <= 4'h0a64;
         4'haf7a 	:	val_out <= 4'h0a64;
         4'haf7b 	:	val_out <= 4'h0a64;
         4'haf80 	:	val_out <= 4'h0a5a;
         4'haf81 	:	val_out <= 4'h0a5a;
         4'haf82 	:	val_out <= 4'h0a5a;
         4'haf83 	:	val_out <= 4'h0a5a;
         4'haf88 	:	val_out <= 4'h0a50;
         4'haf89 	:	val_out <= 4'h0a50;
         4'haf8a 	:	val_out <= 4'h0a50;
         4'haf8b 	:	val_out <= 4'h0a50;
         4'haf90 	:	val_out <= 4'h0a46;
         4'haf91 	:	val_out <= 4'h0a46;
         4'haf92 	:	val_out <= 4'h0a46;
         4'haf93 	:	val_out <= 4'h0a46;
         4'haf98 	:	val_out <= 4'h0a3c;
         4'haf99 	:	val_out <= 4'h0a3c;
         4'haf9a 	:	val_out <= 4'h0a3c;
         4'haf9b 	:	val_out <= 4'h0a3c;
         4'hafa0 	:	val_out <= 4'h0a33;
         4'hafa1 	:	val_out <= 4'h0a33;
         4'hafa2 	:	val_out <= 4'h0a33;
         4'hafa3 	:	val_out <= 4'h0a33;
         4'hafa8 	:	val_out <= 4'h0a29;
         4'hafa9 	:	val_out <= 4'h0a29;
         4'hafaa 	:	val_out <= 4'h0a29;
         4'hafab 	:	val_out <= 4'h0a29;
         4'hafb0 	:	val_out <= 4'h0a1f;
         4'hafb1 	:	val_out <= 4'h0a1f;
         4'hafb2 	:	val_out <= 4'h0a1f;
         4'hafb3 	:	val_out <= 4'h0a1f;
         4'hafb8 	:	val_out <= 4'h0a15;
         4'hafb9 	:	val_out <= 4'h0a15;
         4'hafba 	:	val_out <= 4'h0a15;
         4'hafbb 	:	val_out <= 4'h0a15;
         4'hafc0 	:	val_out <= 4'h0a0b;
         4'hafc1 	:	val_out <= 4'h0a0b;
         4'hafc2 	:	val_out <= 4'h0a0b;
         4'hafc3 	:	val_out <= 4'h0a0b;
         4'hafc8 	:	val_out <= 4'h0a02;
         4'hafc9 	:	val_out <= 4'h0a02;
         4'hafca 	:	val_out <= 4'h0a02;
         4'hafcb 	:	val_out <= 4'h0a02;
         4'hafd0 	:	val_out <= 4'h09f8;
         4'hafd1 	:	val_out <= 4'h09f8;
         4'hafd2 	:	val_out <= 4'h09f8;
         4'hafd3 	:	val_out <= 4'h09f8;
         4'hafd8 	:	val_out <= 4'h09ee;
         4'hafd9 	:	val_out <= 4'h09ee;
         4'hafda 	:	val_out <= 4'h09ee;
         4'hafdb 	:	val_out <= 4'h09ee;
         4'hafe0 	:	val_out <= 4'h09e4;
         4'hafe1 	:	val_out <= 4'h09e4;
         4'hafe2 	:	val_out <= 4'h09e4;
         4'hafe3 	:	val_out <= 4'h09e4;
         4'hafe8 	:	val_out <= 4'h09db;
         4'hafe9 	:	val_out <= 4'h09db;
         4'hafea 	:	val_out <= 4'h09db;
         4'hafeb 	:	val_out <= 4'h09db;
         4'haff0 	:	val_out <= 4'h09d1;
         4'haff1 	:	val_out <= 4'h09d1;
         4'haff2 	:	val_out <= 4'h09d1;
         4'haff3 	:	val_out <= 4'h09d1;
         4'haff8 	:	val_out <= 4'h09c7;
         4'haff9 	:	val_out <= 4'h09c7;
         4'haffa 	:	val_out <= 4'h09c7;
         4'haffb 	:	val_out <= 4'h09c7;
         4'hb000 	:	val_out <= 4'h09be;
         4'hb001 	:	val_out <= 4'h09be;
         4'hb002 	:	val_out <= 4'h09be;
         4'hb003 	:	val_out <= 4'h09be;
         4'hb008 	:	val_out <= 4'h09b4;
         4'hb009 	:	val_out <= 4'h09b4;
         4'hb00a 	:	val_out <= 4'h09b4;
         4'hb00b 	:	val_out <= 4'h09b4;
         4'hb010 	:	val_out <= 4'h09ab;
         4'hb011 	:	val_out <= 4'h09ab;
         4'hb012 	:	val_out <= 4'h09ab;
         4'hb013 	:	val_out <= 4'h09ab;
         4'hb018 	:	val_out <= 4'h09a1;
         4'hb019 	:	val_out <= 4'h09a1;
         4'hb01a 	:	val_out <= 4'h09a1;
         4'hb01b 	:	val_out <= 4'h09a1;
         4'hb020 	:	val_out <= 4'h0997;
         4'hb021 	:	val_out <= 4'h0997;
         4'hb022 	:	val_out <= 4'h0997;
         4'hb023 	:	val_out <= 4'h0997;
         4'hb028 	:	val_out <= 4'h098e;
         4'hb029 	:	val_out <= 4'h098e;
         4'hb02a 	:	val_out <= 4'h098e;
         4'hb02b 	:	val_out <= 4'h098e;
         4'hb030 	:	val_out <= 4'h0984;
         4'hb031 	:	val_out <= 4'h0984;
         4'hb032 	:	val_out <= 4'h0984;
         4'hb033 	:	val_out <= 4'h0984;
         4'hb038 	:	val_out <= 4'h097b;
         4'hb039 	:	val_out <= 4'h097b;
         4'hb03a 	:	val_out <= 4'h097b;
         4'hb03b 	:	val_out <= 4'h097b;
         4'hb040 	:	val_out <= 4'h0971;
         4'hb041 	:	val_out <= 4'h0971;
         4'hb042 	:	val_out <= 4'h0971;
         4'hb043 	:	val_out <= 4'h0971;
         4'hb048 	:	val_out <= 4'h0968;
         4'hb049 	:	val_out <= 4'h0968;
         4'hb04a 	:	val_out <= 4'h0968;
         4'hb04b 	:	val_out <= 4'h0968;
         4'hb050 	:	val_out <= 4'h095f;
         4'hb051 	:	val_out <= 4'h095f;
         4'hb052 	:	val_out <= 4'h095f;
         4'hb053 	:	val_out <= 4'h095f;
         4'hb058 	:	val_out <= 4'h0955;
         4'hb059 	:	val_out <= 4'h0955;
         4'hb05a 	:	val_out <= 4'h0955;
         4'hb05b 	:	val_out <= 4'h0955;
         4'hb060 	:	val_out <= 4'h094c;
         4'hb061 	:	val_out <= 4'h094c;
         4'hb062 	:	val_out <= 4'h094c;
         4'hb063 	:	val_out <= 4'h094c;
         4'hb068 	:	val_out <= 4'h0942;
         4'hb069 	:	val_out <= 4'h0942;
         4'hb06a 	:	val_out <= 4'h0942;
         4'hb06b 	:	val_out <= 4'h0942;
         4'hb070 	:	val_out <= 4'h0939;
         4'hb071 	:	val_out <= 4'h0939;
         4'hb072 	:	val_out <= 4'h0939;
         4'hb073 	:	val_out <= 4'h0939;
         4'hb078 	:	val_out <= 4'h0930;
         4'hb079 	:	val_out <= 4'h0930;
         4'hb07a 	:	val_out <= 4'h0930;
         4'hb07b 	:	val_out <= 4'h0930;
         4'hb080 	:	val_out <= 4'h0926;
         4'hb081 	:	val_out <= 4'h0926;
         4'hb082 	:	val_out <= 4'h0926;
         4'hb083 	:	val_out <= 4'h0926;
         4'hb088 	:	val_out <= 4'h091d;
         4'hb089 	:	val_out <= 4'h091d;
         4'hb08a 	:	val_out <= 4'h091d;
         4'hb08b 	:	val_out <= 4'h091d;
         4'hb090 	:	val_out <= 4'h0914;
         4'hb091 	:	val_out <= 4'h0914;
         4'hb092 	:	val_out <= 4'h0914;
         4'hb093 	:	val_out <= 4'h0914;
         4'hb098 	:	val_out <= 4'h090a;
         4'hb099 	:	val_out <= 4'h090a;
         4'hb09a 	:	val_out <= 4'h090a;
         4'hb09b 	:	val_out <= 4'h090a;
         4'hb0a0 	:	val_out <= 4'h0901;
         4'hb0a1 	:	val_out <= 4'h0901;
         4'hb0a2 	:	val_out <= 4'h0901;
         4'hb0a3 	:	val_out <= 4'h0901;
         4'hb0a8 	:	val_out <= 4'h08f8;
         4'hb0a9 	:	val_out <= 4'h08f8;
         4'hb0aa 	:	val_out <= 4'h08f8;
         4'hb0ab 	:	val_out <= 4'h08f8;
         4'hb0b0 	:	val_out <= 4'h08ef;
         4'hb0b1 	:	val_out <= 4'h08ef;
         4'hb0b2 	:	val_out <= 4'h08ef;
         4'hb0b3 	:	val_out <= 4'h08ef;
         4'hb0b8 	:	val_out <= 4'h08e5;
         4'hb0b9 	:	val_out <= 4'h08e5;
         4'hb0ba 	:	val_out <= 4'h08e5;
         4'hb0bb 	:	val_out <= 4'h08e5;
         4'hb0c0 	:	val_out <= 4'h08dc;
         4'hb0c1 	:	val_out <= 4'h08dc;
         4'hb0c2 	:	val_out <= 4'h08dc;
         4'hb0c3 	:	val_out <= 4'h08dc;
         4'hb0c8 	:	val_out <= 4'h08d3;
         4'hb0c9 	:	val_out <= 4'h08d3;
         4'hb0ca 	:	val_out <= 4'h08d3;
         4'hb0cb 	:	val_out <= 4'h08d3;
         4'hb0d0 	:	val_out <= 4'h08ca;
         4'hb0d1 	:	val_out <= 4'h08ca;
         4'hb0d2 	:	val_out <= 4'h08ca;
         4'hb0d3 	:	val_out <= 4'h08ca;
         4'hb0d8 	:	val_out <= 4'h08c1;
         4'hb0d9 	:	val_out <= 4'h08c1;
         4'hb0da 	:	val_out <= 4'h08c1;
         4'hb0db 	:	val_out <= 4'h08c1;
         4'hb0e0 	:	val_out <= 4'h08b8;
         4'hb0e1 	:	val_out <= 4'h08b8;
         4'hb0e2 	:	val_out <= 4'h08b8;
         4'hb0e3 	:	val_out <= 4'h08b8;
         4'hb0e8 	:	val_out <= 4'h08ae;
         4'hb0e9 	:	val_out <= 4'h08ae;
         4'hb0ea 	:	val_out <= 4'h08ae;
         4'hb0eb 	:	val_out <= 4'h08ae;
         4'hb0f0 	:	val_out <= 4'h08a5;
         4'hb0f1 	:	val_out <= 4'h08a5;
         4'hb0f2 	:	val_out <= 4'h08a5;
         4'hb0f3 	:	val_out <= 4'h08a5;
         4'hb0f8 	:	val_out <= 4'h089c;
         4'hb0f9 	:	val_out <= 4'h089c;
         4'hb0fa 	:	val_out <= 4'h089c;
         4'hb0fb 	:	val_out <= 4'h089c;
         4'hb100 	:	val_out <= 4'h0893;
         4'hb101 	:	val_out <= 4'h0893;
         4'hb102 	:	val_out <= 4'h0893;
         4'hb103 	:	val_out <= 4'h0893;
         4'hb108 	:	val_out <= 4'h088a;
         4'hb109 	:	val_out <= 4'h088a;
         4'hb10a 	:	val_out <= 4'h088a;
         4'hb10b 	:	val_out <= 4'h088a;
         4'hb110 	:	val_out <= 4'h0881;
         4'hb111 	:	val_out <= 4'h0881;
         4'hb112 	:	val_out <= 4'h0881;
         4'hb113 	:	val_out <= 4'h0881;
         4'hb118 	:	val_out <= 4'h0878;
         4'hb119 	:	val_out <= 4'h0878;
         4'hb11a 	:	val_out <= 4'h0878;
         4'hb11b 	:	val_out <= 4'h0878;
         4'hb120 	:	val_out <= 4'h086f;
         4'hb121 	:	val_out <= 4'h086f;
         4'hb122 	:	val_out <= 4'h086f;
         4'hb123 	:	val_out <= 4'h086f;
         4'hb128 	:	val_out <= 4'h0866;
         4'hb129 	:	val_out <= 4'h0866;
         4'hb12a 	:	val_out <= 4'h0866;
         4'hb12b 	:	val_out <= 4'h0866;
         4'hb130 	:	val_out <= 4'h085d;
         4'hb131 	:	val_out <= 4'h085d;
         4'hb132 	:	val_out <= 4'h085d;
         4'hb133 	:	val_out <= 4'h085d;
         4'hb138 	:	val_out <= 4'h0854;
         4'hb139 	:	val_out <= 4'h0854;
         4'hb13a 	:	val_out <= 4'h0854;
         4'hb13b 	:	val_out <= 4'h0854;
         4'hb140 	:	val_out <= 4'h084b;
         4'hb141 	:	val_out <= 4'h084b;
         4'hb142 	:	val_out <= 4'h084b;
         4'hb143 	:	val_out <= 4'h084b;
         4'hb148 	:	val_out <= 4'h0843;
         4'hb149 	:	val_out <= 4'h0843;
         4'hb14a 	:	val_out <= 4'h0843;
         4'hb14b 	:	val_out <= 4'h0843;
         4'hb150 	:	val_out <= 4'h083a;
         4'hb151 	:	val_out <= 4'h083a;
         4'hb152 	:	val_out <= 4'h083a;
         4'hb153 	:	val_out <= 4'h083a;
         4'hb158 	:	val_out <= 4'h0831;
         4'hb159 	:	val_out <= 4'h0831;
         4'hb15a 	:	val_out <= 4'h0831;
         4'hb15b 	:	val_out <= 4'h0831;
         4'hb160 	:	val_out <= 4'h0828;
         4'hb161 	:	val_out <= 4'h0828;
         4'hb162 	:	val_out <= 4'h0828;
         4'hb163 	:	val_out <= 4'h0828;
         4'hb168 	:	val_out <= 4'h081f;
         4'hb169 	:	val_out <= 4'h081f;
         4'hb16a 	:	val_out <= 4'h081f;
         4'hb16b 	:	val_out <= 4'h081f;
         4'hb170 	:	val_out <= 4'h0816;
         4'hb171 	:	val_out <= 4'h0816;
         4'hb172 	:	val_out <= 4'h0816;
         4'hb173 	:	val_out <= 4'h0816;
         4'hb178 	:	val_out <= 4'h080e;
         4'hb179 	:	val_out <= 4'h080e;
         4'hb17a 	:	val_out <= 4'h080e;
         4'hb17b 	:	val_out <= 4'h080e;
         4'hb180 	:	val_out <= 4'h0805;
         4'hb181 	:	val_out <= 4'h0805;
         4'hb182 	:	val_out <= 4'h0805;
         4'hb183 	:	val_out <= 4'h0805;
         4'hb188 	:	val_out <= 4'h07fc;
         4'hb189 	:	val_out <= 4'h07fc;
         4'hb18a 	:	val_out <= 4'h07fc;
         4'hb18b 	:	val_out <= 4'h07fc;
         4'hb190 	:	val_out <= 4'h07f3;
         4'hb191 	:	val_out <= 4'h07f3;
         4'hb192 	:	val_out <= 4'h07f3;
         4'hb193 	:	val_out <= 4'h07f3;
         4'hb198 	:	val_out <= 4'h07eb;
         4'hb199 	:	val_out <= 4'h07eb;
         4'hb19a 	:	val_out <= 4'h07eb;
         4'hb19b 	:	val_out <= 4'h07eb;
         4'hb1a0 	:	val_out <= 4'h07e2;
         4'hb1a1 	:	val_out <= 4'h07e2;
         4'hb1a2 	:	val_out <= 4'h07e2;
         4'hb1a3 	:	val_out <= 4'h07e2;
         4'hb1a8 	:	val_out <= 4'h07d9;
         4'hb1a9 	:	val_out <= 4'h07d9;
         4'hb1aa 	:	val_out <= 4'h07d9;
         4'hb1ab 	:	val_out <= 4'h07d9;
         4'hb1b0 	:	val_out <= 4'h07d1;
         4'hb1b1 	:	val_out <= 4'h07d1;
         4'hb1b2 	:	val_out <= 4'h07d1;
         4'hb1b3 	:	val_out <= 4'h07d1;
         4'hb1b8 	:	val_out <= 4'h07c8;
         4'hb1b9 	:	val_out <= 4'h07c8;
         4'hb1ba 	:	val_out <= 4'h07c8;
         4'hb1bb 	:	val_out <= 4'h07c8;
         4'hb1c0 	:	val_out <= 4'h07bf;
         4'hb1c1 	:	val_out <= 4'h07bf;
         4'hb1c2 	:	val_out <= 4'h07bf;
         4'hb1c3 	:	val_out <= 4'h07bf;
         4'hb1c8 	:	val_out <= 4'h07b7;
         4'hb1c9 	:	val_out <= 4'h07b7;
         4'hb1ca 	:	val_out <= 4'h07b7;
         4'hb1cb 	:	val_out <= 4'h07b7;
         4'hb1d0 	:	val_out <= 4'h07ae;
         4'hb1d1 	:	val_out <= 4'h07ae;
         4'hb1d2 	:	val_out <= 4'h07ae;
         4'hb1d3 	:	val_out <= 4'h07ae;
         4'hb1d8 	:	val_out <= 4'h07a6;
         4'hb1d9 	:	val_out <= 4'h07a6;
         4'hb1da 	:	val_out <= 4'h07a6;
         4'hb1db 	:	val_out <= 4'h07a6;
         4'hb1e0 	:	val_out <= 4'h079d;
         4'hb1e1 	:	val_out <= 4'h079d;
         4'hb1e2 	:	val_out <= 4'h079d;
         4'hb1e3 	:	val_out <= 4'h079d;
         4'hb1e8 	:	val_out <= 4'h0794;
         4'hb1e9 	:	val_out <= 4'h0794;
         4'hb1ea 	:	val_out <= 4'h0794;
         4'hb1eb 	:	val_out <= 4'h0794;
         4'hb1f0 	:	val_out <= 4'h078c;
         4'hb1f1 	:	val_out <= 4'h078c;
         4'hb1f2 	:	val_out <= 4'h078c;
         4'hb1f3 	:	val_out <= 4'h078c;
         4'hb1f8 	:	val_out <= 4'h0783;
         4'hb1f9 	:	val_out <= 4'h0783;
         4'hb1fa 	:	val_out <= 4'h0783;
         4'hb1fb 	:	val_out <= 4'h0783;
         4'hb200 	:	val_out <= 4'h077b;
         4'hb201 	:	val_out <= 4'h077b;
         4'hb202 	:	val_out <= 4'h077b;
         4'hb203 	:	val_out <= 4'h077b;
         4'hb208 	:	val_out <= 4'h0773;
         4'hb209 	:	val_out <= 4'h0773;
         4'hb20a 	:	val_out <= 4'h0773;
         4'hb20b 	:	val_out <= 4'h0773;
         4'hb210 	:	val_out <= 4'h076a;
         4'hb211 	:	val_out <= 4'h076a;
         4'hb212 	:	val_out <= 4'h076a;
         4'hb213 	:	val_out <= 4'h076a;
         4'hb218 	:	val_out <= 4'h0762;
         4'hb219 	:	val_out <= 4'h0762;
         4'hb21a 	:	val_out <= 4'h0762;
         4'hb21b 	:	val_out <= 4'h0762;
         4'hb220 	:	val_out <= 4'h0759;
         4'hb221 	:	val_out <= 4'h0759;
         4'hb222 	:	val_out <= 4'h0759;
         4'hb223 	:	val_out <= 4'h0759;
         4'hb228 	:	val_out <= 4'h0751;
         4'hb229 	:	val_out <= 4'h0751;
         4'hb22a 	:	val_out <= 4'h0751;
         4'hb22b 	:	val_out <= 4'h0751;
         4'hb230 	:	val_out <= 4'h0749;
         4'hb231 	:	val_out <= 4'h0749;
         4'hb232 	:	val_out <= 4'h0749;
         4'hb233 	:	val_out <= 4'h0749;
         4'hb238 	:	val_out <= 4'h0740;
         4'hb239 	:	val_out <= 4'h0740;
         4'hb23a 	:	val_out <= 4'h0740;
         4'hb23b 	:	val_out <= 4'h0740;
         4'hb240 	:	val_out <= 4'h0738;
         4'hb241 	:	val_out <= 4'h0738;
         4'hb242 	:	val_out <= 4'h0738;
         4'hb243 	:	val_out <= 4'h0738;
         4'hb248 	:	val_out <= 4'h0730;
         4'hb249 	:	val_out <= 4'h0730;
         4'hb24a 	:	val_out <= 4'h0730;
         4'hb24b 	:	val_out <= 4'h0730;
         4'hb250 	:	val_out <= 4'h0727;
         4'hb251 	:	val_out <= 4'h0727;
         4'hb252 	:	val_out <= 4'h0727;
         4'hb253 	:	val_out <= 4'h0727;
         4'hb258 	:	val_out <= 4'h071f;
         4'hb259 	:	val_out <= 4'h071f;
         4'hb25a 	:	val_out <= 4'h071f;
         4'hb25b 	:	val_out <= 4'h071f;
         4'hb260 	:	val_out <= 4'h0717;
         4'hb261 	:	val_out <= 4'h0717;
         4'hb262 	:	val_out <= 4'h0717;
         4'hb263 	:	val_out <= 4'h0717;
         4'hb268 	:	val_out <= 4'h070e;
         4'hb269 	:	val_out <= 4'h070e;
         4'hb26a 	:	val_out <= 4'h070e;
         4'hb26b 	:	val_out <= 4'h070e;
         4'hb270 	:	val_out <= 4'h0706;
         4'hb271 	:	val_out <= 4'h0706;
         4'hb272 	:	val_out <= 4'h0706;
         4'hb273 	:	val_out <= 4'h0706;
         4'hb278 	:	val_out <= 4'h06fe;
         4'hb279 	:	val_out <= 4'h06fe;
         4'hb27a 	:	val_out <= 4'h06fe;
         4'hb27b 	:	val_out <= 4'h06fe;
         4'hb280 	:	val_out <= 4'h06f6;
         4'hb281 	:	val_out <= 4'h06f6;
         4'hb282 	:	val_out <= 4'h06f6;
         4'hb283 	:	val_out <= 4'h06f6;
         4'hb288 	:	val_out <= 4'h06ee;
         4'hb289 	:	val_out <= 4'h06ee;
         4'hb28a 	:	val_out <= 4'h06ee;
         4'hb28b 	:	val_out <= 4'h06ee;
         4'hb290 	:	val_out <= 4'h06e6;
         4'hb291 	:	val_out <= 4'h06e6;
         4'hb292 	:	val_out <= 4'h06e6;
         4'hb293 	:	val_out <= 4'h06e6;
         4'hb298 	:	val_out <= 4'h06dd;
         4'hb299 	:	val_out <= 4'h06dd;
         4'hb29a 	:	val_out <= 4'h06dd;
         4'hb29b 	:	val_out <= 4'h06dd;
         4'hb2a0 	:	val_out <= 4'h06d5;
         4'hb2a1 	:	val_out <= 4'h06d5;
         4'hb2a2 	:	val_out <= 4'h06d5;
         4'hb2a3 	:	val_out <= 4'h06d5;
         4'hb2a8 	:	val_out <= 4'h06cd;
         4'hb2a9 	:	val_out <= 4'h06cd;
         4'hb2aa 	:	val_out <= 4'h06cd;
         4'hb2ab 	:	val_out <= 4'h06cd;
         4'hb2b0 	:	val_out <= 4'h06c5;
         4'hb2b1 	:	val_out <= 4'h06c5;
         4'hb2b2 	:	val_out <= 4'h06c5;
         4'hb2b3 	:	val_out <= 4'h06c5;
         4'hb2b8 	:	val_out <= 4'h06bd;
         4'hb2b9 	:	val_out <= 4'h06bd;
         4'hb2ba 	:	val_out <= 4'h06bd;
         4'hb2bb 	:	val_out <= 4'h06bd;
         4'hb2c0 	:	val_out <= 4'h06b5;
         4'hb2c1 	:	val_out <= 4'h06b5;
         4'hb2c2 	:	val_out <= 4'h06b5;
         4'hb2c3 	:	val_out <= 4'h06b5;
         4'hb2c8 	:	val_out <= 4'h06ad;
         4'hb2c9 	:	val_out <= 4'h06ad;
         4'hb2ca 	:	val_out <= 4'h06ad;
         4'hb2cb 	:	val_out <= 4'h06ad;
         4'hb2d0 	:	val_out <= 4'h06a5;
         4'hb2d1 	:	val_out <= 4'h06a5;
         4'hb2d2 	:	val_out <= 4'h06a5;
         4'hb2d3 	:	val_out <= 4'h06a5;
         4'hb2d8 	:	val_out <= 4'h069d;
         4'hb2d9 	:	val_out <= 4'h069d;
         4'hb2da 	:	val_out <= 4'h069d;
         4'hb2db 	:	val_out <= 4'h069d;
         4'hb2e0 	:	val_out <= 4'h0695;
         4'hb2e1 	:	val_out <= 4'h0695;
         4'hb2e2 	:	val_out <= 4'h0695;
         4'hb2e3 	:	val_out <= 4'h0695;
         4'hb2e8 	:	val_out <= 4'h068d;
         4'hb2e9 	:	val_out <= 4'h068d;
         4'hb2ea 	:	val_out <= 4'h068d;
         4'hb2eb 	:	val_out <= 4'h068d;
         4'hb2f0 	:	val_out <= 4'h0685;
         4'hb2f1 	:	val_out <= 4'h0685;
         4'hb2f2 	:	val_out <= 4'h0685;
         4'hb2f3 	:	val_out <= 4'h0685;
         4'hb2f8 	:	val_out <= 4'h067d;
         4'hb2f9 	:	val_out <= 4'h067d;
         4'hb2fa 	:	val_out <= 4'h067d;
         4'hb2fb 	:	val_out <= 4'h067d;
         4'hb300 	:	val_out <= 4'h0675;
         4'hb301 	:	val_out <= 4'h0675;
         4'hb302 	:	val_out <= 4'h0675;
         4'hb303 	:	val_out <= 4'h0675;
         4'hb308 	:	val_out <= 4'h066d;
         4'hb309 	:	val_out <= 4'h066d;
         4'hb30a 	:	val_out <= 4'h066d;
         4'hb30b 	:	val_out <= 4'h066d;
         4'hb310 	:	val_out <= 4'h0666;
         4'hb311 	:	val_out <= 4'h0666;
         4'hb312 	:	val_out <= 4'h0666;
         4'hb313 	:	val_out <= 4'h0666;
         4'hb318 	:	val_out <= 4'h065e;
         4'hb319 	:	val_out <= 4'h065e;
         4'hb31a 	:	val_out <= 4'h065e;
         4'hb31b 	:	val_out <= 4'h065e;
         4'hb320 	:	val_out <= 4'h0656;
         4'hb321 	:	val_out <= 4'h0656;
         4'hb322 	:	val_out <= 4'h0656;
         4'hb323 	:	val_out <= 4'h0656;
         4'hb328 	:	val_out <= 4'h064e;
         4'hb329 	:	val_out <= 4'h064e;
         4'hb32a 	:	val_out <= 4'h064e;
         4'hb32b 	:	val_out <= 4'h064e;
         4'hb330 	:	val_out <= 4'h0646;
         4'hb331 	:	val_out <= 4'h0646;
         4'hb332 	:	val_out <= 4'h0646;
         4'hb333 	:	val_out <= 4'h0646;
         4'hb338 	:	val_out <= 4'h063f;
         4'hb339 	:	val_out <= 4'h063f;
         4'hb33a 	:	val_out <= 4'h063f;
         4'hb33b 	:	val_out <= 4'h063f;
         4'hb340 	:	val_out <= 4'h0637;
         4'hb341 	:	val_out <= 4'h0637;
         4'hb342 	:	val_out <= 4'h0637;
         4'hb343 	:	val_out <= 4'h0637;
         4'hb348 	:	val_out <= 4'h062f;
         4'hb349 	:	val_out <= 4'h062f;
         4'hb34a 	:	val_out <= 4'h062f;
         4'hb34b 	:	val_out <= 4'h062f;
         4'hb350 	:	val_out <= 4'h0627;
         4'hb351 	:	val_out <= 4'h0627;
         4'hb352 	:	val_out <= 4'h0627;
         4'hb353 	:	val_out <= 4'h0627;
         4'hb358 	:	val_out <= 4'h0620;
         4'hb359 	:	val_out <= 4'h0620;
         4'hb35a 	:	val_out <= 4'h0620;
         4'hb35b 	:	val_out <= 4'h0620;
         4'hb360 	:	val_out <= 4'h0618;
         4'hb361 	:	val_out <= 4'h0618;
         4'hb362 	:	val_out <= 4'h0618;
         4'hb363 	:	val_out <= 4'h0618;
         4'hb368 	:	val_out <= 4'h0610;
         4'hb369 	:	val_out <= 4'h0610;
         4'hb36a 	:	val_out <= 4'h0610;
         4'hb36b 	:	val_out <= 4'h0610;
         4'hb370 	:	val_out <= 4'h0609;
         4'hb371 	:	val_out <= 4'h0609;
         4'hb372 	:	val_out <= 4'h0609;
         4'hb373 	:	val_out <= 4'h0609;
         4'hb378 	:	val_out <= 4'h0601;
         4'hb379 	:	val_out <= 4'h0601;
         4'hb37a 	:	val_out <= 4'h0601;
         4'hb37b 	:	val_out <= 4'h0601;
         4'hb380 	:	val_out <= 4'h05fa;
         4'hb381 	:	val_out <= 4'h05fa;
         4'hb382 	:	val_out <= 4'h05fa;
         4'hb383 	:	val_out <= 4'h05fa;
         4'hb388 	:	val_out <= 4'h05f2;
         4'hb389 	:	val_out <= 4'h05f2;
         4'hb38a 	:	val_out <= 4'h05f2;
         4'hb38b 	:	val_out <= 4'h05f2;
         4'hb390 	:	val_out <= 4'h05ea;
         4'hb391 	:	val_out <= 4'h05ea;
         4'hb392 	:	val_out <= 4'h05ea;
         4'hb393 	:	val_out <= 4'h05ea;
         4'hb398 	:	val_out <= 4'h05e3;
         4'hb399 	:	val_out <= 4'h05e3;
         4'hb39a 	:	val_out <= 4'h05e3;
         4'hb39b 	:	val_out <= 4'h05e3;
         4'hb3a0 	:	val_out <= 4'h05db;
         4'hb3a1 	:	val_out <= 4'h05db;
         4'hb3a2 	:	val_out <= 4'h05db;
         4'hb3a3 	:	val_out <= 4'h05db;
         4'hb3a8 	:	val_out <= 4'h05d4;
         4'hb3a9 	:	val_out <= 4'h05d4;
         4'hb3aa 	:	val_out <= 4'h05d4;
         4'hb3ab 	:	val_out <= 4'h05d4;
         4'hb3b0 	:	val_out <= 4'h05cc;
         4'hb3b1 	:	val_out <= 4'h05cc;
         4'hb3b2 	:	val_out <= 4'h05cc;
         4'hb3b3 	:	val_out <= 4'h05cc;
         4'hb3b8 	:	val_out <= 4'h05c5;
         4'hb3b9 	:	val_out <= 4'h05c5;
         4'hb3ba 	:	val_out <= 4'h05c5;
         4'hb3bb 	:	val_out <= 4'h05c5;
         4'hb3c0 	:	val_out <= 4'h05bd;
         4'hb3c1 	:	val_out <= 4'h05bd;
         4'hb3c2 	:	val_out <= 4'h05bd;
         4'hb3c3 	:	val_out <= 4'h05bd;
         4'hb3c8 	:	val_out <= 4'h05b6;
         4'hb3c9 	:	val_out <= 4'h05b6;
         4'hb3ca 	:	val_out <= 4'h05b6;
         4'hb3cb 	:	val_out <= 4'h05b6;
         4'hb3d0 	:	val_out <= 4'h05af;
         4'hb3d1 	:	val_out <= 4'h05af;
         4'hb3d2 	:	val_out <= 4'h05af;
         4'hb3d3 	:	val_out <= 4'h05af;
         4'hb3d8 	:	val_out <= 4'h05a7;
         4'hb3d9 	:	val_out <= 4'h05a7;
         4'hb3da 	:	val_out <= 4'h05a7;
         4'hb3db 	:	val_out <= 4'h05a7;
         4'hb3e0 	:	val_out <= 4'h05a0;
         4'hb3e1 	:	val_out <= 4'h05a0;
         4'hb3e2 	:	val_out <= 4'h05a0;
         4'hb3e3 	:	val_out <= 4'h05a0;
         4'hb3e8 	:	val_out <= 4'h0598;
         4'hb3e9 	:	val_out <= 4'h0598;
         4'hb3ea 	:	val_out <= 4'h0598;
         4'hb3eb 	:	val_out <= 4'h0598;
         4'hb3f0 	:	val_out <= 4'h0591;
         4'hb3f1 	:	val_out <= 4'h0591;
         4'hb3f2 	:	val_out <= 4'h0591;
         4'hb3f3 	:	val_out <= 4'h0591;
         4'hb3f8 	:	val_out <= 4'h058a;
         4'hb3f9 	:	val_out <= 4'h058a;
         4'hb3fa 	:	val_out <= 4'h058a;
         4'hb3fb 	:	val_out <= 4'h058a;
         4'hb400 	:	val_out <= 4'h0582;
         4'hb401 	:	val_out <= 4'h0582;
         4'hb402 	:	val_out <= 4'h0582;
         4'hb403 	:	val_out <= 4'h0582;
         4'hb408 	:	val_out <= 4'h057b;
         4'hb409 	:	val_out <= 4'h057b;
         4'hb40a 	:	val_out <= 4'h057b;
         4'hb40b 	:	val_out <= 4'h057b;
         4'hb410 	:	val_out <= 4'h0574;
         4'hb411 	:	val_out <= 4'h0574;
         4'hb412 	:	val_out <= 4'h0574;
         4'hb413 	:	val_out <= 4'h0574;
         4'hb418 	:	val_out <= 4'h056d;
         4'hb419 	:	val_out <= 4'h056d;
         4'hb41a 	:	val_out <= 4'h056d;
         4'hb41b 	:	val_out <= 4'h056d;
         4'hb420 	:	val_out <= 4'h0565;
         4'hb421 	:	val_out <= 4'h0565;
         4'hb422 	:	val_out <= 4'h0565;
         4'hb423 	:	val_out <= 4'h0565;
         4'hb428 	:	val_out <= 4'h055e;
         4'hb429 	:	val_out <= 4'h055e;
         4'hb42a 	:	val_out <= 4'h055e;
         4'hb42b 	:	val_out <= 4'h055e;
         4'hb430 	:	val_out <= 4'h0557;
         4'hb431 	:	val_out <= 4'h0557;
         4'hb432 	:	val_out <= 4'h0557;
         4'hb433 	:	val_out <= 4'h0557;
         4'hb438 	:	val_out <= 4'h0550;
         4'hb439 	:	val_out <= 4'h0550;
         4'hb43a 	:	val_out <= 4'h0550;
         4'hb43b 	:	val_out <= 4'h0550;
         4'hb440 	:	val_out <= 4'h0549;
         4'hb441 	:	val_out <= 4'h0549;
         4'hb442 	:	val_out <= 4'h0549;
         4'hb443 	:	val_out <= 4'h0549;
         4'hb448 	:	val_out <= 4'h0542;
         4'hb449 	:	val_out <= 4'h0542;
         4'hb44a 	:	val_out <= 4'h0542;
         4'hb44b 	:	val_out <= 4'h0542;
         4'hb450 	:	val_out <= 4'h053a;
         4'hb451 	:	val_out <= 4'h053a;
         4'hb452 	:	val_out <= 4'h053a;
         4'hb453 	:	val_out <= 4'h053a;
         4'hb458 	:	val_out <= 4'h0533;
         4'hb459 	:	val_out <= 4'h0533;
         4'hb45a 	:	val_out <= 4'h0533;
         4'hb45b 	:	val_out <= 4'h0533;
         4'hb460 	:	val_out <= 4'h052c;
         4'hb461 	:	val_out <= 4'h052c;
         4'hb462 	:	val_out <= 4'h052c;
         4'hb463 	:	val_out <= 4'h052c;
         4'hb468 	:	val_out <= 4'h0525;
         4'hb469 	:	val_out <= 4'h0525;
         4'hb46a 	:	val_out <= 4'h0525;
         4'hb46b 	:	val_out <= 4'h0525;
         4'hb470 	:	val_out <= 4'h051e;
         4'hb471 	:	val_out <= 4'h051e;
         4'hb472 	:	val_out <= 4'h051e;
         4'hb473 	:	val_out <= 4'h051e;
         4'hb478 	:	val_out <= 4'h0517;
         4'hb479 	:	val_out <= 4'h0517;
         4'hb47a 	:	val_out <= 4'h0517;
         4'hb47b 	:	val_out <= 4'h0517;
         4'hb480 	:	val_out <= 4'h0510;
         4'hb481 	:	val_out <= 4'h0510;
         4'hb482 	:	val_out <= 4'h0510;
         4'hb483 	:	val_out <= 4'h0510;
         4'hb488 	:	val_out <= 4'h0509;
         4'hb489 	:	val_out <= 4'h0509;
         4'hb48a 	:	val_out <= 4'h0509;
         4'hb48b 	:	val_out <= 4'h0509;
         4'hb490 	:	val_out <= 4'h0502;
         4'hb491 	:	val_out <= 4'h0502;
         4'hb492 	:	val_out <= 4'h0502;
         4'hb493 	:	val_out <= 4'h0502;
         4'hb498 	:	val_out <= 4'h04fb;
         4'hb499 	:	val_out <= 4'h04fb;
         4'hb49a 	:	val_out <= 4'h04fb;
         4'hb49b 	:	val_out <= 4'h04fb;
         4'hb4a0 	:	val_out <= 4'h04f4;
         4'hb4a1 	:	val_out <= 4'h04f4;
         4'hb4a2 	:	val_out <= 4'h04f4;
         4'hb4a3 	:	val_out <= 4'h04f4;
         4'hb4a8 	:	val_out <= 4'h04ed;
         4'hb4a9 	:	val_out <= 4'h04ed;
         4'hb4aa 	:	val_out <= 4'h04ed;
         4'hb4ab 	:	val_out <= 4'h04ed;
         4'hb4b0 	:	val_out <= 4'h04e6;
         4'hb4b1 	:	val_out <= 4'h04e6;
         4'hb4b2 	:	val_out <= 4'h04e6;
         4'hb4b3 	:	val_out <= 4'h04e6;
         4'hb4b8 	:	val_out <= 4'h04e0;
         4'hb4b9 	:	val_out <= 4'h04e0;
         4'hb4ba 	:	val_out <= 4'h04e0;
         4'hb4bb 	:	val_out <= 4'h04e0;
         4'hb4c0 	:	val_out <= 4'h04d9;
         4'hb4c1 	:	val_out <= 4'h04d9;
         4'hb4c2 	:	val_out <= 4'h04d9;
         4'hb4c3 	:	val_out <= 4'h04d9;
         4'hb4c8 	:	val_out <= 4'h04d2;
         4'hb4c9 	:	val_out <= 4'h04d2;
         4'hb4ca 	:	val_out <= 4'h04d2;
         4'hb4cb 	:	val_out <= 4'h04d2;
         4'hb4d0 	:	val_out <= 4'h04cb;
         4'hb4d1 	:	val_out <= 4'h04cb;
         4'hb4d2 	:	val_out <= 4'h04cb;
         4'hb4d3 	:	val_out <= 4'h04cb;
         4'hb4d8 	:	val_out <= 4'h04c4;
         4'hb4d9 	:	val_out <= 4'h04c4;
         4'hb4da 	:	val_out <= 4'h04c4;
         4'hb4db 	:	val_out <= 4'h04c4;
         4'hb4e0 	:	val_out <= 4'h04bd;
         4'hb4e1 	:	val_out <= 4'h04bd;
         4'hb4e2 	:	val_out <= 4'h04bd;
         4'hb4e3 	:	val_out <= 4'h04bd;
         4'hb4e8 	:	val_out <= 4'h04b7;
         4'hb4e9 	:	val_out <= 4'h04b7;
         4'hb4ea 	:	val_out <= 4'h04b7;
         4'hb4eb 	:	val_out <= 4'h04b7;
         4'hb4f0 	:	val_out <= 4'h04b0;
         4'hb4f1 	:	val_out <= 4'h04b0;
         4'hb4f2 	:	val_out <= 4'h04b0;
         4'hb4f3 	:	val_out <= 4'h04b0;
         4'hb4f8 	:	val_out <= 4'h04a9;
         4'hb4f9 	:	val_out <= 4'h04a9;
         4'hb4fa 	:	val_out <= 4'h04a9;
         4'hb4fb 	:	val_out <= 4'h04a9;
         4'hb500 	:	val_out <= 4'h04a2;
         4'hb501 	:	val_out <= 4'h04a2;
         4'hb502 	:	val_out <= 4'h04a2;
         4'hb503 	:	val_out <= 4'h04a2;
         4'hb508 	:	val_out <= 4'h049c;
         4'hb509 	:	val_out <= 4'h049c;
         4'hb50a 	:	val_out <= 4'h049c;
         4'hb50b 	:	val_out <= 4'h049c;
         4'hb510 	:	val_out <= 4'h0495;
         4'hb511 	:	val_out <= 4'h0495;
         4'hb512 	:	val_out <= 4'h0495;
         4'hb513 	:	val_out <= 4'h0495;
         4'hb518 	:	val_out <= 4'h048e;
         4'hb519 	:	val_out <= 4'h048e;
         4'hb51a 	:	val_out <= 4'h048e;
         4'hb51b 	:	val_out <= 4'h048e;
         4'hb520 	:	val_out <= 4'h0488;
         4'hb521 	:	val_out <= 4'h0488;
         4'hb522 	:	val_out <= 4'h0488;
         4'hb523 	:	val_out <= 4'h0488;
         4'hb528 	:	val_out <= 4'h0481;
         4'hb529 	:	val_out <= 4'h0481;
         4'hb52a 	:	val_out <= 4'h0481;
         4'hb52b 	:	val_out <= 4'h0481;
         4'hb530 	:	val_out <= 4'h047b;
         4'hb531 	:	val_out <= 4'h047b;
         4'hb532 	:	val_out <= 4'h047b;
         4'hb533 	:	val_out <= 4'h047b;
         4'hb538 	:	val_out <= 4'h0474;
         4'hb539 	:	val_out <= 4'h0474;
         4'hb53a 	:	val_out <= 4'h0474;
         4'hb53b 	:	val_out <= 4'h0474;
         4'hb540 	:	val_out <= 4'h046d;
         4'hb541 	:	val_out <= 4'h046d;
         4'hb542 	:	val_out <= 4'h046d;
         4'hb543 	:	val_out <= 4'h046d;
         4'hb548 	:	val_out <= 4'h0467;
         4'hb549 	:	val_out <= 4'h0467;
         4'hb54a 	:	val_out <= 4'h0467;
         4'hb54b 	:	val_out <= 4'h0467;
         4'hb550 	:	val_out <= 4'h0460;
         4'hb551 	:	val_out <= 4'h0460;
         4'hb552 	:	val_out <= 4'h0460;
         4'hb553 	:	val_out <= 4'h0460;
         4'hb558 	:	val_out <= 4'h045a;
         4'hb559 	:	val_out <= 4'h045a;
         4'hb55a 	:	val_out <= 4'h045a;
         4'hb55b 	:	val_out <= 4'h045a;
         4'hb560 	:	val_out <= 4'h0453;
         4'hb561 	:	val_out <= 4'h0453;
         4'hb562 	:	val_out <= 4'h0453;
         4'hb563 	:	val_out <= 4'h0453;
         4'hb568 	:	val_out <= 4'h044d;
         4'hb569 	:	val_out <= 4'h044d;
         4'hb56a 	:	val_out <= 4'h044d;
         4'hb56b 	:	val_out <= 4'h044d;
         4'hb570 	:	val_out <= 4'h0446;
         4'hb571 	:	val_out <= 4'h0446;
         4'hb572 	:	val_out <= 4'h0446;
         4'hb573 	:	val_out <= 4'h0446;
         4'hb578 	:	val_out <= 4'h0440;
         4'hb579 	:	val_out <= 4'h0440;
         4'hb57a 	:	val_out <= 4'h0440;
         4'hb57b 	:	val_out <= 4'h0440;
         4'hb580 	:	val_out <= 4'h043a;
         4'hb581 	:	val_out <= 4'h043a;
         4'hb582 	:	val_out <= 4'h043a;
         4'hb583 	:	val_out <= 4'h043a;
         4'hb588 	:	val_out <= 4'h0433;
         4'hb589 	:	val_out <= 4'h0433;
         4'hb58a 	:	val_out <= 4'h0433;
         4'hb58b 	:	val_out <= 4'h0433;
         4'hb590 	:	val_out <= 4'h042d;
         4'hb591 	:	val_out <= 4'h042d;
         4'hb592 	:	val_out <= 4'h042d;
         4'hb593 	:	val_out <= 4'h042d;
         4'hb598 	:	val_out <= 4'h0426;
         4'hb599 	:	val_out <= 4'h0426;
         4'hb59a 	:	val_out <= 4'h0426;
         4'hb59b 	:	val_out <= 4'h0426;
         4'hb5a0 	:	val_out <= 4'h0420;
         4'hb5a1 	:	val_out <= 4'h0420;
         4'hb5a2 	:	val_out <= 4'h0420;
         4'hb5a3 	:	val_out <= 4'h0420;
         4'hb5a8 	:	val_out <= 4'h041a;
         4'hb5a9 	:	val_out <= 4'h041a;
         4'hb5aa 	:	val_out <= 4'h041a;
         4'hb5ab 	:	val_out <= 4'h041a;
         4'hb5b0 	:	val_out <= 4'h0414;
         4'hb5b1 	:	val_out <= 4'h0414;
         4'hb5b2 	:	val_out <= 4'h0414;
         4'hb5b3 	:	val_out <= 4'h0414;
         4'hb5b8 	:	val_out <= 4'h040d;
         4'hb5b9 	:	val_out <= 4'h040d;
         4'hb5ba 	:	val_out <= 4'h040d;
         4'hb5bb 	:	val_out <= 4'h040d;
         4'hb5c0 	:	val_out <= 4'h0407;
         4'hb5c1 	:	val_out <= 4'h0407;
         4'hb5c2 	:	val_out <= 4'h0407;
         4'hb5c3 	:	val_out <= 4'h0407;
         4'hb5c8 	:	val_out <= 4'h0401;
         4'hb5c9 	:	val_out <= 4'h0401;
         4'hb5ca 	:	val_out <= 4'h0401;
         4'hb5cb 	:	val_out <= 4'h0401;
         4'hb5d0 	:	val_out <= 4'h03fa;
         4'hb5d1 	:	val_out <= 4'h03fa;
         4'hb5d2 	:	val_out <= 4'h03fa;
         4'hb5d3 	:	val_out <= 4'h03fa;
         4'hb5d8 	:	val_out <= 4'h03f4;
         4'hb5d9 	:	val_out <= 4'h03f4;
         4'hb5da 	:	val_out <= 4'h03f4;
         4'hb5db 	:	val_out <= 4'h03f4;
         4'hb5e0 	:	val_out <= 4'h03ee;
         4'hb5e1 	:	val_out <= 4'h03ee;
         4'hb5e2 	:	val_out <= 4'h03ee;
         4'hb5e3 	:	val_out <= 4'h03ee;
         4'hb5e8 	:	val_out <= 4'h03e8;
         4'hb5e9 	:	val_out <= 4'h03e8;
         4'hb5ea 	:	val_out <= 4'h03e8;
         4'hb5eb 	:	val_out <= 4'h03e8;
         4'hb5f0 	:	val_out <= 4'h03e2;
         4'hb5f1 	:	val_out <= 4'h03e2;
         4'hb5f2 	:	val_out <= 4'h03e2;
         4'hb5f3 	:	val_out <= 4'h03e2;
         4'hb5f8 	:	val_out <= 4'h03dc;
         4'hb5f9 	:	val_out <= 4'h03dc;
         4'hb5fa 	:	val_out <= 4'h03dc;
         4'hb5fb 	:	val_out <= 4'h03dc;
         4'hb600 	:	val_out <= 4'h03d6;
         4'hb601 	:	val_out <= 4'h03d6;
         4'hb602 	:	val_out <= 4'h03d6;
         4'hb603 	:	val_out <= 4'h03d6;
         4'hb608 	:	val_out <= 4'h03cf;
         4'hb609 	:	val_out <= 4'h03cf;
         4'hb60a 	:	val_out <= 4'h03cf;
         4'hb60b 	:	val_out <= 4'h03cf;
         4'hb610 	:	val_out <= 4'h03c9;
         4'hb611 	:	val_out <= 4'h03c9;
         4'hb612 	:	val_out <= 4'h03c9;
         4'hb613 	:	val_out <= 4'h03c9;
         4'hb618 	:	val_out <= 4'h03c3;
         4'hb619 	:	val_out <= 4'h03c3;
         4'hb61a 	:	val_out <= 4'h03c3;
         4'hb61b 	:	val_out <= 4'h03c3;
         4'hb620 	:	val_out <= 4'h03bd;
         4'hb621 	:	val_out <= 4'h03bd;
         4'hb622 	:	val_out <= 4'h03bd;
         4'hb623 	:	val_out <= 4'h03bd;
         4'hb628 	:	val_out <= 4'h03b7;
         4'hb629 	:	val_out <= 4'h03b7;
         4'hb62a 	:	val_out <= 4'h03b7;
         4'hb62b 	:	val_out <= 4'h03b7;
         4'hb630 	:	val_out <= 4'h03b1;
         4'hb631 	:	val_out <= 4'h03b1;
         4'hb632 	:	val_out <= 4'h03b1;
         4'hb633 	:	val_out <= 4'h03b1;
         4'hb638 	:	val_out <= 4'h03ab;
         4'hb639 	:	val_out <= 4'h03ab;
         4'hb63a 	:	val_out <= 4'h03ab;
         4'hb63b 	:	val_out <= 4'h03ab;
         4'hb640 	:	val_out <= 4'h03a5;
         4'hb641 	:	val_out <= 4'h03a5;
         4'hb642 	:	val_out <= 4'h03a5;
         4'hb643 	:	val_out <= 4'h03a5;
         4'hb648 	:	val_out <= 4'h039f;
         4'hb649 	:	val_out <= 4'h039f;
         4'hb64a 	:	val_out <= 4'h039f;
         4'hb64b 	:	val_out <= 4'h039f;
         4'hb650 	:	val_out <= 4'h0399;
         4'hb651 	:	val_out <= 4'h0399;
         4'hb652 	:	val_out <= 4'h0399;
         4'hb653 	:	val_out <= 4'h0399;
         4'hb658 	:	val_out <= 4'h0393;
         4'hb659 	:	val_out <= 4'h0393;
         4'hb65a 	:	val_out <= 4'h0393;
         4'hb65b 	:	val_out <= 4'h0393;
         4'hb660 	:	val_out <= 4'h038e;
         4'hb661 	:	val_out <= 4'h038e;
         4'hb662 	:	val_out <= 4'h038e;
         4'hb663 	:	val_out <= 4'h038e;
         4'hb668 	:	val_out <= 4'h0388;
         4'hb669 	:	val_out <= 4'h0388;
         4'hb66a 	:	val_out <= 4'h0388;
         4'hb66b 	:	val_out <= 4'h0388;
         4'hb670 	:	val_out <= 4'h0382;
         4'hb671 	:	val_out <= 4'h0382;
         4'hb672 	:	val_out <= 4'h0382;
         4'hb673 	:	val_out <= 4'h0382;
         4'hb678 	:	val_out <= 4'h037c;
         4'hb679 	:	val_out <= 4'h037c;
         4'hb67a 	:	val_out <= 4'h037c;
         4'hb67b 	:	val_out <= 4'h037c;
         4'hb680 	:	val_out <= 4'h0376;
         4'hb681 	:	val_out <= 4'h0376;
         4'hb682 	:	val_out <= 4'h0376;
         4'hb683 	:	val_out <= 4'h0376;
         4'hb688 	:	val_out <= 4'h0370;
         4'hb689 	:	val_out <= 4'h0370;
         4'hb68a 	:	val_out <= 4'h0370;
         4'hb68b 	:	val_out <= 4'h0370;
         4'hb690 	:	val_out <= 4'h036b;
         4'hb691 	:	val_out <= 4'h036b;
         4'hb692 	:	val_out <= 4'h036b;
         4'hb693 	:	val_out <= 4'h036b;
         4'hb698 	:	val_out <= 4'h0365;
         4'hb699 	:	val_out <= 4'h0365;
         4'hb69a 	:	val_out <= 4'h0365;
         4'hb69b 	:	val_out <= 4'h0365;
         4'hb6a0 	:	val_out <= 4'h035f;
         4'hb6a1 	:	val_out <= 4'h035f;
         4'hb6a2 	:	val_out <= 4'h035f;
         4'hb6a3 	:	val_out <= 4'h035f;
         4'hb6a8 	:	val_out <= 4'h0359;
         4'hb6a9 	:	val_out <= 4'h0359;
         4'hb6aa 	:	val_out <= 4'h0359;
         4'hb6ab 	:	val_out <= 4'h0359;
         4'hb6b0 	:	val_out <= 4'h0354;
         4'hb6b1 	:	val_out <= 4'h0354;
         4'hb6b2 	:	val_out <= 4'h0354;
         4'hb6b3 	:	val_out <= 4'h0354;
         4'hb6b8 	:	val_out <= 4'h034e;
         4'hb6b9 	:	val_out <= 4'h034e;
         4'hb6ba 	:	val_out <= 4'h034e;
         4'hb6bb 	:	val_out <= 4'h034e;
         4'hb6c0 	:	val_out <= 4'h0348;
         4'hb6c1 	:	val_out <= 4'h0348;
         4'hb6c2 	:	val_out <= 4'h0348;
         4'hb6c3 	:	val_out <= 4'h0348;
         4'hb6c8 	:	val_out <= 4'h0343;
         4'hb6c9 	:	val_out <= 4'h0343;
         4'hb6ca 	:	val_out <= 4'h0343;
         4'hb6cb 	:	val_out <= 4'h0343;
         4'hb6d0 	:	val_out <= 4'h033d;
         4'hb6d1 	:	val_out <= 4'h033d;
         4'hb6d2 	:	val_out <= 4'h033d;
         4'hb6d3 	:	val_out <= 4'h033d;
         4'hb6d8 	:	val_out <= 4'h0337;
         4'hb6d9 	:	val_out <= 4'h0337;
         4'hb6da 	:	val_out <= 4'h0337;
         4'hb6db 	:	val_out <= 4'h0337;
         4'hb6e0 	:	val_out <= 4'h0332;
         4'hb6e1 	:	val_out <= 4'h0332;
         4'hb6e2 	:	val_out <= 4'h0332;
         4'hb6e3 	:	val_out <= 4'h0332;
         4'hb6e8 	:	val_out <= 4'h032c;
         4'hb6e9 	:	val_out <= 4'h032c;
         4'hb6ea 	:	val_out <= 4'h032c;
         4'hb6eb 	:	val_out <= 4'h032c;
         4'hb6f0 	:	val_out <= 4'h0327;
         4'hb6f1 	:	val_out <= 4'h0327;
         4'hb6f2 	:	val_out <= 4'h0327;
         4'hb6f3 	:	val_out <= 4'h0327;
         4'hb6f8 	:	val_out <= 4'h0321;
         4'hb6f9 	:	val_out <= 4'h0321;
         4'hb6fa 	:	val_out <= 4'h0321;
         4'hb6fb 	:	val_out <= 4'h0321;
         4'hb700 	:	val_out <= 4'h031c;
         4'hb701 	:	val_out <= 4'h031c;
         4'hb702 	:	val_out <= 4'h031c;
         4'hb703 	:	val_out <= 4'h031c;
         4'hb708 	:	val_out <= 4'h0316;
         4'hb709 	:	val_out <= 4'h0316;
         4'hb70a 	:	val_out <= 4'h0316;
         4'hb70b 	:	val_out <= 4'h0316;
         4'hb710 	:	val_out <= 4'h0311;
         4'hb711 	:	val_out <= 4'h0311;
         4'hb712 	:	val_out <= 4'h0311;
         4'hb713 	:	val_out <= 4'h0311;
         4'hb718 	:	val_out <= 4'h030b;
         4'hb719 	:	val_out <= 4'h030b;
         4'hb71a 	:	val_out <= 4'h030b;
         4'hb71b 	:	val_out <= 4'h030b;
         4'hb720 	:	val_out <= 4'h0306;
         4'hb721 	:	val_out <= 4'h0306;
         4'hb722 	:	val_out <= 4'h0306;
         4'hb723 	:	val_out <= 4'h0306;
         4'hb728 	:	val_out <= 4'h0300;
         4'hb729 	:	val_out <= 4'h0300;
         4'hb72a 	:	val_out <= 4'h0300;
         4'hb72b 	:	val_out <= 4'h0300;
         4'hb730 	:	val_out <= 4'h02fb;
         4'hb731 	:	val_out <= 4'h02fb;
         4'hb732 	:	val_out <= 4'h02fb;
         4'hb733 	:	val_out <= 4'h02fb;
         4'hb738 	:	val_out <= 4'h02f6;
         4'hb739 	:	val_out <= 4'h02f6;
         4'hb73a 	:	val_out <= 4'h02f6;
         4'hb73b 	:	val_out <= 4'h02f6;
         4'hb740 	:	val_out <= 4'h02f0;
         4'hb741 	:	val_out <= 4'h02f0;
         4'hb742 	:	val_out <= 4'h02f0;
         4'hb743 	:	val_out <= 4'h02f0;
         4'hb748 	:	val_out <= 4'h02eb;
         4'hb749 	:	val_out <= 4'h02eb;
         4'hb74a 	:	val_out <= 4'h02eb;
         4'hb74b 	:	val_out <= 4'h02eb;
         4'hb750 	:	val_out <= 4'h02e6;
         4'hb751 	:	val_out <= 4'h02e6;
         4'hb752 	:	val_out <= 4'h02e6;
         4'hb753 	:	val_out <= 4'h02e6;
         4'hb758 	:	val_out <= 4'h02e0;
         4'hb759 	:	val_out <= 4'h02e0;
         4'hb75a 	:	val_out <= 4'h02e0;
         4'hb75b 	:	val_out <= 4'h02e0;
         4'hb760 	:	val_out <= 4'h02db;
         4'hb761 	:	val_out <= 4'h02db;
         4'hb762 	:	val_out <= 4'h02db;
         4'hb763 	:	val_out <= 4'h02db;
         4'hb768 	:	val_out <= 4'h02d6;
         4'hb769 	:	val_out <= 4'h02d6;
         4'hb76a 	:	val_out <= 4'h02d6;
         4'hb76b 	:	val_out <= 4'h02d6;
         4'hb770 	:	val_out <= 4'h02d0;
         4'hb771 	:	val_out <= 4'h02d0;
         4'hb772 	:	val_out <= 4'h02d0;
         4'hb773 	:	val_out <= 4'h02d0;
         4'hb778 	:	val_out <= 4'h02cb;
         4'hb779 	:	val_out <= 4'h02cb;
         4'hb77a 	:	val_out <= 4'h02cb;
         4'hb77b 	:	val_out <= 4'h02cb;
         4'hb780 	:	val_out <= 4'h02c6;
         4'hb781 	:	val_out <= 4'h02c6;
         4'hb782 	:	val_out <= 4'h02c6;
         4'hb783 	:	val_out <= 4'h02c6;
         4'hb788 	:	val_out <= 4'h02c1;
         4'hb789 	:	val_out <= 4'h02c1;
         4'hb78a 	:	val_out <= 4'h02c1;
         4'hb78b 	:	val_out <= 4'h02c1;
         4'hb790 	:	val_out <= 4'h02bc;
         4'hb791 	:	val_out <= 4'h02bc;
         4'hb792 	:	val_out <= 4'h02bc;
         4'hb793 	:	val_out <= 4'h02bc;
         4'hb798 	:	val_out <= 4'h02b6;
         4'hb799 	:	val_out <= 4'h02b6;
         4'hb79a 	:	val_out <= 4'h02b6;
         4'hb79b 	:	val_out <= 4'h02b6;
         4'hb7a0 	:	val_out <= 4'h02b1;
         4'hb7a1 	:	val_out <= 4'h02b1;
         4'hb7a2 	:	val_out <= 4'h02b1;
         4'hb7a3 	:	val_out <= 4'h02b1;
         4'hb7a8 	:	val_out <= 4'h02ac;
         4'hb7a9 	:	val_out <= 4'h02ac;
         4'hb7aa 	:	val_out <= 4'h02ac;
         4'hb7ab 	:	val_out <= 4'h02ac;
         4'hb7b0 	:	val_out <= 4'h02a7;
         4'hb7b1 	:	val_out <= 4'h02a7;
         4'hb7b2 	:	val_out <= 4'h02a7;
         4'hb7b3 	:	val_out <= 4'h02a7;
         4'hb7b8 	:	val_out <= 4'h02a2;
         4'hb7b9 	:	val_out <= 4'h02a2;
         4'hb7ba 	:	val_out <= 4'h02a2;
         4'hb7bb 	:	val_out <= 4'h02a2;
         4'hb7c0 	:	val_out <= 4'h029d;
         4'hb7c1 	:	val_out <= 4'h029d;
         4'hb7c2 	:	val_out <= 4'h029d;
         4'hb7c3 	:	val_out <= 4'h029d;
         4'hb7c8 	:	val_out <= 4'h0298;
         4'hb7c9 	:	val_out <= 4'h0298;
         4'hb7ca 	:	val_out <= 4'h0298;
         4'hb7cb 	:	val_out <= 4'h0298;
         4'hb7d0 	:	val_out <= 4'h0293;
         4'hb7d1 	:	val_out <= 4'h0293;
         4'hb7d2 	:	val_out <= 4'h0293;
         4'hb7d3 	:	val_out <= 4'h0293;
         4'hb7d8 	:	val_out <= 4'h028e;
         4'hb7d9 	:	val_out <= 4'h028e;
         4'hb7da 	:	val_out <= 4'h028e;
         4'hb7db 	:	val_out <= 4'h028e;
         4'hb7e0 	:	val_out <= 4'h0289;
         4'hb7e1 	:	val_out <= 4'h0289;
         4'hb7e2 	:	val_out <= 4'h0289;
         4'hb7e3 	:	val_out <= 4'h0289;
         4'hb7e8 	:	val_out <= 4'h0284;
         4'hb7e9 	:	val_out <= 4'h0284;
         4'hb7ea 	:	val_out <= 4'h0284;
         4'hb7eb 	:	val_out <= 4'h0284;
         4'hb7f0 	:	val_out <= 4'h027f;
         4'hb7f1 	:	val_out <= 4'h027f;
         4'hb7f2 	:	val_out <= 4'h027f;
         4'hb7f3 	:	val_out <= 4'h027f;
         4'hb7f8 	:	val_out <= 4'h027a;
         4'hb7f9 	:	val_out <= 4'h027a;
         4'hb7fa 	:	val_out <= 4'h027a;
         4'hb7fb 	:	val_out <= 4'h027a;
         4'hb800 	:	val_out <= 4'h0275;
         4'hb801 	:	val_out <= 4'h0275;
         4'hb802 	:	val_out <= 4'h0275;
         4'hb803 	:	val_out <= 4'h0275;
         4'hb808 	:	val_out <= 4'h0270;
         4'hb809 	:	val_out <= 4'h0270;
         4'hb80a 	:	val_out <= 4'h0270;
         4'hb80b 	:	val_out <= 4'h0270;
         4'hb810 	:	val_out <= 4'h026b;
         4'hb811 	:	val_out <= 4'h026b;
         4'hb812 	:	val_out <= 4'h026b;
         4'hb813 	:	val_out <= 4'h026b;
         4'hb818 	:	val_out <= 4'h0267;
         4'hb819 	:	val_out <= 4'h0267;
         4'hb81a 	:	val_out <= 4'h0267;
         4'hb81b 	:	val_out <= 4'h0267;
         4'hb820 	:	val_out <= 4'h0262;
         4'hb821 	:	val_out <= 4'h0262;
         4'hb822 	:	val_out <= 4'h0262;
         4'hb823 	:	val_out <= 4'h0262;
         4'hb828 	:	val_out <= 4'h025d;
         4'hb829 	:	val_out <= 4'h025d;
         4'hb82a 	:	val_out <= 4'h025d;
         4'hb82b 	:	val_out <= 4'h025d;
         4'hb830 	:	val_out <= 4'h0258;
         4'hb831 	:	val_out <= 4'h0258;
         4'hb832 	:	val_out <= 4'h0258;
         4'hb833 	:	val_out <= 4'h0258;
         4'hb838 	:	val_out <= 4'h0253;
         4'hb839 	:	val_out <= 4'h0253;
         4'hb83a 	:	val_out <= 4'h0253;
         4'hb83b 	:	val_out <= 4'h0253;
         4'hb840 	:	val_out <= 4'h024f;
         4'hb841 	:	val_out <= 4'h024f;
         4'hb842 	:	val_out <= 4'h024f;
         4'hb843 	:	val_out <= 4'h024f;
         4'hb848 	:	val_out <= 4'h024a;
         4'hb849 	:	val_out <= 4'h024a;
         4'hb84a 	:	val_out <= 4'h024a;
         4'hb84b 	:	val_out <= 4'h024a;
         4'hb850 	:	val_out <= 4'h0245;
         4'hb851 	:	val_out <= 4'h0245;
         4'hb852 	:	val_out <= 4'h0245;
         4'hb853 	:	val_out <= 4'h0245;
         4'hb858 	:	val_out <= 4'h0240;
         4'hb859 	:	val_out <= 4'h0240;
         4'hb85a 	:	val_out <= 4'h0240;
         4'hb85b 	:	val_out <= 4'h0240;
         4'hb860 	:	val_out <= 4'h023c;
         4'hb861 	:	val_out <= 4'h023c;
         4'hb862 	:	val_out <= 4'h023c;
         4'hb863 	:	val_out <= 4'h023c;
         4'hb868 	:	val_out <= 4'h0237;
         4'hb869 	:	val_out <= 4'h0237;
         4'hb86a 	:	val_out <= 4'h0237;
         4'hb86b 	:	val_out <= 4'h0237;
         4'hb870 	:	val_out <= 4'h0232;
         4'hb871 	:	val_out <= 4'h0232;
         4'hb872 	:	val_out <= 4'h0232;
         4'hb873 	:	val_out <= 4'h0232;
         4'hb878 	:	val_out <= 4'h022e;
         4'hb879 	:	val_out <= 4'h022e;
         4'hb87a 	:	val_out <= 4'h022e;
         4'hb87b 	:	val_out <= 4'h022e;
         4'hb880 	:	val_out <= 4'h0229;
         4'hb881 	:	val_out <= 4'h0229;
         4'hb882 	:	val_out <= 4'h0229;
         4'hb883 	:	val_out <= 4'h0229;
         4'hb888 	:	val_out <= 4'h0225;
         4'hb889 	:	val_out <= 4'h0225;
         4'hb88a 	:	val_out <= 4'h0225;
         4'hb88b 	:	val_out <= 4'h0225;
         4'hb890 	:	val_out <= 4'h0220;
         4'hb891 	:	val_out <= 4'h0220;
         4'hb892 	:	val_out <= 4'h0220;
         4'hb893 	:	val_out <= 4'h0220;
         4'hb898 	:	val_out <= 4'h021b;
         4'hb899 	:	val_out <= 4'h021b;
         4'hb89a 	:	val_out <= 4'h021b;
         4'hb89b 	:	val_out <= 4'h021b;
         4'hb8a0 	:	val_out <= 4'h0217;
         4'hb8a1 	:	val_out <= 4'h0217;
         4'hb8a2 	:	val_out <= 4'h0217;
         4'hb8a3 	:	val_out <= 4'h0217;
         4'hb8a8 	:	val_out <= 4'h0212;
         4'hb8a9 	:	val_out <= 4'h0212;
         4'hb8aa 	:	val_out <= 4'h0212;
         4'hb8ab 	:	val_out <= 4'h0212;
         4'hb8b0 	:	val_out <= 4'h020e;
         4'hb8b1 	:	val_out <= 4'h020e;
         4'hb8b2 	:	val_out <= 4'h020e;
         4'hb8b3 	:	val_out <= 4'h020e;
         4'hb8b8 	:	val_out <= 4'h0209;
         4'hb8b9 	:	val_out <= 4'h0209;
         4'hb8ba 	:	val_out <= 4'h0209;
         4'hb8bb 	:	val_out <= 4'h0209;
         4'hb8c0 	:	val_out <= 4'h0205;
         4'hb8c1 	:	val_out <= 4'h0205;
         4'hb8c2 	:	val_out <= 4'h0205;
         4'hb8c3 	:	val_out <= 4'h0205;
         4'hb8c8 	:	val_out <= 4'h0200;
         4'hb8c9 	:	val_out <= 4'h0200;
         4'hb8ca 	:	val_out <= 4'h0200;
         4'hb8cb 	:	val_out <= 4'h0200;
         4'hb8d0 	:	val_out <= 4'h01fc;
         4'hb8d1 	:	val_out <= 4'h01fc;
         4'hb8d2 	:	val_out <= 4'h01fc;
         4'hb8d3 	:	val_out <= 4'h01fc;
         4'hb8d8 	:	val_out <= 4'h01f8;
         4'hb8d9 	:	val_out <= 4'h01f8;
         4'hb8da 	:	val_out <= 4'h01f8;
         4'hb8db 	:	val_out <= 4'h01f8;
         4'hb8e0 	:	val_out <= 4'h01f3;
         4'hb8e1 	:	val_out <= 4'h01f3;
         4'hb8e2 	:	val_out <= 4'h01f3;
         4'hb8e3 	:	val_out <= 4'h01f3;
         4'hb8e8 	:	val_out <= 4'h01ef;
         4'hb8e9 	:	val_out <= 4'h01ef;
         4'hb8ea 	:	val_out <= 4'h01ef;
         4'hb8eb 	:	val_out <= 4'h01ef;
         4'hb8f0 	:	val_out <= 4'h01eb;
         4'hb8f1 	:	val_out <= 4'h01eb;
         4'hb8f2 	:	val_out <= 4'h01eb;
         4'hb8f3 	:	val_out <= 4'h01eb;
         4'hb8f8 	:	val_out <= 4'h01e6;
         4'hb8f9 	:	val_out <= 4'h01e6;
         4'hb8fa 	:	val_out <= 4'h01e6;
         4'hb8fb 	:	val_out <= 4'h01e6;
         4'hb900 	:	val_out <= 4'h01e2;
         4'hb901 	:	val_out <= 4'h01e2;
         4'hb902 	:	val_out <= 4'h01e2;
         4'hb903 	:	val_out <= 4'h01e2;
         4'hb908 	:	val_out <= 4'h01de;
         4'hb909 	:	val_out <= 4'h01de;
         4'hb90a 	:	val_out <= 4'h01de;
         4'hb90b 	:	val_out <= 4'h01de;
         4'hb910 	:	val_out <= 4'h01d9;
         4'hb911 	:	val_out <= 4'h01d9;
         4'hb912 	:	val_out <= 4'h01d9;
         4'hb913 	:	val_out <= 4'h01d9;
         4'hb918 	:	val_out <= 4'h01d5;
         4'hb919 	:	val_out <= 4'h01d5;
         4'hb91a 	:	val_out <= 4'h01d5;
         4'hb91b 	:	val_out <= 4'h01d5;
         4'hb920 	:	val_out <= 4'h01d1;
         4'hb921 	:	val_out <= 4'h01d1;
         4'hb922 	:	val_out <= 4'h01d1;
         4'hb923 	:	val_out <= 4'h01d1;
         4'hb928 	:	val_out <= 4'h01cd;
         4'hb929 	:	val_out <= 4'h01cd;
         4'hb92a 	:	val_out <= 4'h01cd;
         4'hb92b 	:	val_out <= 4'h01cd;
         4'hb930 	:	val_out <= 4'h01c8;
         4'hb931 	:	val_out <= 4'h01c8;
         4'hb932 	:	val_out <= 4'h01c8;
         4'hb933 	:	val_out <= 4'h01c8;
         4'hb938 	:	val_out <= 4'h01c4;
         4'hb939 	:	val_out <= 4'h01c4;
         4'hb93a 	:	val_out <= 4'h01c4;
         4'hb93b 	:	val_out <= 4'h01c4;
         4'hb940 	:	val_out <= 4'h01c0;
         4'hb941 	:	val_out <= 4'h01c0;
         4'hb942 	:	val_out <= 4'h01c0;
         4'hb943 	:	val_out <= 4'h01c0;
         4'hb948 	:	val_out <= 4'h01bc;
         4'hb949 	:	val_out <= 4'h01bc;
         4'hb94a 	:	val_out <= 4'h01bc;
         4'hb94b 	:	val_out <= 4'h01bc;
         4'hb950 	:	val_out <= 4'h01b8;
         4'hb951 	:	val_out <= 4'h01b8;
         4'hb952 	:	val_out <= 4'h01b8;
         4'hb953 	:	val_out <= 4'h01b8;
         4'hb958 	:	val_out <= 4'h01b4;
         4'hb959 	:	val_out <= 4'h01b4;
         4'hb95a 	:	val_out <= 4'h01b4;
         4'hb95b 	:	val_out <= 4'h01b4;
         4'hb960 	:	val_out <= 4'h01b0;
         4'hb961 	:	val_out <= 4'h01b0;
         4'hb962 	:	val_out <= 4'h01b0;
         4'hb963 	:	val_out <= 4'h01b0;
         4'hb968 	:	val_out <= 4'h01ac;
         4'hb969 	:	val_out <= 4'h01ac;
         4'hb96a 	:	val_out <= 4'h01ac;
         4'hb96b 	:	val_out <= 4'h01ac;
         4'hb970 	:	val_out <= 4'h01a8;
         4'hb971 	:	val_out <= 4'h01a8;
         4'hb972 	:	val_out <= 4'h01a8;
         4'hb973 	:	val_out <= 4'h01a8;
         4'hb978 	:	val_out <= 4'h01a4;
         4'hb979 	:	val_out <= 4'h01a4;
         4'hb97a 	:	val_out <= 4'h01a4;
         4'hb97b 	:	val_out <= 4'h01a4;
         4'hb980 	:	val_out <= 4'h01a0;
         4'hb981 	:	val_out <= 4'h01a0;
         4'hb982 	:	val_out <= 4'h01a0;
         4'hb983 	:	val_out <= 4'h01a0;
         4'hb988 	:	val_out <= 4'h019c;
         4'hb989 	:	val_out <= 4'h019c;
         4'hb98a 	:	val_out <= 4'h019c;
         4'hb98b 	:	val_out <= 4'h019c;
         4'hb990 	:	val_out <= 4'h0198;
         4'hb991 	:	val_out <= 4'h0198;
         4'hb992 	:	val_out <= 4'h0198;
         4'hb993 	:	val_out <= 4'h0198;
         4'hb998 	:	val_out <= 4'h0194;
         4'hb999 	:	val_out <= 4'h0194;
         4'hb99a 	:	val_out <= 4'h0194;
         4'hb99b 	:	val_out <= 4'h0194;
         4'hb9a0 	:	val_out <= 4'h0190;
         4'hb9a1 	:	val_out <= 4'h0190;
         4'hb9a2 	:	val_out <= 4'h0190;
         4'hb9a3 	:	val_out <= 4'h0190;
         4'hb9a8 	:	val_out <= 4'h018c;
         4'hb9a9 	:	val_out <= 4'h018c;
         4'hb9aa 	:	val_out <= 4'h018c;
         4'hb9ab 	:	val_out <= 4'h018c;
         4'hb9b0 	:	val_out <= 4'h0188;
         4'hb9b1 	:	val_out <= 4'h0188;
         4'hb9b2 	:	val_out <= 4'h0188;
         4'hb9b3 	:	val_out <= 4'h0188;
         4'hb9b8 	:	val_out <= 4'h0184;
         4'hb9b9 	:	val_out <= 4'h0184;
         4'hb9ba 	:	val_out <= 4'h0184;
         4'hb9bb 	:	val_out <= 4'h0184;
         4'hb9c0 	:	val_out <= 4'h0180;
         4'hb9c1 	:	val_out <= 4'h0180;
         4'hb9c2 	:	val_out <= 4'h0180;
         4'hb9c3 	:	val_out <= 4'h0180;
         4'hb9c8 	:	val_out <= 4'h017c;
         4'hb9c9 	:	val_out <= 4'h017c;
         4'hb9ca 	:	val_out <= 4'h017c;
         4'hb9cb 	:	val_out <= 4'h017c;
         4'hb9d0 	:	val_out <= 4'h0179;
         4'hb9d1 	:	val_out <= 4'h0179;
         4'hb9d2 	:	val_out <= 4'h0179;
         4'hb9d3 	:	val_out <= 4'h0179;
         4'hb9d8 	:	val_out <= 4'h0175;
         4'hb9d9 	:	val_out <= 4'h0175;
         4'hb9da 	:	val_out <= 4'h0175;
         4'hb9db 	:	val_out <= 4'h0175;
         4'hb9e0 	:	val_out <= 4'h0171;
         4'hb9e1 	:	val_out <= 4'h0171;
         4'hb9e2 	:	val_out <= 4'h0171;
         4'hb9e3 	:	val_out <= 4'h0171;
         4'hb9e8 	:	val_out <= 4'h016d;
         4'hb9e9 	:	val_out <= 4'h016d;
         4'hb9ea 	:	val_out <= 4'h016d;
         4'hb9eb 	:	val_out <= 4'h016d;
         4'hb9f0 	:	val_out <= 4'h016a;
         4'hb9f1 	:	val_out <= 4'h016a;
         4'hb9f2 	:	val_out <= 4'h016a;
         4'hb9f3 	:	val_out <= 4'h016a;
         4'hb9f8 	:	val_out <= 4'h0166;
         4'hb9f9 	:	val_out <= 4'h0166;
         4'hb9fa 	:	val_out <= 4'h0166;
         4'hb9fb 	:	val_out <= 4'h0166;
         4'hba00 	:	val_out <= 4'h0162;
         4'hba01 	:	val_out <= 4'h0162;
         4'hba02 	:	val_out <= 4'h0162;
         4'hba03 	:	val_out <= 4'h0162;
         4'hba08 	:	val_out <= 4'h015e;
         4'hba09 	:	val_out <= 4'h015e;
         4'hba0a 	:	val_out <= 4'h015e;
         4'hba0b 	:	val_out <= 4'h015e;
         4'hba10 	:	val_out <= 4'h015b;
         4'hba11 	:	val_out <= 4'h015b;
         4'hba12 	:	val_out <= 4'h015b;
         4'hba13 	:	val_out <= 4'h015b;
         4'hba18 	:	val_out <= 4'h0157;
         4'hba19 	:	val_out <= 4'h0157;
         4'hba1a 	:	val_out <= 4'h0157;
         4'hba1b 	:	val_out <= 4'h0157;
         4'hba20 	:	val_out <= 4'h0154;
         4'hba21 	:	val_out <= 4'h0154;
         4'hba22 	:	val_out <= 4'h0154;
         4'hba23 	:	val_out <= 4'h0154;
         4'hba28 	:	val_out <= 4'h0150;
         4'hba29 	:	val_out <= 4'h0150;
         4'hba2a 	:	val_out <= 4'h0150;
         4'hba2b 	:	val_out <= 4'h0150;
         4'hba30 	:	val_out <= 4'h014c;
         4'hba31 	:	val_out <= 4'h014c;
         4'hba32 	:	val_out <= 4'h014c;
         4'hba33 	:	val_out <= 4'h014c;
         4'hba38 	:	val_out <= 4'h0149;
         4'hba39 	:	val_out <= 4'h0149;
         4'hba3a 	:	val_out <= 4'h0149;
         4'hba3b 	:	val_out <= 4'h0149;
         4'hba40 	:	val_out <= 4'h0145;
         4'hba41 	:	val_out <= 4'h0145;
         4'hba42 	:	val_out <= 4'h0145;
         4'hba43 	:	val_out <= 4'h0145;
         4'hba48 	:	val_out <= 4'h0142;
         4'hba49 	:	val_out <= 4'h0142;
         4'hba4a 	:	val_out <= 4'h0142;
         4'hba4b 	:	val_out <= 4'h0142;
         4'hba50 	:	val_out <= 4'h013e;
         4'hba51 	:	val_out <= 4'h013e;
         4'hba52 	:	val_out <= 4'h013e;
         4'hba53 	:	val_out <= 4'h013e;
         4'hba58 	:	val_out <= 4'h013b;
         4'hba59 	:	val_out <= 4'h013b;
         4'hba5a 	:	val_out <= 4'h013b;
         4'hba5b 	:	val_out <= 4'h013b;
         4'hba60 	:	val_out <= 4'h0137;
         4'hba61 	:	val_out <= 4'h0137;
         4'hba62 	:	val_out <= 4'h0137;
         4'hba63 	:	val_out <= 4'h0137;
         4'hba68 	:	val_out <= 4'h0134;
         4'hba69 	:	val_out <= 4'h0134;
         4'hba6a 	:	val_out <= 4'h0134;
         4'hba6b 	:	val_out <= 4'h0134;
         4'hba70 	:	val_out <= 4'h0130;
         4'hba71 	:	val_out <= 4'h0130;
         4'hba72 	:	val_out <= 4'h0130;
         4'hba73 	:	val_out <= 4'h0130;
         4'hba78 	:	val_out <= 4'h012d;
         4'hba79 	:	val_out <= 4'h012d;
         4'hba7a 	:	val_out <= 4'h012d;
         4'hba7b 	:	val_out <= 4'h012d;
         4'hba80 	:	val_out <= 4'h012a;
         4'hba81 	:	val_out <= 4'h012a;
         4'hba82 	:	val_out <= 4'h012a;
         4'hba83 	:	val_out <= 4'h012a;
         4'hba88 	:	val_out <= 4'h0126;
         4'hba89 	:	val_out <= 4'h0126;
         4'hba8a 	:	val_out <= 4'h0126;
         4'hba8b 	:	val_out <= 4'h0126;
         4'hba90 	:	val_out <= 4'h0123;
         4'hba91 	:	val_out <= 4'h0123;
         4'hba92 	:	val_out <= 4'h0123;
         4'hba93 	:	val_out <= 4'h0123;
         4'hba98 	:	val_out <= 4'h0120;
         4'hba99 	:	val_out <= 4'h0120;
         4'hba9a 	:	val_out <= 4'h0120;
         4'hba9b 	:	val_out <= 4'h0120;
         4'hbaa0 	:	val_out <= 4'h011c;
         4'hbaa1 	:	val_out <= 4'h011c;
         4'hbaa2 	:	val_out <= 4'h011c;
         4'hbaa3 	:	val_out <= 4'h011c;
         4'hbaa8 	:	val_out <= 4'h0119;
         4'hbaa9 	:	val_out <= 4'h0119;
         4'hbaaa 	:	val_out <= 4'h0119;
         4'hbaab 	:	val_out <= 4'h0119;
         4'hbab0 	:	val_out <= 4'h0116;
         4'hbab1 	:	val_out <= 4'h0116;
         4'hbab2 	:	val_out <= 4'h0116;
         4'hbab3 	:	val_out <= 4'h0116;
         4'hbab8 	:	val_out <= 4'h0112;
         4'hbab9 	:	val_out <= 4'h0112;
         4'hbaba 	:	val_out <= 4'h0112;
         4'hbabb 	:	val_out <= 4'h0112;
         4'hbac0 	:	val_out <= 4'h010f;
         4'hbac1 	:	val_out <= 4'h010f;
         4'hbac2 	:	val_out <= 4'h010f;
         4'hbac3 	:	val_out <= 4'h010f;
         4'hbac8 	:	val_out <= 4'h010c;
         4'hbac9 	:	val_out <= 4'h010c;
         4'hbaca 	:	val_out <= 4'h010c;
         4'hbacb 	:	val_out <= 4'h010c;
         4'hbad0 	:	val_out <= 4'h0109;
         4'hbad1 	:	val_out <= 4'h0109;
         4'hbad2 	:	val_out <= 4'h0109;
         4'hbad3 	:	val_out <= 4'h0109;
         4'hbad8 	:	val_out <= 4'h0106;
         4'hbad9 	:	val_out <= 4'h0106;
         4'hbada 	:	val_out <= 4'h0106;
         4'hbadb 	:	val_out <= 4'h0106;
         4'hbae0 	:	val_out <= 4'h0102;
         4'hbae1 	:	val_out <= 4'h0102;
         4'hbae2 	:	val_out <= 4'h0102;
         4'hbae3 	:	val_out <= 4'h0102;
         4'hbae8 	:	val_out <= 4'h00ff;
         4'hbae9 	:	val_out <= 4'h00ff;
         4'hbaea 	:	val_out <= 4'h00ff;
         4'hbaeb 	:	val_out <= 4'h00ff;
         4'hbaf0 	:	val_out <= 4'h00fc;
         4'hbaf1 	:	val_out <= 4'h00fc;
         4'hbaf2 	:	val_out <= 4'h00fc;
         4'hbaf3 	:	val_out <= 4'h00fc;
         4'hbaf8 	:	val_out <= 4'h00f9;
         4'hbaf9 	:	val_out <= 4'h00f9;
         4'hbafa 	:	val_out <= 4'h00f9;
         4'hbafb 	:	val_out <= 4'h00f9;
         4'hbb00 	:	val_out <= 4'h00f6;
         4'hbb01 	:	val_out <= 4'h00f6;
         4'hbb02 	:	val_out <= 4'h00f6;
         4'hbb03 	:	val_out <= 4'h00f6;
         4'hbb08 	:	val_out <= 4'h00f3;
         4'hbb09 	:	val_out <= 4'h00f3;
         4'hbb0a 	:	val_out <= 4'h00f3;
         4'hbb0b 	:	val_out <= 4'h00f3;
         4'hbb10 	:	val_out <= 4'h00f0;
         4'hbb11 	:	val_out <= 4'h00f0;
         4'hbb12 	:	val_out <= 4'h00f0;
         4'hbb13 	:	val_out <= 4'h00f0;
         4'hbb18 	:	val_out <= 4'h00ed;
         4'hbb19 	:	val_out <= 4'h00ed;
         4'hbb1a 	:	val_out <= 4'h00ed;
         4'hbb1b 	:	val_out <= 4'h00ed;
         4'hbb20 	:	val_out <= 4'h00ea;
         4'hbb21 	:	val_out <= 4'h00ea;
         4'hbb22 	:	val_out <= 4'h00ea;
         4'hbb23 	:	val_out <= 4'h00ea;
         4'hbb28 	:	val_out <= 4'h00e7;
         4'hbb29 	:	val_out <= 4'h00e7;
         4'hbb2a 	:	val_out <= 4'h00e7;
         4'hbb2b 	:	val_out <= 4'h00e7;
         4'hbb30 	:	val_out <= 4'h00e4;
         4'hbb31 	:	val_out <= 4'h00e4;
         4'hbb32 	:	val_out <= 4'h00e4;
         4'hbb33 	:	val_out <= 4'h00e4;
         4'hbb38 	:	val_out <= 4'h00e1;
         4'hbb39 	:	val_out <= 4'h00e1;
         4'hbb3a 	:	val_out <= 4'h00e1;
         4'hbb3b 	:	val_out <= 4'h00e1;
         4'hbb40 	:	val_out <= 4'h00de;
         4'hbb41 	:	val_out <= 4'h00de;
         4'hbb42 	:	val_out <= 4'h00de;
         4'hbb43 	:	val_out <= 4'h00de;
         4'hbb48 	:	val_out <= 4'h00db;
         4'hbb49 	:	val_out <= 4'h00db;
         4'hbb4a 	:	val_out <= 4'h00db;
         4'hbb4b 	:	val_out <= 4'h00db;
         4'hbb50 	:	val_out <= 4'h00d8;
         4'hbb51 	:	val_out <= 4'h00d8;
         4'hbb52 	:	val_out <= 4'h00d8;
         4'hbb53 	:	val_out <= 4'h00d8;
         4'hbb58 	:	val_out <= 4'h00d5;
         4'hbb59 	:	val_out <= 4'h00d5;
         4'hbb5a 	:	val_out <= 4'h00d5;
         4'hbb5b 	:	val_out <= 4'h00d5;
         4'hbb60 	:	val_out <= 4'h00d2;
         4'hbb61 	:	val_out <= 4'h00d2;
         4'hbb62 	:	val_out <= 4'h00d2;
         4'hbb63 	:	val_out <= 4'h00d2;
         4'hbb68 	:	val_out <= 4'h00d0;
         4'hbb69 	:	val_out <= 4'h00d0;
         4'hbb6a 	:	val_out <= 4'h00d0;
         4'hbb6b 	:	val_out <= 4'h00d0;
         4'hbb70 	:	val_out <= 4'h00cd;
         4'hbb71 	:	val_out <= 4'h00cd;
         4'hbb72 	:	val_out <= 4'h00cd;
         4'hbb73 	:	val_out <= 4'h00cd;
         4'hbb78 	:	val_out <= 4'h00ca;
         4'hbb79 	:	val_out <= 4'h00ca;
         4'hbb7a 	:	val_out <= 4'h00ca;
         4'hbb7b 	:	val_out <= 4'h00ca;
         4'hbb80 	:	val_out <= 4'h00c7;
         4'hbb81 	:	val_out <= 4'h00c7;
         4'hbb82 	:	val_out <= 4'h00c7;
         4'hbb83 	:	val_out <= 4'h00c7;
         4'hbb88 	:	val_out <= 4'h00c4;
         4'hbb89 	:	val_out <= 4'h00c4;
         4'hbb8a 	:	val_out <= 4'h00c4;
         4'hbb8b 	:	val_out <= 4'h00c4;
         4'hbb90 	:	val_out <= 4'h00c2;
         4'hbb91 	:	val_out <= 4'h00c2;
         4'hbb92 	:	val_out <= 4'h00c2;
         4'hbb93 	:	val_out <= 4'h00c2;
         4'hbb98 	:	val_out <= 4'h00bf;
         4'hbb99 	:	val_out <= 4'h00bf;
         4'hbb9a 	:	val_out <= 4'h00bf;
         4'hbb9b 	:	val_out <= 4'h00bf;
         4'hbba0 	:	val_out <= 4'h00bc;
         4'hbba1 	:	val_out <= 4'h00bc;
         4'hbba2 	:	val_out <= 4'h00bc;
         4'hbba3 	:	val_out <= 4'h00bc;
         4'hbba8 	:	val_out <= 4'h00ba;
         4'hbba9 	:	val_out <= 4'h00ba;
         4'hbbaa 	:	val_out <= 4'h00ba;
         4'hbbab 	:	val_out <= 4'h00ba;
         4'hbbb0 	:	val_out <= 4'h00b7;
         4'hbbb1 	:	val_out <= 4'h00b7;
         4'hbbb2 	:	val_out <= 4'h00b7;
         4'hbbb3 	:	val_out <= 4'h00b7;
         4'hbbb8 	:	val_out <= 4'h00b4;
         4'hbbb9 	:	val_out <= 4'h00b4;
         4'hbbba 	:	val_out <= 4'h00b4;
         4'hbbbb 	:	val_out <= 4'h00b4;
         4'hbbc0 	:	val_out <= 4'h00b2;
         4'hbbc1 	:	val_out <= 4'h00b2;
         4'hbbc2 	:	val_out <= 4'h00b2;
         4'hbbc3 	:	val_out <= 4'h00b2;
         4'hbbc8 	:	val_out <= 4'h00af;
         4'hbbc9 	:	val_out <= 4'h00af;
         4'hbbca 	:	val_out <= 4'h00af;
         4'hbbcb 	:	val_out <= 4'h00af;
         4'hbbd0 	:	val_out <= 4'h00ac;
         4'hbbd1 	:	val_out <= 4'h00ac;
         4'hbbd2 	:	val_out <= 4'h00ac;
         4'hbbd3 	:	val_out <= 4'h00ac;
         4'hbbd8 	:	val_out <= 4'h00aa;
         4'hbbd9 	:	val_out <= 4'h00aa;
         4'hbbda 	:	val_out <= 4'h00aa;
         4'hbbdb 	:	val_out <= 4'h00aa;
         4'hbbe0 	:	val_out <= 4'h00a7;
         4'hbbe1 	:	val_out <= 4'h00a7;
         4'hbbe2 	:	val_out <= 4'h00a7;
         4'hbbe3 	:	val_out <= 4'h00a7;
         4'hbbe8 	:	val_out <= 4'h00a5;
         4'hbbe9 	:	val_out <= 4'h00a5;
         4'hbbea 	:	val_out <= 4'h00a5;
         4'hbbeb 	:	val_out <= 4'h00a5;
         4'hbbf0 	:	val_out <= 4'h00a2;
         4'hbbf1 	:	val_out <= 4'h00a2;
         4'hbbf2 	:	val_out <= 4'h00a2;
         4'hbbf3 	:	val_out <= 4'h00a2;
         4'hbbf8 	:	val_out <= 4'h00a0;
         4'hbbf9 	:	val_out <= 4'h00a0;
         4'hbbfa 	:	val_out <= 4'h00a0;
         4'hbbfb 	:	val_out <= 4'h00a0;
         4'hbc00 	:	val_out <= 4'h009d;
         4'hbc01 	:	val_out <= 4'h009d;
         4'hbc02 	:	val_out <= 4'h009d;
         4'hbc03 	:	val_out <= 4'h009d;
         4'hbc08 	:	val_out <= 4'h009b;
         4'hbc09 	:	val_out <= 4'h009b;
         4'hbc0a 	:	val_out <= 4'h009b;
         4'hbc0b 	:	val_out <= 4'h009b;
         4'hbc10 	:	val_out <= 4'h0098;
         4'hbc11 	:	val_out <= 4'h0098;
         4'hbc12 	:	val_out <= 4'h0098;
         4'hbc13 	:	val_out <= 4'h0098;
         4'hbc18 	:	val_out <= 4'h0096;
         4'hbc19 	:	val_out <= 4'h0096;
         4'hbc1a 	:	val_out <= 4'h0096;
         4'hbc1b 	:	val_out <= 4'h0096;
         4'hbc20 	:	val_out <= 4'h0094;
         4'hbc21 	:	val_out <= 4'h0094;
         4'hbc22 	:	val_out <= 4'h0094;
         4'hbc23 	:	val_out <= 4'h0094;
         4'hbc28 	:	val_out <= 4'h0091;
         4'hbc29 	:	val_out <= 4'h0091;
         4'hbc2a 	:	val_out <= 4'h0091;
         4'hbc2b 	:	val_out <= 4'h0091;
         4'hbc30 	:	val_out <= 4'h008f;
         4'hbc31 	:	val_out <= 4'h008f;
         4'hbc32 	:	val_out <= 4'h008f;
         4'hbc33 	:	val_out <= 4'h008f;
         4'hbc38 	:	val_out <= 4'h008d;
         4'hbc39 	:	val_out <= 4'h008d;
         4'hbc3a 	:	val_out <= 4'h008d;
         4'hbc3b 	:	val_out <= 4'h008d;
         4'hbc40 	:	val_out <= 4'h008a;
         4'hbc41 	:	val_out <= 4'h008a;
         4'hbc42 	:	val_out <= 4'h008a;
         4'hbc43 	:	val_out <= 4'h008a;
         4'hbc48 	:	val_out <= 4'h0088;
         4'hbc49 	:	val_out <= 4'h0088;
         4'hbc4a 	:	val_out <= 4'h0088;
         4'hbc4b 	:	val_out <= 4'h0088;
         4'hbc50 	:	val_out <= 4'h0086;
         4'hbc51 	:	val_out <= 4'h0086;
         4'hbc52 	:	val_out <= 4'h0086;
         4'hbc53 	:	val_out <= 4'h0086;
         4'hbc58 	:	val_out <= 4'h0083;
         4'hbc59 	:	val_out <= 4'h0083;
         4'hbc5a 	:	val_out <= 4'h0083;
         4'hbc5b 	:	val_out <= 4'h0083;
         4'hbc60 	:	val_out <= 4'h0081;
         4'hbc61 	:	val_out <= 4'h0081;
         4'hbc62 	:	val_out <= 4'h0081;
         4'hbc63 	:	val_out <= 4'h0081;
         4'hbc68 	:	val_out <= 4'h007f;
         4'hbc69 	:	val_out <= 4'h007f;
         4'hbc6a 	:	val_out <= 4'h007f;
         4'hbc6b 	:	val_out <= 4'h007f;
         4'hbc70 	:	val_out <= 4'h007d;
         4'hbc71 	:	val_out <= 4'h007d;
         4'hbc72 	:	val_out <= 4'h007d;
         4'hbc73 	:	val_out <= 4'h007d;
         4'hbc78 	:	val_out <= 4'h007a;
         4'hbc79 	:	val_out <= 4'h007a;
         4'hbc7a 	:	val_out <= 4'h007a;
         4'hbc7b 	:	val_out <= 4'h007a;
         4'hbc80 	:	val_out <= 4'h0078;
         4'hbc81 	:	val_out <= 4'h0078;
         4'hbc82 	:	val_out <= 4'h0078;
         4'hbc83 	:	val_out <= 4'h0078;
         4'hbc88 	:	val_out <= 4'h0076;
         4'hbc89 	:	val_out <= 4'h0076;
         4'hbc8a 	:	val_out <= 4'h0076;
         4'hbc8b 	:	val_out <= 4'h0076;
         4'hbc90 	:	val_out <= 4'h0074;
         4'hbc91 	:	val_out <= 4'h0074;
         4'hbc92 	:	val_out <= 4'h0074;
         4'hbc93 	:	val_out <= 4'h0074;
         4'hbc98 	:	val_out <= 4'h0072;
         4'hbc99 	:	val_out <= 4'h0072;
         4'hbc9a 	:	val_out <= 4'h0072;
         4'hbc9b 	:	val_out <= 4'h0072;
         4'hbca0 	:	val_out <= 4'h0070;
         4'hbca1 	:	val_out <= 4'h0070;
         4'hbca2 	:	val_out <= 4'h0070;
         4'hbca3 	:	val_out <= 4'h0070;
         4'hbca8 	:	val_out <= 4'h006e;
         4'hbca9 	:	val_out <= 4'h006e;
         4'hbcaa 	:	val_out <= 4'h006e;
         4'hbcab 	:	val_out <= 4'h006e;
         4'hbcb0 	:	val_out <= 4'h006c;
         4'hbcb1 	:	val_out <= 4'h006c;
         4'hbcb2 	:	val_out <= 4'h006c;
         4'hbcb3 	:	val_out <= 4'h006c;
         4'hbcb8 	:	val_out <= 4'h006a;
         4'hbcb9 	:	val_out <= 4'h006a;
         4'hbcba 	:	val_out <= 4'h006a;
         4'hbcbb 	:	val_out <= 4'h006a;
         4'hbcc0 	:	val_out <= 4'h0068;
         4'hbcc1 	:	val_out <= 4'h0068;
         4'hbcc2 	:	val_out <= 4'h0068;
         4'hbcc3 	:	val_out <= 4'h0068;
         4'hbcc8 	:	val_out <= 4'h0066;
         4'hbcc9 	:	val_out <= 4'h0066;
         4'hbcca 	:	val_out <= 4'h0066;
         4'hbccb 	:	val_out <= 4'h0066;
         4'hbcd0 	:	val_out <= 4'h0064;
         4'hbcd1 	:	val_out <= 4'h0064;
         4'hbcd2 	:	val_out <= 4'h0064;
         4'hbcd3 	:	val_out <= 4'h0064;
         4'hbcd8 	:	val_out <= 4'h0062;
         4'hbcd9 	:	val_out <= 4'h0062;
         4'hbcda 	:	val_out <= 4'h0062;
         4'hbcdb 	:	val_out <= 4'h0062;
         4'hbce0 	:	val_out <= 4'h0060;
         4'hbce1 	:	val_out <= 4'h0060;
         4'hbce2 	:	val_out <= 4'h0060;
         4'hbce3 	:	val_out <= 4'h0060;
         4'hbce8 	:	val_out <= 4'h005e;
         4'hbce9 	:	val_out <= 4'h005e;
         4'hbcea 	:	val_out <= 4'h005e;
         4'hbceb 	:	val_out <= 4'h005e;
         4'hbcf0 	:	val_out <= 4'h005c;
         4'hbcf1 	:	val_out <= 4'h005c;
         4'hbcf2 	:	val_out <= 4'h005c;
         4'hbcf3 	:	val_out <= 4'h005c;
         4'hbcf8 	:	val_out <= 4'h005a;
         4'hbcf9 	:	val_out <= 4'h005a;
         4'hbcfa 	:	val_out <= 4'h005a;
         4'hbcfb 	:	val_out <= 4'h005a;
         4'hbd00 	:	val_out <= 4'h0058;
         4'hbd01 	:	val_out <= 4'h0058;
         4'hbd02 	:	val_out <= 4'h0058;
         4'hbd03 	:	val_out <= 4'h0058;
         4'hbd08 	:	val_out <= 4'h0056;
         4'hbd09 	:	val_out <= 4'h0056;
         4'hbd0a 	:	val_out <= 4'h0056;
         4'hbd0b 	:	val_out <= 4'h0056;
         4'hbd10 	:	val_out <= 4'h0055;
         4'hbd11 	:	val_out <= 4'h0055;
         4'hbd12 	:	val_out <= 4'h0055;
         4'hbd13 	:	val_out <= 4'h0055;
         4'hbd18 	:	val_out <= 4'h0053;
         4'hbd19 	:	val_out <= 4'h0053;
         4'hbd1a 	:	val_out <= 4'h0053;
         4'hbd1b 	:	val_out <= 4'h0053;
         4'hbd20 	:	val_out <= 4'h0051;
         4'hbd21 	:	val_out <= 4'h0051;
         4'hbd22 	:	val_out <= 4'h0051;
         4'hbd23 	:	val_out <= 4'h0051;
         4'hbd28 	:	val_out <= 4'h004f;
         4'hbd29 	:	val_out <= 4'h004f;
         4'hbd2a 	:	val_out <= 4'h004f;
         4'hbd2b 	:	val_out <= 4'h004f;
         4'hbd30 	:	val_out <= 4'h004e;
         4'hbd31 	:	val_out <= 4'h004e;
         4'hbd32 	:	val_out <= 4'h004e;
         4'hbd33 	:	val_out <= 4'h004e;
         4'hbd38 	:	val_out <= 4'h004c;
         4'hbd39 	:	val_out <= 4'h004c;
         4'hbd3a 	:	val_out <= 4'h004c;
         4'hbd3b 	:	val_out <= 4'h004c;
         4'hbd40 	:	val_out <= 4'h004a;
         4'hbd41 	:	val_out <= 4'h004a;
         4'hbd42 	:	val_out <= 4'h004a;
         4'hbd43 	:	val_out <= 4'h004a;
         4'hbd48 	:	val_out <= 4'h0048;
         4'hbd49 	:	val_out <= 4'h0048;
         4'hbd4a 	:	val_out <= 4'h0048;
         4'hbd4b 	:	val_out <= 4'h0048;
         4'hbd50 	:	val_out <= 4'h0047;
         4'hbd51 	:	val_out <= 4'h0047;
         4'hbd52 	:	val_out <= 4'h0047;
         4'hbd53 	:	val_out <= 4'h0047;
         4'hbd58 	:	val_out <= 4'h0045;
         4'hbd59 	:	val_out <= 4'h0045;
         4'hbd5a 	:	val_out <= 4'h0045;
         4'hbd5b 	:	val_out <= 4'h0045;
         4'hbd60 	:	val_out <= 4'h0043;
         4'hbd61 	:	val_out <= 4'h0043;
         4'hbd62 	:	val_out <= 4'h0043;
         4'hbd63 	:	val_out <= 4'h0043;
         4'hbd68 	:	val_out <= 4'h0042;
         4'hbd69 	:	val_out <= 4'h0042;
         4'hbd6a 	:	val_out <= 4'h0042;
         4'hbd6b 	:	val_out <= 4'h0042;
         4'hbd70 	:	val_out <= 4'h0040;
         4'hbd71 	:	val_out <= 4'h0040;
         4'hbd72 	:	val_out <= 4'h0040;
         4'hbd73 	:	val_out <= 4'h0040;
         4'hbd78 	:	val_out <= 4'h003f;
         4'hbd79 	:	val_out <= 4'h003f;
         4'hbd7a 	:	val_out <= 4'h003f;
         4'hbd7b 	:	val_out <= 4'h003f;
         4'hbd80 	:	val_out <= 4'h003d;
         4'hbd81 	:	val_out <= 4'h003d;
         4'hbd82 	:	val_out <= 4'h003d;
         4'hbd83 	:	val_out <= 4'h003d;
         4'hbd88 	:	val_out <= 4'h003c;
         4'hbd89 	:	val_out <= 4'h003c;
         4'hbd8a 	:	val_out <= 4'h003c;
         4'hbd8b 	:	val_out <= 4'h003c;
         4'hbd90 	:	val_out <= 4'h003a;
         4'hbd91 	:	val_out <= 4'h003a;
         4'hbd92 	:	val_out <= 4'h003a;
         4'hbd93 	:	val_out <= 4'h003a;
         4'hbd98 	:	val_out <= 4'h0039;
         4'hbd99 	:	val_out <= 4'h0039;
         4'hbd9a 	:	val_out <= 4'h0039;
         4'hbd9b 	:	val_out <= 4'h0039;
         4'hbda0 	:	val_out <= 4'h0037;
         4'hbda1 	:	val_out <= 4'h0037;
         4'hbda2 	:	val_out <= 4'h0037;
         4'hbda3 	:	val_out <= 4'h0037;
         4'hbda8 	:	val_out <= 4'h0036;
         4'hbda9 	:	val_out <= 4'h0036;
         4'hbdaa 	:	val_out <= 4'h0036;
         4'hbdab 	:	val_out <= 4'h0036;
         4'hbdb0 	:	val_out <= 4'h0034;
         4'hbdb1 	:	val_out <= 4'h0034;
         4'hbdb2 	:	val_out <= 4'h0034;
         4'hbdb3 	:	val_out <= 4'h0034;
         4'hbdb8 	:	val_out <= 4'h0033;
         4'hbdb9 	:	val_out <= 4'h0033;
         4'hbdba 	:	val_out <= 4'h0033;
         4'hbdbb 	:	val_out <= 4'h0033;
         4'hbdc0 	:	val_out <= 4'h0031;
         4'hbdc1 	:	val_out <= 4'h0031;
         4'hbdc2 	:	val_out <= 4'h0031;
         4'hbdc3 	:	val_out <= 4'h0031;
         4'hbdc8 	:	val_out <= 4'h0030;
         4'hbdc9 	:	val_out <= 4'h0030;
         4'hbdca 	:	val_out <= 4'h0030;
         4'hbdcb 	:	val_out <= 4'h0030;
         4'hbdd0 	:	val_out <= 4'h002f;
         4'hbdd1 	:	val_out <= 4'h002f;
         4'hbdd2 	:	val_out <= 4'h002f;
         4'hbdd3 	:	val_out <= 4'h002f;
         4'hbdd8 	:	val_out <= 4'h002d;
         4'hbdd9 	:	val_out <= 4'h002d;
         4'hbdda 	:	val_out <= 4'h002d;
         4'hbddb 	:	val_out <= 4'h002d;
         4'hbde0 	:	val_out <= 4'h002c;
         4'hbde1 	:	val_out <= 4'h002c;
         4'hbde2 	:	val_out <= 4'h002c;
         4'hbde3 	:	val_out <= 4'h002c;
         4'hbde8 	:	val_out <= 4'h002b;
         4'hbde9 	:	val_out <= 4'h002b;
         4'hbdea 	:	val_out <= 4'h002b;
         4'hbdeb 	:	val_out <= 4'h002b;
         4'hbdf0 	:	val_out <= 4'h0029;
         4'hbdf1 	:	val_out <= 4'h0029;
         4'hbdf2 	:	val_out <= 4'h0029;
         4'hbdf3 	:	val_out <= 4'h0029;
         4'hbdf8 	:	val_out <= 4'h0028;
         4'hbdf9 	:	val_out <= 4'h0028;
         4'hbdfa 	:	val_out <= 4'h0028;
         4'hbdfb 	:	val_out <= 4'h0028;
         4'hbe00 	:	val_out <= 4'h0027;
         4'hbe01 	:	val_out <= 4'h0027;
         4'hbe02 	:	val_out <= 4'h0027;
         4'hbe03 	:	val_out <= 4'h0027;
         4'hbe08 	:	val_out <= 4'h0026;
         4'hbe09 	:	val_out <= 4'h0026;
         4'hbe0a 	:	val_out <= 4'h0026;
         4'hbe0b 	:	val_out <= 4'h0026;
         4'hbe10 	:	val_out <= 4'h0025;
         4'hbe11 	:	val_out <= 4'h0025;
         4'hbe12 	:	val_out <= 4'h0025;
         4'hbe13 	:	val_out <= 4'h0025;
         4'hbe18 	:	val_out <= 4'h0023;
         4'hbe19 	:	val_out <= 4'h0023;
         4'hbe1a 	:	val_out <= 4'h0023;
         4'hbe1b 	:	val_out <= 4'h0023;
         4'hbe20 	:	val_out <= 4'h0022;
         4'hbe21 	:	val_out <= 4'h0022;
         4'hbe22 	:	val_out <= 4'h0022;
         4'hbe23 	:	val_out <= 4'h0022;
         4'hbe28 	:	val_out <= 4'h0021;
         4'hbe29 	:	val_out <= 4'h0021;
         4'hbe2a 	:	val_out <= 4'h0021;
         4'hbe2b 	:	val_out <= 4'h0021;
         4'hbe30 	:	val_out <= 4'h0020;
         4'hbe31 	:	val_out <= 4'h0020;
         4'hbe32 	:	val_out <= 4'h0020;
         4'hbe33 	:	val_out <= 4'h0020;
         4'hbe38 	:	val_out <= 4'h001f;
         4'hbe39 	:	val_out <= 4'h001f;
         4'hbe3a 	:	val_out <= 4'h001f;
         4'hbe3b 	:	val_out <= 4'h001f;
         4'hbe40 	:	val_out <= 4'h001e;
         4'hbe41 	:	val_out <= 4'h001e;
         4'hbe42 	:	val_out <= 4'h001e;
         4'hbe43 	:	val_out <= 4'h001e;
         4'hbe48 	:	val_out <= 4'h001d;
         4'hbe49 	:	val_out <= 4'h001d;
         4'hbe4a 	:	val_out <= 4'h001d;
         4'hbe4b 	:	val_out <= 4'h001d;
         4'hbe50 	:	val_out <= 4'h001c;
         4'hbe51 	:	val_out <= 4'h001c;
         4'hbe52 	:	val_out <= 4'h001c;
         4'hbe53 	:	val_out <= 4'h001c;
         4'hbe58 	:	val_out <= 4'h001b;
         4'hbe59 	:	val_out <= 4'h001b;
         4'hbe5a 	:	val_out <= 4'h001b;
         4'hbe5b 	:	val_out <= 4'h001b;
         4'hbe60 	:	val_out <= 4'h001a;
         4'hbe61 	:	val_out <= 4'h001a;
         4'hbe62 	:	val_out <= 4'h001a;
         4'hbe63 	:	val_out <= 4'h001a;
         4'hbe68 	:	val_out <= 4'h0019;
         4'hbe69 	:	val_out <= 4'h0019;
         4'hbe6a 	:	val_out <= 4'h0019;
         4'hbe6b 	:	val_out <= 4'h0019;
         4'hbe70 	:	val_out <= 4'h0018;
         4'hbe71 	:	val_out <= 4'h0018;
         4'hbe72 	:	val_out <= 4'h0018;
         4'hbe73 	:	val_out <= 4'h0018;
         4'hbe78 	:	val_out <= 4'h0017;
         4'hbe79 	:	val_out <= 4'h0017;
         4'hbe7a 	:	val_out <= 4'h0017;
         4'hbe7b 	:	val_out <= 4'h0017;
         4'hbe80 	:	val_out <= 4'h0016;
         4'hbe81 	:	val_out <= 4'h0016;
         4'hbe82 	:	val_out <= 4'h0016;
         4'hbe83 	:	val_out <= 4'h0016;
         4'hbe88 	:	val_out <= 4'h0015;
         4'hbe89 	:	val_out <= 4'h0015;
         4'hbe8a 	:	val_out <= 4'h0015;
         4'hbe8b 	:	val_out <= 4'h0015;
         4'hbe90 	:	val_out <= 4'h0014;
         4'hbe91 	:	val_out <= 4'h0014;
         4'hbe92 	:	val_out <= 4'h0014;
         4'hbe93 	:	val_out <= 4'h0014;
         4'hbe98 	:	val_out <= 4'h0013;
         4'hbe99 	:	val_out <= 4'h0013;
         4'hbe9a 	:	val_out <= 4'h0013;
         4'hbe9b 	:	val_out <= 4'h0013;
         4'hbea0 	:	val_out <= 4'h0012;
         4'hbea1 	:	val_out <= 4'h0012;
         4'hbea2 	:	val_out <= 4'h0012;
         4'hbea3 	:	val_out <= 4'h0012;
         4'hbea8 	:	val_out <= 4'h0011;
         4'hbea9 	:	val_out <= 4'h0011;
         4'hbeaa 	:	val_out <= 4'h0011;
         4'hbeab 	:	val_out <= 4'h0011;
         4'hbeb0 	:	val_out <= 4'h0011;
         4'hbeb1 	:	val_out <= 4'h0011;
         4'hbeb2 	:	val_out <= 4'h0011;
         4'hbeb3 	:	val_out <= 4'h0011;
         4'hbeb8 	:	val_out <= 4'h0010;
         4'hbeb9 	:	val_out <= 4'h0010;
         4'hbeba 	:	val_out <= 4'h0010;
         4'hbebb 	:	val_out <= 4'h0010;
         4'hbec0 	:	val_out <= 4'h000f;
         4'hbec1 	:	val_out <= 4'h000f;
         4'hbec2 	:	val_out <= 4'h000f;
         4'hbec3 	:	val_out <= 4'h000f;
         4'hbec8 	:	val_out <= 4'h000e;
         4'hbec9 	:	val_out <= 4'h000e;
         4'hbeca 	:	val_out <= 4'h000e;
         4'hbecb 	:	val_out <= 4'h000e;
         4'hbed0 	:	val_out <= 4'h000d;
         4'hbed1 	:	val_out <= 4'h000d;
         4'hbed2 	:	val_out <= 4'h000d;
         4'hbed3 	:	val_out <= 4'h000d;
         4'hbed8 	:	val_out <= 4'h000d;
         4'hbed9 	:	val_out <= 4'h000d;
         4'hbeda 	:	val_out <= 4'h000d;
         4'hbedb 	:	val_out <= 4'h000d;
         4'hbee0 	:	val_out <= 4'h000c;
         4'hbee1 	:	val_out <= 4'h000c;
         4'hbee2 	:	val_out <= 4'h000c;
         4'hbee3 	:	val_out <= 4'h000c;
         4'hbee8 	:	val_out <= 4'h000b;
         4'hbee9 	:	val_out <= 4'h000b;
         4'hbeea 	:	val_out <= 4'h000b;
         4'hbeeb 	:	val_out <= 4'h000b;
         4'hbef0 	:	val_out <= 4'h000b;
         4'hbef1 	:	val_out <= 4'h000b;
         4'hbef2 	:	val_out <= 4'h000b;
         4'hbef3 	:	val_out <= 4'h000b;
         4'hbef8 	:	val_out <= 4'h000a;
         4'hbef9 	:	val_out <= 4'h000a;
         4'hbefa 	:	val_out <= 4'h000a;
         4'hbefb 	:	val_out <= 4'h000a;
         4'hbf00 	:	val_out <= 4'h0009;
         4'hbf01 	:	val_out <= 4'h0009;
         4'hbf02 	:	val_out <= 4'h0009;
         4'hbf03 	:	val_out <= 4'h0009;
         4'hbf08 	:	val_out <= 4'h0009;
         4'hbf09 	:	val_out <= 4'h0009;
         4'hbf0a 	:	val_out <= 4'h0009;
         4'hbf0b 	:	val_out <= 4'h0009;
         4'hbf10 	:	val_out <= 4'h0008;
         4'hbf11 	:	val_out <= 4'h0008;
         4'hbf12 	:	val_out <= 4'h0008;
         4'hbf13 	:	val_out <= 4'h0008;
         4'hbf18 	:	val_out <= 4'h0008;
         4'hbf19 	:	val_out <= 4'h0008;
         4'hbf1a 	:	val_out <= 4'h0008;
         4'hbf1b 	:	val_out <= 4'h0008;
         4'hbf20 	:	val_out <= 4'h0007;
         4'hbf21 	:	val_out <= 4'h0007;
         4'hbf22 	:	val_out <= 4'h0007;
         4'hbf23 	:	val_out <= 4'h0007;
         4'hbf28 	:	val_out <= 4'h0007;
         4'hbf29 	:	val_out <= 4'h0007;
         4'hbf2a 	:	val_out <= 4'h0007;
         4'hbf2b 	:	val_out <= 4'h0007;
         4'hbf30 	:	val_out <= 4'h0006;
         4'hbf31 	:	val_out <= 4'h0006;
         4'hbf32 	:	val_out <= 4'h0006;
         4'hbf33 	:	val_out <= 4'h0006;
         4'hbf38 	:	val_out <= 4'h0006;
         4'hbf39 	:	val_out <= 4'h0006;
         4'hbf3a 	:	val_out <= 4'h0006;
         4'hbf3b 	:	val_out <= 4'h0006;
         4'hbf40 	:	val_out <= 4'h0005;
         4'hbf41 	:	val_out <= 4'h0005;
         4'hbf42 	:	val_out <= 4'h0005;
         4'hbf43 	:	val_out <= 4'h0005;
         4'hbf48 	:	val_out <= 4'h0005;
         4'hbf49 	:	val_out <= 4'h0005;
         4'hbf4a 	:	val_out <= 4'h0005;
         4'hbf4b 	:	val_out <= 4'h0005;
         4'hbf50 	:	val_out <= 4'h0004;
         4'hbf51 	:	val_out <= 4'h0004;
         4'hbf52 	:	val_out <= 4'h0004;
         4'hbf53 	:	val_out <= 4'h0004;
         4'hbf58 	:	val_out <= 4'h0004;
         4'hbf59 	:	val_out <= 4'h0004;
         4'hbf5a 	:	val_out <= 4'h0004;
         4'hbf5b 	:	val_out <= 4'h0004;
         4'hbf60 	:	val_out <= 4'h0003;
         4'hbf61 	:	val_out <= 4'h0003;
         4'hbf62 	:	val_out <= 4'h0003;
         4'hbf63 	:	val_out <= 4'h0003;
         4'hbf68 	:	val_out <= 4'h0003;
         4'hbf69 	:	val_out <= 4'h0003;
         4'hbf6a 	:	val_out <= 4'h0003;
         4'hbf6b 	:	val_out <= 4'h0003;
         4'hbf70 	:	val_out <= 4'h0003;
         4'hbf71 	:	val_out <= 4'h0003;
         4'hbf72 	:	val_out <= 4'h0003;
         4'hbf73 	:	val_out <= 4'h0003;
         4'hbf78 	:	val_out <= 4'h0002;
         4'hbf79 	:	val_out <= 4'h0002;
         4'hbf7a 	:	val_out <= 4'h0002;
         4'hbf7b 	:	val_out <= 4'h0002;
         4'hbf80 	:	val_out <= 4'h0002;
         4'hbf81 	:	val_out <= 4'h0002;
         4'hbf82 	:	val_out <= 4'h0002;
         4'hbf83 	:	val_out <= 4'h0002;
         4'hbf88 	:	val_out <= 4'h0002;
         4'hbf89 	:	val_out <= 4'h0002;
         4'hbf8a 	:	val_out <= 4'h0002;
         4'hbf8b 	:	val_out <= 4'h0002;
         4'hbf90 	:	val_out <= 4'h0001;
         4'hbf91 	:	val_out <= 4'h0001;
         4'hbf92 	:	val_out <= 4'h0001;
         4'hbf93 	:	val_out <= 4'h0001;
         4'hbf98 	:	val_out <= 4'h0001;
         4'hbf99 	:	val_out <= 4'h0001;
         4'hbf9a 	:	val_out <= 4'h0001;
         4'hbf9b 	:	val_out <= 4'h0001;
         4'hbfa0 	:	val_out <= 4'h0001;
         4'hbfa1 	:	val_out <= 4'h0001;
         4'hbfa2 	:	val_out <= 4'h0001;
         4'hbfa3 	:	val_out <= 4'h0001;
         4'hbfa8 	:	val_out <= 4'h0001;
         4'hbfa9 	:	val_out <= 4'h0001;
         4'hbfaa 	:	val_out <= 4'h0001;
         4'hbfab 	:	val_out <= 4'h0001;
         4'hbfb0 	:	val_out <= 4'h0000;
         4'hbfb1 	:	val_out <= 4'h0000;
         4'hbfb2 	:	val_out <= 4'h0000;
         4'hbfb3 	:	val_out <= 4'h0000;
         4'hbfb8 	:	val_out <= 4'h0000;
         4'hbfb9 	:	val_out <= 4'h0000;
         4'hbfba 	:	val_out <= 4'h0000;
         4'hbfbb 	:	val_out <= 4'h0000;
         4'hbfc0 	:	val_out <= 4'h0000;
         4'hbfc1 	:	val_out <= 4'h0000;
         4'hbfc2 	:	val_out <= 4'h0000;
         4'hbfc3 	:	val_out <= 4'h0000;
         4'hbfc8 	:	val_out <= 4'h0000;
         4'hbfc9 	:	val_out <= 4'h0000;
         4'hbfca 	:	val_out <= 4'h0000;
         4'hbfcb 	:	val_out <= 4'h0000;
         4'hbfd0 	:	val_out <= 4'h0000;
         4'hbfd1 	:	val_out <= 4'h0000;
         4'hbfd2 	:	val_out <= 4'h0000;
         4'hbfd3 	:	val_out <= 4'h0000;
         4'hbfd8 	:	val_out <= 4'h0000;
         4'hbfd9 	:	val_out <= 4'h0000;
         4'hbfda 	:	val_out <= 4'h0000;
         4'hbfdb 	:	val_out <= 4'h0000;
         4'hbfe0 	:	val_out <= 4'h0000;
         4'hbfe1 	:	val_out <= 4'h0000;
         4'hbfe2 	:	val_out <= 4'h0000;
         4'hbfe3 	:	val_out <= 4'h0000;
         4'hbfe8 	:	val_out <= 4'h0000;
         4'hbfe9 	:	val_out <= 4'h0000;
         4'hbfea 	:	val_out <= 4'h0000;
         4'hbfeb 	:	val_out <= 4'h0000;
         4'hbff0 	:	val_out <= 4'h0000;
         4'hbff1 	:	val_out <= 4'h0000;
         4'hbff2 	:	val_out <= 4'h0000;
         4'hbff3 	:	val_out <= 4'h0000;
         4'hbff8 	:	val_out <= 4'h0000;
         4'hbff9 	:	val_out <= 4'h0000;
         4'hbffa 	:	val_out <= 4'h0000;
         4'hbffb 	:	val_out <= 4'h0000;
         4'hc000 	:	val_out <= 4'h0000;
         4'hc001 	:	val_out <= 4'h0000;
         4'hc002 	:	val_out <= 4'h0000;
         4'hc003 	:	val_out <= 4'h0000;
         4'hc008 	:	val_out <= 4'h0000;
         4'hc009 	:	val_out <= 4'h0000;
         4'hc00a 	:	val_out <= 4'h0000;
         4'hc00b 	:	val_out <= 4'h0000;
         4'hc010 	:	val_out <= 4'h0000;
         4'hc011 	:	val_out <= 4'h0000;
         4'hc012 	:	val_out <= 4'h0000;
         4'hc013 	:	val_out <= 4'h0000;
         4'hc018 	:	val_out <= 4'h0000;
         4'hc019 	:	val_out <= 4'h0000;
         4'hc01a 	:	val_out <= 4'h0000;
         4'hc01b 	:	val_out <= 4'h0000;
         4'hc020 	:	val_out <= 4'h0000;
         4'hc021 	:	val_out <= 4'h0000;
         4'hc022 	:	val_out <= 4'h0000;
         4'hc023 	:	val_out <= 4'h0000;
         4'hc028 	:	val_out <= 4'h0000;
         4'hc029 	:	val_out <= 4'h0000;
         4'hc02a 	:	val_out <= 4'h0000;
         4'hc02b 	:	val_out <= 4'h0000;
         4'hc030 	:	val_out <= 4'h0000;
         4'hc031 	:	val_out <= 4'h0000;
         4'hc032 	:	val_out <= 4'h0000;
         4'hc033 	:	val_out <= 4'h0000;
         4'hc038 	:	val_out <= 4'h0000;
         4'hc039 	:	val_out <= 4'h0000;
         4'hc03a 	:	val_out <= 4'h0000;
         4'hc03b 	:	val_out <= 4'h0000;
         4'hc040 	:	val_out <= 4'h0000;
         4'hc041 	:	val_out <= 4'h0000;
         4'hc042 	:	val_out <= 4'h0000;
         4'hc043 	:	val_out <= 4'h0000;
         4'hc048 	:	val_out <= 4'h0000;
         4'hc049 	:	val_out <= 4'h0000;
         4'hc04a 	:	val_out <= 4'h0000;
         4'hc04b 	:	val_out <= 4'h0000;
         4'hc050 	:	val_out <= 4'h0000;
         4'hc051 	:	val_out <= 4'h0000;
         4'hc052 	:	val_out <= 4'h0000;
         4'hc053 	:	val_out <= 4'h0000;
         4'hc058 	:	val_out <= 4'h0001;
         4'hc059 	:	val_out <= 4'h0001;
         4'hc05a 	:	val_out <= 4'h0001;
         4'hc05b 	:	val_out <= 4'h0001;
         4'hc060 	:	val_out <= 4'h0001;
         4'hc061 	:	val_out <= 4'h0001;
         4'hc062 	:	val_out <= 4'h0001;
         4'hc063 	:	val_out <= 4'h0001;
         4'hc068 	:	val_out <= 4'h0001;
         4'hc069 	:	val_out <= 4'h0001;
         4'hc06a 	:	val_out <= 4'h0001;
         4'hc06b 	:	val_out <= 4'h0001;
         4'hc070 	:	val_out <= 4'h0001;
         4'hc071 	:	val_out <= 4'h0001;
         4'hc072 	:	val_out <= 4'h0001;
         4'hc073 	:	val_out <= 4'h0001;
         4'hc078 	:	val_out <= 4'h0002;
         4'hc079 	:	val_out <= 4'h0002;
         4'hc07a 	:	val_out <= 4'h0002;
         4'hc07b 	:	val_out <= 4'h0002;
         4'hc080 	:	val_out <= 4'h0002;
         4'hc081 	:	val_out <= 4'h0002;
         4'hc082 	:	val_out <= 4'h0002;
         4'hc083 	:	val_out <= 4'h0002;
         4'hc088 	:	val_out <= 4'h0002;
         4'hc089 	:	val_out <= 4'h0002;
         4'hc08a 	:	val_out <= 4'h0002;
         4'hc08b 	:	val_out <= 4'h0002;
         4'hc090 	:	val_out <= 4'h0003;
         4'hc091 	:	val_out <= 4'h0003;
         4'hc092 	:	val_out <= 4'h0003;
         4'hc093 	:	val_out <= 4'h0003;
         4'hc098 	:	val_out <= 4'h0003;
         4'hc099 	:	val_out <= 4'h0003;
         4'hc09a 	:	val_out <= 4'h0003;
         4'hc09b 	:	val_out <= 4'h0003;
         4'hc0a0 	:	val_out <= 4'h0003;
         4'hc0a1 	:	val_out <= 4'h0003;
         4'hc0a2 	:	val_out <= 4'h0003;
         4'hc0a3 	:	val_out <= 4'h0003;
         4'hc0a8 	:	val_out <= 4'h0004;
         4'hc0a9 	:	val_out <= 4'h0004;
         4'hc0aa 	:	val_out <= 4'h0004;
         4'hc0ab 	:	val_out <= 4'h0004;
         4'hc0b0 	:	val_out <= 4'h0004;
         4'hc0b1 	:	val_out <= 4'h0004;
         4'hc0b2 	:	val_out <= 4'h0004;
         4'hc0b3 	:	val_out <= 4'h0004;
         4'hc0b8 	:	val_out <= 4'h0005;
         4'hc0b9 	:	val_out <= 4'h0005;
         4'hc0ba 	:	val_out <= 4'h0005;
         4'hc0bb 	:	val_out <= 4'h0005;
         4'hc0c0 	:	val_out <= 4'h0005;
         4'hc0c1 	:	val_out <= 4'h0005;
         4'hc0c2 	:	val_out <= 4'h0005;
         4'hc0c3 	:	val_out <= 4'h0005;
         4'hc0c8 	:	val_out <= 4'h0006;
         4'hc0c9 	:	val_out <= 4'h0006;
         4'hc0ca 	:	val_out <= 4'h0006;
         4'hc0cb 	:	val_out <= 4'h0006;
         4'hc0d0 	:	val_out <= 4'h0006;
         4'hc0d1 	:	val_out <= 4'h0006;
         4'hc0d2 	:	val_out <= 4'h0006;
         4'hc0d3 	:	val_out <= 4'h0006;
         4'hc0d8 	:	val_out <= 4'h0007;
         4'hc0d9 	:	val_out <= 4'h0007;
         4'hc0da 	:	val_out <= 4'h0007;
         4'hc0db 	:	val_out <= 4'h0007;
         4'hc0e0 	:	val_out <= 4'h0007;
         4'hc0e1 	:	val_out <= 4'h0007;
         4'hc0e2 	:	val_out <= 4'h0007;
         4'hc0e3 	:	val_out <= 4'h0007;
         4'hc0e8 	:	val_out <= 4'h0008;
         4'hc0e9 	:	val_out <= 4'h0008;
         4'hc0ea 	:	val_out <= 4'h0008;
         4'hc0eb 	:	val_out <= 4'h0008;
         4'hc0f0 	:	val_out <= 4'h0008;
         4'hc0f1 	:	val_out <= 4'h0008;
         4'hc0f2 	:	val_out <= 4'h0008;
         4'hc0f3 	:	val_out <= 4'h0008;
         4'hc0f8 	:	val_out <= 4'h0009;
         4'hc0f9 	:	val_out <= 4'h0009;
         4'hc0fa 	:	val_out <= 4'h0009;
         4'hc0fb 	:	val_out <= 4'h0009;
         4'hc100 	:	val_out <= 4'h0009;
         4'hc101 	:	val_out <= 4'h0009;
         4'hc102 	:	val_out <= 4'h0009;
         4'hc103 	:	val_out <= 4'h0009;
         4'hc108 	:	val_out <= 4'h000a;
         4'hc109 	:	val_out <= 4'h000a;
         4'hc10a 	:	val_out <= 4'h000a;
         4'hc10b 	:	val_out <= 4'h000a;
         4'hc110 	:	val_out <= 4'h000b;
         4'hc111 	:	val_out <= 4'h000b;
         4'hc112 	:	val_out <= 4'h000b;
         4'hc113 	:	val_out <= 4'h000b;
         4'hc118 	:	val_out <= 4'h000b;
         4'hc119 	:	val_out <= 4'h000b;
         4'hc11a 	:	val_out <= 4'h000b;
         4'hc11b 	:	val_out <= 4'h000b;
         4'hc120 	:	val_out <= 4'h000c;
         4'hc121 	:	val_out <= 4'h000c;
         4'hc122 	:	val_out <= 4'h000c;
         4'hc123 	:	val_out <= 4'h000c;
         4'hc128 	:	val_out <= 4'h000d;
         4'hc129 	:	val_out <= 4'h000d;
         4'hc12a 	:	val_out <= 4'h000d;
         4'hc12b 	:	val_out <= 4'h000d;
         4'hc130 	:	val_out <= 4'h000d;
         4'hc131 	:	val_out <= 4'h000d;
         4'hc132 	:	val_out <= 4'h000d;
         4'hc133 	:	val_out <= 4'h000d;
         4'hc138 	:	val_out <= 4'h000e;
         4'hc139 	:	val_out <= 4'h000e;
         4'hc13a 	:	val_out <= 4'h000e;
         4'hc13b 	:	val_out <= 4'h000e;
         4'hc140 	:	val_out <= 4'h000f;
         4'hc141 	:	val_out <= 4'h000f;
         4'hc142 	:	val_out <= 4'h000f;
         4'hc143 	:	val_out <= 4'h000f;
         4'hc148 	:	val_out <= 4'h0010;
         4'hc149 	:	val_out <= 4'h0010;
         4'hc14a 	:	val_out <= 4'h0010;
         4'hc14b 	:	val_out <= 4'h0010;
         4'hc150 	:	val_out <= 4'h0011;
         4'hc151 	:	val_out <= 4'h0011;
         4'hc152 	:	val_out <= 4'h0011;
         4'hc153 	:	val_out <= 4'h0011;
         4'hc158 	:	val_out <= 4'h0011;
         4'hc159 	:	val_out <= 4'h0011;
         4'hc15a 	:	val_out <= 4'h0011;
         4'hc15b 	:	val_out <= 4'h0011;
         4'hc160 	:	val_out <= 4'h0012;
         4'hc161 	:	val_out <= 4'h0012;
         4'hc162 	:	val_out <= 4'h0012;
         4'hc163 	:	val_out <= 4'h0012;
         4'hc168 	:	val_out <= 4'h0013;
         4'hc169 	:	val_out <= 4'h0013;
         4'hc16a 	:	val_out <= 4'h0013;
         4'hc16b 	:	val_out <= 4'h0013;
         4'hc170 	:	val_out <= 4'h0014;
         4'hc171 	:	val_out <= 4'h0014;
         4'hc172 	:	val_out <= 4'h0014;
         4'hc173 	:	val_out <= 4'h0014;
         4'hc178 	:	val_out <= 4'h0015;
         4'hc179 	:	val_out <= 4'h0015;
         4'hc17a 	:	val_out <= 4'h0015;
         4'hc17b 	:	val_out <= 4'h0015;
         4'hc180 	:	val_out <= 4'h0016;
         4'hc181 	:	val_out <= 4'h0016;
         4'hc182 	:	val_out <= 4'h0016;
         4'hc183 	:	val_out <= 4'h0016;
         4'hc188 	:	val_out <= 4'h0017;
         4'hc189 	:	val_out <= 4'h0017;
         4'hc18a 	:	val_out <= 4'h0017;
         4'hc18b 	:	val_out <= 4'h0017;
         4'hc190 	:	val_out <= 4'h0018;
         4'hc191 	:	val_out <= 4'h0018;
         4'hc192 	:	val_out <= 4'h0018;
         4'hc193 	:	val_out <= 4'h0018;
         4'hc198 	:	val_out <= 4'h0019;
         4'hc199 	:	val_out <= 4'h0019;
         4'hc19a 	:	val_out <= 4'h0019;
         4'hc19b 	:	val_out <= 4'h0019;
         4'hc1a0 	:	val_out <= 4'h001a;
         4'hc1a1 	:	val_out <= 4'h001a;
         4'hc1a2 	:	val_out <= 4'h001a;
         4'hc1a3 	:	val_out <= 4'h001a;
         4'hc1a8 	:	val_out <= 4'h001b;
         4'hc1a9 	:	val_out <= 4'h001b;
         4'hc1aa 	:	val_out <= 4'h001b;
         4'hc1ab 	:	val_out <= 4'h001b;
         4'hc1b0 	:	val_out <= 4'h001c;
         4'hc1b1 	:	val_out <= 4'h001c;
         4'hc1b2 	:	val_out <= 4'h001c;
         4'hc1b3 	:	val_out <= 4'h001c;
         4'hc1b8 	:	val_out <= 4'h001d;
         4'hc1b9 	:	val_out <= 4'h001d;
         4'hc1ba 	:	val_out <= 4'h001d;
         4'hc1bb 	:	val_out <= 4'h001d;
         4'hc1c0 	:	val_out <= 4'h001e;
         4'hc1c1 	:	val_out <= 4'h001e;
         4'hc1c2 	:	val_out <= 4'h001e;
         4'hc1c3 	:	val_out <= 4'h001e;
         4'hc1c8 	:	val_out <= 4'h001f;
         4'hc1c9 	:	val_out <= 4'h001f;
         4'hc1ca 	:	val_out <= 4'h001f;
         4'hc1cb 	:	val_out <= 4'h001f;
         4'hc1d0 	:	val_out <= 4'h0020;
         4'hc1d1 	:	val_out <= 4'h0020;
         4'hc1d2 	:	val_out <= 4'h0020;
         4'hc1d3 	:	val_out <= 4'h0020;
         4'hc1d8 	:	val_out <= 4'h0021;
         4'hc1d9 	:	val_out <= 4'h0021;
         4'hc1da 	:	val_out <= 4'h0021;
         4'hc1db 	:	val_out <= 4'h0021;
         4'hc1e0 	:	val_out <= 4'h0022;
         4'hc1e1 	:	val_out <= 4'h0022;
         4'hc1e2 	:	val_out <= 4'h0022;
         4'hc1e3 	:	val_out <= 4'h0022;
         4'hc1e8 	:	val_out <= 4'h0023;
         4'hc1e9 	:	val_out <= 4'h0023;
         4'hc1ea 	:	val_out <= 4'h0023;
         4'hc1eb 	:	val_out <= 4'h0023;
         4'hc1f0 	:	val_out <= 4'h0025;
         4'hc1f1 	:	val_out <= 4'h0025;
         4'hc1f2 	:	val_out <= 4'h0025;
         4'hc1f3 	:	val_out <= 4'h0025;
         4'hc1f8 	:	val_out <= 4'h0026;
         4'hc1f9 	:	val_out <= 4'h0026;
         4'hc1fa 	:	val_out <= 4'h0026;
         4'hc1fb 	:	val_out <= 4'h0026;
         4'hc200 	:	val_out <= 4'h0027;
         4'hc201 	:	val_out <= 4'h0027;
         4'hc202 	:	val_out <= 4'h0027;
         4'hc203 	:	val_out <= 4'h0027;
         4'hc208 	:	val_out <= 4'h0028;
         4'hc209 	:	val_out <= 4'h0028;
         4'hc20a 	:	val_out <= 4'h0028;
         4'hc20b 	:	val_out <= 4'h0028;
         4'hc210 	:	val_out <= 4'h0029;
         4'hc211 	:	val_out <= 4'h0029;
         4'hc212 	:	val_out <= 4'h0029;
         4'hc213 	:	val_out <= 4'h0029;
         4'hc218 	:	val_out <= 4'h002b;
         4'hc219 	:	val_out <= 4'h002b;
         4'hc21a 	:	val_out <= 4'h002b;
         4'hc21b 	:	val_out <= 4'h002b;
         4'hc220 	:	val_out <= 4'h002c;
         4'hc221 	:	val_out <= 4'h002c;
         4'hc222 	:	val_out <= 4'h002c;
         4'hc223 	:	val_out <= 4'h002c;
         4'hc228 	:	val_out <= 4'h002d;
         4'hc229 	:	val_out <= 4'h002d;
         4'hc22a 	:	val_out <= 4'h002d;
         4'hc22b 	:	val_out <= 4'h002d;
         4'hc230 	:	val_out <= 4'h002f;
         4'hc231 	:	val_out <= 4'h002f;
         4'hc232 	:	val_out <= 4'h002f;
         4'hc233 	:	val_out <= 4'h002f;
         4'hc238 	:	val_out <= 4'h0030;
         4'hc239 	:	val_out <= 4'h0030;
         4'hc23a 	:	val_out <= 4'h0030;
         4'hc23b 	:	val_out <= 4'h0030;
         4'hc240 	:	val_out <= 4'h0031;
         4'hc241 	:	val_out <= 4'h0031;
         4'hc242 	:	val_out <= 4'h0031;
         4'hc243 	:	val_out <= 4'h0031;
         4'hc248 	:	val_out <= 4'h0033;
         4'hc249 	:	val_out <= 4'h0033;
         4'hc24a 	:	val_out <= 4'h0033;
         4'hc24b 	:	val_out <= 4'h0033;
         4'hc250 	:	val_out <= 4'h0034;
         4'hc251 	:	val_out <= 4'h0034;
         4'hc252 	:	val_out <= 4'h0034;
         4'hc253 	:	val_out <= 4'h0034;
         4'hc258 	:	val_out <= 4'h0036;
         4'hc259 	:	val_out <= 4'h0036;
         4'hc25a 	:	val_out <= 4'h0036;
         4'hc25b 	:	val_out <= 4'h0036;
         4'hc260 	:	val_out <= 4'h0037;
         4'hc261 	:	val_out <= 4'h0037;
         4'hc262 	:	val_out <= 4'h0037;
         4'hc263 	:	val_out <= 4'h0037;
         4'hc268 	:	val_out <= 4'h0039;
         4'hc269 	:	val_out <= 4'h0039;
         4'hc26a 	:	val_out <= 4'h0039;
         4'hc26b 	:	val_out <= 4'h0039;
         4'hc270 	:	val_out <= 4'h003a;
         4'hc271 	:	val_out <= 4'h003a;
         4'hc272 	:	val_out <= 4'h003a;
         4'hc273 	:	val_out <= 4'h003a;
         4'hc278 	:	val_out <= 4'h003c;
         4'hc279 	:	val_out <= 4'h003c;
         4'hc27a 	:	val_out <= 4'h003c;
         4'hc27b 	:	val_out <= 4'h003c;
         4'hc280 	:	val_out <= 4'h003d;
         4'hc281 	:	val_out <= 4'h003d;
         4'hc282 	:	val_out <= 4'h003d;
         4'hc283 	:	val_out <= 4'h003d;
         4'hc288 	:	val_out <= 4'h003f;
         4'hc289 	:	val_out <= 4'h003f;
         4'hc28a 	:	val_out <= 4'h003f;
         4'hc28b 	:	val_out <= 4'h003f;
         4'hc290 	:	val_out <= 4'h0040;
         4'hc291 	:	val_out <= 4'h0040;
         4'hc292 	:	val_out <= 4'h0040;
         4'hc293 	:	val_out <= 4'h0040;
         4'hc298 	:	val_out <= 4'h0042;
         4'hc299 	:	val_out <= 4'h0042;
         4'hc29a 	:	val_out <= 4'h0042;
         4'hc29b 	:	val_out <= 4'h0042;
         4'hc2a0 	:	val_out <= 4'h0043;
         4'hc2a1 	:	val_out <= 4'h0043;
         4'hc2a2 	:	val_out <= 4'h0043;
         4'hc2a3 	:	val_out <= 4'h0043;
         4'hc2a8 	:	val_out <= 4'h0045;
         4'hc2a9 	:	val_out <= 4'h0045;
         4'hc2aa 	:	val_out <= 4'h0045;
         4'hc2ab 	:	val_out <= 4'h0045;
         4'hc2b0 	:	val_out <= 4'h0047;
         4'hc2b1 	:	val_out <= 4'h0047;
         4'hc2b2 	:	val_out <= 4'h0047;
         4'hc2b3 	:	val_out <= 4'h0047;
         4'hc2b8 	:	val_out <= 4'h0048;
         4'hc2b9 	:	val_out <= 4'h0048;
         4'hc2ba 	:	val_out <= 4'h0048;
         4'hc2bb 	:	val_out <= 4'h0048;
         4'hc2c0 	:	val_out <= 4'h004a;
         4'hc2c1 	:	val_out <= 4'h004a;
         4'hc2c2 	:	val_out <= 4'h004a;
         4'hc2c3 	:	val_out <= 4'h004a;
         4'hc2c8 	:	val_out <= 4'h004c;
         4'hc2c9 	:	val_out <= 4'h004c;
         4'hc2ca 	:	val_out <= 4'h004c;
         4'hc2cb 	:	val_out <= 4'h004c;
         4'hc2d0 	:	val_out <= 4'h004e;
         4'hc2d1 	:	val_out <= 4'h004e;
         4'hc2d2 	:	val_out <= 4'h004e;
         4'hc2d3 	:	val_out <= 4'h004e;
         4'hc2d8 	:	val_out <= 4'h004f;
         4'hc2d9 	:	val_out <= 4'h004f;
         4'hc2da 	:	val_out <= 4'h004f;
         4'hc2db 	:	val_out <= 4'h004f;
         4'hc2e0 	:	val_out <= 4'h0051;
         4'hc2e1 	:	val_out <= 4'h0051;
         4'hc2e2 	:	val_out <= 4'h0051;
         4'hc2e3 	:	val_out <= 4'h0051;
         4'hc2e8 	:	val_out <= 4'h0053;
         4'hc2e9 	:	val_out <= 4'h0053;
         4'hc2ea 	:	val_out <= 4'h0053;
         4'hc2eb 	:	val_out <= 4'h0053;
         4'hc2f0 	:	val_out <= 4'h0055;
         4'hc2f1 	:	val_out <= 4'h0055;
         4'hc2f2 	:	val_out <= 4'h0055;
         4'hc2f3 	:	val_out <= 4'h0055;
         4'hc2f8 	:	val_out <= 4'h0056;
         4'hc2f9 	:	val_out <= 4'h0056;
         4'hc2fa 	:	val_out <= 4'h0056;
         4'hc2fb 	:	val_out <= 4'h0056;
         4'hc300 	:	val_out <= 4'h0058;
         4'hc301 	:	val_out <= 4'h0058;
         4'hc302 	:	val_out <= 4'h0058;
         4'hc303 	:	val_out <= 4'h0058;
         4'hc308 	:	val_out <= 4'h005a;
         4'hc309 	:	val_out <= 4'h005a;
         4'hc30a 	:	val_out <= 4'h005a;
         4'hc30b 	:	val_out <= 4'h005a;
         4'hc310 	:	val_out <= 4'h005c;
         4'hc311 	:	val_out <= 4'h005c;
         4'hc312 	:	val_out <= 4'h005c;
         4'hc313 	:	val_out <= 4'h005c;
         4'hc318 	:	val_out <= 4'h005e;
         4'hc319 	:	val_out <= 4'h005e;
         4'hc31a 	:	val_out <= 4'h005e;
         4'hc31b 	:	val_out <= 4'h005e;
         4'hc320 	:	val_out <= 4'h0060;
         4'hc321 	:	val_out <= 4'h0060;
         4'hc322 	:	val_out <= 4'h0060;
         4'hc323 	:	val_out <= 4'h0060;
         4'hc328 	:	val_out <= 4'h0062;
         4'hc329 	:	val_out <= 4'h0062;
         4'hc32a 	:	val_out <= 4'h0062;
         4'hc32b 	:	val_out <= 4'h0062;
         4'hc330 	:	val_out <= 4'h0064;
         4'hc331 	:	val_out <= 4'h0064;
         4'hc332 	:	val_out <= 4'h0064;
         4'hc333 	:	val_out <= 4'h0064;
         4'hc338 	:	val_out <= 4'h0066;
         4'hc339 	:	val_out <= 4'h0066;
         4'hc33a 	:	val_out <= 4'h0066;
         4'hc33b 	:	val_out <= 4'h0066;
         4'hc340 	:	val_out <= 4'h0068;
         4'hc341 	:	val_out <= 4'h0068;
         4'hc342 	:	val_out <= 4'h0068;
         4'hc343 	:	val_out <= 4'h0068;
         4'hc348 	:	val_out <= 4'h006a;
         4'hc349 	:	val_out <= 4'h006a;
         4'hc34a 	:	val_out <= 4'h006a;
         4'hc34b 	:	val_out <= 4'h006a;
         4'hc350 	:	val_out <= 4'h006c;
         4'hc351 	:	val_out <= 4'h006c;
         4'hc352 	:	val_out <= 4'h006c;
         4'hc353 	:	val_out <= 4'h006c;
         4'hc358 	:	val_out <= 4'h006e;
         4'hc359 	:	val_out <= 4'h006e;
         4'hc35a 	:	val_out <= 4'h006e;
         4'hc35b 	:	val_out <= 4'h006e;
         4'hc360 	:	val_out <= 4'h0070;
         4'hc361 	:	val_out <= 4'h0070;
         4'hc362 	:	val_out <= 4'h0070;
         4'hc363 	:	val_out <= 4'h0070;
         4'hc368 	:	val_out <= 4'h0072;
         4'hc369 	:	val_out <= 4'h0072;
         4'hc36a 	:	val_out <= 4'h0072;
         4'hc36b 	:	val_out <= 4'h0072;
         4'hc370 	:	val_out <= 4'h0074;
         4'hc371 	:	val_out <= 4'h0074;
         4'hc372 	:	val_out <= 4'h0074;
         4'hc373 	:	val_out <= 4'h0074;
         4'hc378 	:	val_out <= 4'h0076;
         4'hc379 	:	val_out <= 4'h0076;
         4'hc37a 	:	val_out <= 4'h0076;
         4'hc37b 	:	val_out <= 4'h0076;
         4'hc380 	:	val_out <= 4'h0078;
         4'hc381 	:	val_out <= 4'h0078;
         4'hc382 	:	val_out <= 4'h0078;
         4'hc383 	:	val_out <= 4'h0078;
         4'hc388 	:	val_out <= 4'h007a;
         4'hc389 	:	val_out <= 4'h007a;
         4'hc38a 	:	val_out <= 4'h007a;
         4'hc38b 	:	val_out <= 4'h007a;
         4'hc390 	:	val_out <= 4'h007d;
         4'hc391 	:	val_out <= 4'h007d;
         4'hc392 	:	val_out <= 4'h007d;
         4'hc393 	:	val_out <= 4'h007d;
         4'hc398 	:	val_out <= 4'h007f;
         4'hc399 	:	val_out <= 4'h007f;
         4'hc39a 	:	val_out <= 4'h007f;
         4'hc39b 	:	val_out <= 4'h007f;
         4'hc3a0 	:	val_out <= 4'h0081;
         4'hc3a1 	:	val_out <= 4'h0081;
         4'hc3a2 	:	val_out <= 4'h0081;
         4'hc3a3 	:	val_out <= 4'h0081;
         4'hc3a8 	:	val_out <= 4'h0083;
         4'hc3a9 	:	val_out <= 4'h0083;
         4'hc3aa 	:	val_out <= 4'h0083;
         4'hc3ab 	:	val_out <= 4'h0083;
         4'hc3b0 	:	val_out <= 4'h0086;
         4'hc3b1 	:	val_out <= 4'h0086;
         4'hc3b2 	:	val_out <= 4'h0086;
         4'hc3b3 	:	val_out <= 4'h0086;
         4'hc3b8 	:	val_out <= 4'h0088;
         4'hc3b9 	:	val_out <= 4'h0088;
         4'hc3ba 	:	val_out <= 4'h0088;
         4'hc3bb 	:	val_out <= 4'h0088;
         4'hc3c0 	:	val_out <= 4'h008a;
         4'hc3c1 	:	val_out <= 4'h008a;
         4'hc3c2 	:	val_out <= 4'h008a;
         4'hc3c3 	:	val_out <= 4'h008a;
         4'hc3c8 	:	val_out <= 4'h008d;
         4'hc3c9 	:	val_out <= 4'h008d;
         4'hc3ca 	:	val_out <= 4'h008d;
         4'hc3cb 	:	val_out <= 4'h008d;
         4'hc3d0 	:	val_out <= 4'h008f;
         4'hc3d1 	:	val_out <= 4'h008f;
         4'hc3d2 	:	val_out <= 4'h008f;
         4'hc3d3 	:	val_out <= 4'h008f;
         4'hc3d8 	:	val_out <= 4'h0091;
         4'hc3d9 	:	val_out <= 4'h0091;
         4'hc3da 	:	val_out <= 4'h0091;
         4'hc3db 	:	val_out <= 4'h0091;
         4'hc3e0 	:	val_out <= 4'h0094;
         4'hc3e1 	:	val_out <= 4'h0094;
         4'hc3e2 	:	val_out <= 4'h0094;
         4'hc3e3 	:	val_out <= 4'h0094;
         4'hc3e8 	:	val_out <= 4'h0096;
         4'hc3e9 	:	val_out <= 4'h0096;
         4'hc3ea 	:	val_out <= 4'h0096;
         4'hc3eb 	:	val_out <= 4'h0096;
         4'hc3f0 	:	val_out <= 4'h0098;
         4'hc3f1 	:	val_out <= 4'h0098;
         4'hc3f2 	:	val_out <= 4'h0098;
         4'hc3f3 	:	val_out <= 4'h0098;
         4'hc3f8 	:	val_out <= 4'h009b;
         4'hc3f9 	:	val_out <= 4'h009b;
         4'hc3fa 	:	val_out <= 4'h009b;
         4'hc3fb 	:	val_out <= 4'h009b;
         4'hc400 	:	val_out <= 4'h009d;
         4'hc401 	:	val_out <= 4'h009d;
         4'hc402 	:	val_out <= 4'h009d;
         4'hc403 	:	val_out <= 4'h009d;
         4'hc408 	:	val_out <= 4'h00a0;
         4'hc409 	:	val_out <= 4'h00a0;
         4'hc40a 	:	val_out <= 4'h00a0;
         4'hc40b 	:	val_out <= 4'h00a0;
         4'hc410 	:	val_out <= 4'h00a2;
         4'hc411 	:	val_out <= 4'h00a2;
         4'hc412 	:	val_out <= 4'h00a2;
         4'hc413 	:	val_out <= 4'h00a2;
         4'hc418 	:	val_out <= 4'h00a5;
         4'hc419 	:	val_out <= 4'h00a5;
         4'hc41a 	:	val_out <= 4'h00a5;
         4'hc41b 	:	val_out <= 4'h00a5;
         4'hc420 	:	val_out <= 4'h00a7;
         4'hc421 	:	val_out <= 4'h00a7;
         4'hc422 	:	val_out <= 4'h00a7;
         4'hc423 	:	val_out <= 4'h00a7;
         4'hc428 	:	val_out <= 4'h00aa;
         4'hc429 	:	val_out <= 4'h00aa;
         4'hc42a 	:	val_out <= 4'h00aa;
         4'hc42b 	:	val_out <= 4'h00aa;
         4'hc430 	:	val_out <= 4'h00ac;
         4'hc431 	:	val_out <= 4'h00ac;
         4'hc432 	:	val_out <= 4'h00ac;
         4'hc433 	:	val_out <= 4'h00ac;
         4'hc438 	:	val_out <= 4'h00af;
         4'hc439 	:	val_out <= 4'h00af;
         4'hc43a 	:	val_out <= 4'h00af;
         4'hc43b 	:	val_out <= 4'h00af;
         4'hc440 	:	val_out <= 4'h00b2;
         4'hc441 	:	val_out <= 4'h00b2;
         4'hc442 	:	val_out <= 4'h00b2;
         4'hc443 	:	val_out <= 4'h00b2;
         4'hc448 	:	val_out <= 4'h00b4;
         4'hc449 	:	val_out <= 4'h00b4;
         4'hc44a 	:	val_out <= 4'h00b4;
         4'hc44b 	:	val_out <= 4'h00b4;
         4'hc450 	:	val_out <= 4'h00b7;
         4'hc451 	:	val_out <= 4'h00b7;
         4'hc452 	:	val_out <= 4'h00b7;
         4'hc453 	:	val_out <= 4'h00b7;
         4'hc458 	:	val_out <= 4'h00ba;
         4'hc459 	:	val_out <= 4'h00ba;
         4'hc45a 	:	val_out <= 4'h00ba;
         4'hc45b 	:	val_out <= 4'h00ba;
         4'hc460 	:	val_out <= 4'h00bc;
         4'hc461 	:	val_out <= 4'h00bc;
         4'hc462 	:	val_out <= 4'h00bc;
         4'hc463 	:	val_out <= 4'h00bc;
         4'hc468 	:	val_out <= 4'h00bf;
         4'hc469 	:	val_out <= 4'h00bf;
         4'hc46a 	:	val_out <= 4'h00bf;
         4'hc46b 	:	val_out <= 4'h00bf;
         4'hc470 	:	val_out <= 4'h00c2;
         4'hc471 	:	val_out <= 4'h00c2;
         4'hc472 	:	val_out <= 4'h00c2;
         4'hc473 	:	val_out <= 4'h00c2;
         4'hc478 	:	val_out <= 4'h00c4;
         4'hc479 	:	val_out <= 4'h00c4;
         4'hc47a 	:	val_out <= 4'h00c4;
         4'hc47b 	:	val_out <= 4'h00c4;
         4'hc480 	:	val_out <= 4'h00c7;
         4'hc481 	:	val_out <= 4'h00c7;
         4'hc482 	:	val_out <= 4'h00c7;
         4'hc483 	:	val_out <= 4'h00c7;
         4'hc488 	:	val_out <= 4'h00ca;
         4'hc489 	:	val_out <= 4'h00ca;
         4'hc48a 	:	val_out <= 4'h00ca;
         4'hc48b 	:	val_out <= 4'h00ca;
         4'hc490 	:	val_out <= 4'h00cd;
         4'hc491 	:	val_out <= 4'h00cd;
         4'hc492 	:	val_out <= 4'h00cd;
         4'hc493 	:	val_out <= 4'h00cd;
         4'hc498 	:	val_out <= 4'h00d0;
         4'hc499 	:	val_out <= 4'h00d0;
         4'hc49a 	:	val_out <= 4'h00d0;
         4'hc49b 	:	val_out <= 4'h00d0;
         4'hc4a0 	:	val_out <= 4'h00d2;
         4'hc4a1 	:	val_out <= 4'h00d2;
         4'hc4a2 	:	val_out <= 4'h00d2;
         4'hc4a3 	:	val_out <= 4'h00d2;
         4'hc4a8 	:	val_out <= 4'h00d5;
         4'hc4a9 	:	val_out <= 4'h00d5;
         4'hc4aa 	:	val_out <= 4'h00d5;
         4'hc4ab 	:	val_out <= 4'h00d5;
         4'hc4b0 	:	val_out <= 4'h00d8;
         4'hc4b1 	:	val_out <= 4'h00d8;
         4'hc4b2 	:	val_out <= 4'h00d8;
         4'hc4b3 	:	val_out <= 4'h00d8;
         4'hc4b8 	:	val_out <= 4'h00db;
         4'hc4b9 	:	val_out <= 4'h00db;
         4'hc4ba 	:	val_out <= 4'h00db;
         4'hc4bb 	:	val_out <= 4'h00db;
         4'hc4c0 	:	val_out <= 4'h00de;
         4'hc4c1 	:	val_out <= 4'h00de;
         4'hc4c2 	:	val_out <= 4'h00de;
         4'hc4c3 	:	val_out <= 4'h00de;
         4'hc4c8 	:	val_out <= 4'h00e1;
         4'hc4c9 	:	val_out <= 4'h00e1;
         4'hc4ca 	:	val_out <= 4'h00e1;
         4'hc4cb 	:	val_out <= 4'h00e1;
         4'hc4d0 	:	val_out <= 4'h00e4;
         4'hc4d1 	:	val_out <= 4'h00e4;
         4'hc4d2 	:	val_out <= 4'h00e4;
         4'hc4d3 	:	val_out <= 4'h00e4;
         4'hc4d8 	:	val_out <= 4'h00e7;
         4'hc4d9 	:	val_out <= 4'h00e7;
         4'hc4da 	:	val_out <= 4'h00e7;
         4'hc4db 	:	val_out <= 4'h00e7;
         4'hc4e0 	:	val_out <= 4'h00ea;
         4'hc4e1 	:	val_out <= 4'h00ea;
         4'hc4e2 	:	val_out <= 4'h00ea;
         4'hc4e3 	:	val_out <= 4'h00ea;
         4'hc4e8 	:	val_out <= 4'h00ed;
         4'hc4e9 	:	val_out <= 4'h00ed;
         4'hc4ea 	:	val_out <= 4'h00ed;
         4'hc4eb 	:	val_out <= 4'h00ed;
         4'hc4f0 	:	val_out <= 4'h00f0;
         4'hc4f1 	:	val_out <= 4'h00f0;
         4'hc4f2 	:	val_out <= 4'h00f0;
         4'hc4f3 	:	val_out <= 4'h00f0;
         4'hc4f8 	:	val_out <= 4'h00f3;
         4'hc4f9 	:	val_out <= 4'h00f3;
         4'hc4fa 	:	val_out <= 4'h00f3;
         4'hc4fb 	:	val_out <= 4'h00f3;
         4'hc500 	:	val_out <= 4'h00f6;
         4'hc501 	:	val_out <= 4'h00f6;
         4'hc502 	:	val_out <= 4'h00f6;
         4'hc503 	:	val_out <= 4'h00f6;
         4'hc508 	:	val_out <= 4'h00f9;
         4'hc509 	:	val_out <= 4'h00f9;
         4'hc50a 	:	val_out <= 4'h00f9;
         4'hc50b 	:	val_out <= 4'h00f9;
         4'hc510 	:	val_out <= 4'h00fc;
         4'hc511 	:	val_out <= 4'h00fc;
         4'hc512 	:	val_out <= 4'h00fc;
         4'hc513 	:	val_out <= 4'h00fc;
         4'hc518 	:	val_out <= 4'h00ff;
         4'hc519 	:	val_out <= 4'h00ff;
         4'hc51a 	:	val_out <= 4'h00ff;
         4'hc51b 	:	val_out <= 4'h00ff;
         4'hc520 	:	val_out <= 4'h0102;
         4'hc521 	:	val_out <= 4'h0102;
         4'hc522 	:	val_out <= 4'h0102;
         4'hc523 	:	val_out <= 4'h0102;
         4'hc528 	:	val_out <= 4'h0106;
         4'hc529 	:	val_out <= 4'h0106;
         4'hc52a 	:	val_out <= 4'h0106;
         4'hc52b 	:	val_out <= 4'h0106;
         4'hc530 	:	val_out <= 4'h0109;
         4'hc531 	:	val_out <= 4'h0109;
         4'hc532 	:	val_out <= 4'h0109;
         4'hc533 	:	val_out <= 4'h0109;
         4'hc538 	:	val_out <= 4'h010c;
         4'hc539 	:	val_out <= 4'h010c;
         4'hc53a 	:	val_out <= 4'h010c;
         4'hc53b 	:	val_out <= 4'h010c;
         4'hc540 	:	val_out <= 4'h010f;
         4'hc541 	:	val_out <= 4'h010f;
         4'hc542 	:	val_out <= 4'h010f;
         4'hc543 	:	val_out <= 4'h010f;
         4'hc548 	:	val_out <= 4'h0112;
         4'hc549 	:	val_out <= 4'h0112;
         4'hc54a 	:	val_out <= 4'h0112;
         4'hc54b 	:	val_out <= 4'h0112;
         4'hc550 	:	val_out <= 4'h0116;
         4'hc551 	:	val_out <= 4'h0116;
         4'hc552 	:	val_out <= 4'h0116;
         4'hc553 	:	val_out <= 4'h0116;
         4'hc558 	:	val_out <= 4'h0119;
         4'hc559 	:	val_out <= 4'h0119;
         4'hc55a 	:	val_out <= 4'h0119;
         4'hc55b 	:	val_out <= 4'h0119;
         4'hc560 	:	val_out <= 4'h011c;
         4'hc561 	:	val_out <= 4'h011c;
         4'hc562 	:	val_out <= 4'h011c;
         4'hc563 	:	val_out <= 4'h011c;
         4'hc568 	:	val_out <= 4'h0120;
         4'hc569 	:	val_out <= 4'h0120;
         4'hc56a 	:	val_out <= 4'h0120;
         4'hc56b 	:	val_out <= 4'h0120;
         4'hc570 	:	val_out <= 4'h0123;
         4'hc571 	:	val_out <= 4'h0123;
         4'hc572 	:	val_out <= 4'h0123;
         4'hc573 	:	val_out <= 4'h0123;
         4'hc578 	:	val_out <= 4'h0126;
         4'hc579 	:	val_out <= 4'h0126;
         4'hc57a 	:	val_out <= 4'h0126;
         4'hc57b 	:	val_out <= 4'h0126;
         4'hc580 	:	val_out <= 4'h012a;
         4'hc581 	:	val_out <= 4'h012a;
         4'hc582 	:	val_out <= 4'h012a;
         4'hc583 	:	val_out <= 4'h012a;
         4'hc588 	:	val_out <= 4'h012d;
         4'hc589 	:	val_out <= 4'h012d;
         4'hc58a 	:	val_out <= 4'h012d;
         4'hc58b 	:	val_out <= 4'h012d;
         4'hc590 	:	val_out <= 4'h0130;
         4'hc591 	:	val_out <= 4'h0130;
         4'hc592 	:	val_out <= 4'h0130;
         4'hc593 	:	val_out <= 4'h0130;
         4'hc598 	:	val_out <= 4'h0134;
         4'hc599 	:	val_out <= 4'h0134;
         4'hc59a 	:	val_out <= 4'h0134;
         4'hc59b 	:	val_out <= 4'h0134;
         4'hc5a0 	:	val_out <= 4'h0137;
         4'hc5a1 	:	val_out <= 4'h0137;
         4'hc5a2 	:	val_out <= 4'h0137;
         4'hc5a3 	:	val_out <= 4'h0137;
         4'hc5a8 	:	val_out <= 4'h013b;
         4'hc5a9 	:	val_out <= 4'h013b;
         4'hc5aa 	:	val_out <= 4'h013b;
         4'hc5ab 	:	val_out <= 4'h013b;
         4'hc5b0 	:	val_out <= 4'h013e;
         4'hc5b1 	:	val_out <= 4'h013e;
         4'hc5b2 	:	val_out <= 4'h013e;
         4'hc5b3 	:	val_out <= 4'h013e;
         4'hc5b8 	:	val_out <= 4'h0142;
         4'hc5b9 	:	val_out <= 4'h0142;
         4'hc5ba 	:	val_out <= 4'h0142;
         4'hc5bb 	:	val_out <= 4'h0142;
         4'hc5c0 	:	val_out <= 4'h0145;
         4'hc5c1 	:	val_out <= 4'h0145;
         4'hc5c2 	:	val_out <= 4'h0145;
         4'hc5c3 	:	val_out <= 4'h0145;
         4'hc5c8 	:	val_out <= 4'h0149;
         4'hc5c9 	:	val_out <= 4'h0149;
         4'hc5ca 	:	val_out <= 4'h0149;
         4'hc5cb 	:	val_out <= 4'h0149;
         4'hc5d0 	:	val_out <= 4'h014c;
         4'hc5d1 	:	val_out <= 4'h014c;
         4'hc5d2 	:	val_out <= 4'h014c;
         4'hc5d3 	:	val_out <= 4'h014c;
         4'hc5d8 	:	val_out <= 4'h0150;
         4'hc5d9 	:	val_out <= 4'h0150;
         4'hc5da 	:	val_out <= 4'h0150;
         4'hc5db 	:	val_out <= 4'h0150;
         4'hc5e0 	:	val_out <= 4'h0154;
         4'hc5e1 	:	val_out <= 4'h0154;
         4'hc5e2 	:	val_out <= 4'h0154;
         4'hc5e3 	:	val_out <= 4'h0154;
         4'hc5e8 	:	val_out <= 4'h0157;
         4'hc5e9 	:	val_out <= 4'h0157;
         4'hc5ea 	:	val_out <= 4'h0157;
         4'hc5eb 	:	val_out <= 4'h0157;
         4'hc5f0 	:	val_out <= 4'h015b;
         4'hc5f1 	:	val_out <= 4'h015b;
         4'hc5f2 	:	val_out <= 4'h015b;
         4'hc5f3 	:	val_out <= 4'h015b;
         4'hc5f8 	:	val_out <= 4'h015e;
         4'hc5f9 	:	val_out <= 4'h015e;
         4'hc5fa 	:	val_out <= 4'h015e;
         4'hc5fb 	:	val_out <= 4'h015e;
         4'hc600 	:	val_out <= 4'h0162;
         4'hc601 	:	val_out <= 4'h0162;
         4'hc602 	:	val_out <= 4'h0162;
         4'hc603 	:	val_out <= 4'h0162;
         4'hc608 	:	val_out <= 4'h0166;
         4'hc609 	:	val_out <= 4'h0166;
         4'hc60a 	:	val_out <= 4'h0166;
         4'hc60b 	:	val_out <= 4'h0166;
         4'hc610 	:	val_out <= 4'h016a;
         4'hc611 	:	val_out <= 4'h016a;
         4'hc612 	:	val_out <= 4'h016a;
         4'hc613 	:	val_out <= 4'h016a;
         4'hc618 	:	val_out <= 4'h016d;
         4'hc619 	:	val_out <= 4'h016d;
         4'hc61a 	:	val_out <= 4'h016d;
         4'hc61b 	:	val_out <= 4'h016d;
         4'hc620 	:	val_out <= 4'h0171;
         4'hc621 	:	val_out <= 4'h0171;
         4'hc622 	:	val_out <= 4'h0171;
         4'hc623 	:	val_out <= 4'h0171;
         4'hc628 	:	val_out <= 4'h0175;
         4'hc629 	:	val_out <= 4'h0175;
         4'hc62a 	:	val_out <= 4'h0175;
         4'hc62b 	:	val_out <= 4'h0175;
         4'hc630 	:	val_out <= 4'h0179;
         4'hc631 	:	val_out <= 4'h0179;
         4'hc632 	:	val_out <= 4'h0179;
         4'hc633 	:	val_out <= 4'h0179;
         4'hc638 	:	val_out <= 4'h017c;
         4'hc639 	:	val_out <= 4'h017c;
         4'hc63a 	:	val_out <= 4'h017c;
         4'hc63b 	:	val_out <= 4'h017c;
         4'hc640 	:	val_out <= 4'h0180;
         4'hc641 	:	val_out <= 4'h0180;
         4'hc642 	:	val_out <= 4'h0180;
         4'hc643 	:	val_out <= 4'h0180;
         4'hc648 	:	val_out <= 4'h0184;
         4'hc649 	:	val_out <= 4'h0184;
         4'hc64a 	:	val_out <= 4'h0184;
         4'hc64b 	:	val_out <= 4'h0184;
         4'hc650 	:	val_out <= 4'h0188;
         4'hc651 	:	val_out <= 4'h0188;
         4'hc652 	:	val_out <= 4'h0188;
         4'hc653 	:	val_out <= 4'h0188;
         4'hc658 	:	val_out <= 4'h018c;
         4'hc659 	:	val_out <= 4'h018c;
         4'hc65a 	:	val_out <= 4'h018c;
         4'hc65b 	:	val_out <= 4'h018c;
         4'hc660 	:	val_out <= 4'h0190;
         4'hc661 	:	val_out <= 4'h0190;
         4'hc662 	:	val_out <= 4'h0190;
         4'hc663 	:	val_out <= 4'h0190;
         4'hc668 	:	val_out <= 4'h0194;
         4'hc669 	:	val_out <= 4'h0194;
         4'hc66a 	:	val_out <= 4'h0194;
         4'hc66b 	:	val_out <= 4'h0194;
         4'hc670 	:	val_out <= 4'h0198;
         4'hc671 	:	val_out <= 4'h0198;
         4'hc672 	:	val_out <= 4'h0198;
         4'hc673 	:	val_out <= 4'h0198;
         4'hc678 	:	val_out <= 4'h019c;
         4'hc679 	:	val_out <= 4'h019c;
         4'hc67a 	:	val_out <= 4'h019c;
         4'hc67b 	:	val_out <= 4'h019c;
         4'hc680 	:	val_out <= 4'h01a0;
         4'hc681 	:	val_out <= 4'h01a0;
         4'hc682 	:	val_out <= 4'h01a0;
         4'hc683 	:	val_out <= 4'h01a0;
         4'hc688 	:	val_out <= 4'h01a4;
         4'hc689 	:	val_out <= 4'h01a4;
         4'hc68a 	:	val_out <= 4'h01a4;
         4'hc68b 	:	val_out <= 4'h01a4;
         4'hc690 	:	val_out <= 4'h01a8;
         4'hc691 	:	val_out <= 4'h01a8;
         4'hc692 	:	val_out <= 4'h01a8;
         4'hc693 	:	val_out <= 4'h01a8;
         4'hc698 	:	val_out <= 4'h01ac;
         4'hc699 	:	val_out <= 4'h01ac;
         4'hc69a 	:	val_out <= 4'h01ac;
         4'hc69b 	:	val_out <= 4'h01ac;
         4'hc6a0 	:	val_out <= 4'h01b0;
         4'hc6a1 	:	val_out <= 4'h01b0;
         4'hc6a2 	:	val_out <= 4'h01b0;
         4'hc6a3 	:	val_out <= 4'h01b0;
         4'hc6a8 	:	val_out <= 4'h01b4;
         4'hc6a9 	:	val_out <= 4'h01b4;
         4'hc6aa 	:	val_out <= 4'h01b4;
         4'hc6ab 	:	val_out <= 4'h01b4;
         4'hc6b0 	:	val_out <= 4'h01b8;
         4'hc6b1 	:	val_out <= 4'h01b8;
         4'hc6b2 	:	val_out <= 4'h01b8;
         4'hc6b3 	:	val_out <= 4'h01b8;
         4'hc6b8 	:	val_out <= 4'h01bc;
         4'hc6b9 	:	val_out <= 4'h01bc;
         4'hc6ba 	:	val_out <= 4'h01bc;
         4'hc6bb 	:	val_out <= 4'h01bc;
         4'hc6c0 	:	val_out <= 4'h01c0;
         4'hc6c1 	:	val_out <= 4'h01c0;
         4'hc6c2 	:	val_out <= 4'h01c0;
         4'hc6c3 	:	val_out <= 4'h01c0;
         4'hc6c8 	:	val_out <= 4'h01c4;
         4'hc6c9 	:	val_out <= 4'h01c4;
         4'hc6ca 	:	val_out <= 4'h01c4;
         4'hc6cb 	:	val_out <= 4'h01c4;
         4'hc6d0 	:	val_out <= 4'h01c8;
         4'hc6d1 	:	val_out <= 4'h01c8;
         4'hc6d2 	:	val_out <= 4'h01c8;
         4'hc6d3 	:	val_out <= 4'h01c8;
         4'hc6d8 	:	val_out <= 4'h01cd;
         4'hc6d9 	:	val_out <= 4'h01cd;
         4'hc6da 	:	val_out <= 4'h01cd;
         4'hc6db 	:	val_out <= 4'h01cd;
         4'hc6e0 	:	val_out <= 4'h01d1;
         4'hc6e1 	:	val_out <= 4'h01d1;
         4'hc6e2 	:	val_out <= 4'h01d1;
         4'hc6e3 	:	val_out <= 4'h01d1;
         4'hc6e8 	:	val_out <= 4'h01d5;
         4'hc6e9 	:	val_out <= 4'h01d5;
         4'hc6ea 	:	val_out <= 4'h01d5;
         4'hc6eb 	:	val_out <= 4'h01d5;
         4'hc6f0 	:	val_out <= 4'h01d9;
         4'hc6f1 	:	val_out <= 4'h01d9;
         4'hc6f2 	:	val_out <= 4'h01d9;
         4'hc6f3 	:	val_out <= 4'h01d9;
         4'hc6f8 	:	val_out <= 4'h01de;
         4'hc6f9 	:	val_out <= 4'h01de;
         4'hc6fa 	:	val_out <= 4'h01de;
         4'hc6fb 	:	val_out <= 4'h01de;
         4'hc700 	:	val_out <= 4'h01e2;
         4'hc701 	:	val_out <= 4'h01e2;
         4'hc702 	:	val_out <= 4'h01e2;
         4'hc703 	:	val_out <= 4'h01e2;
         4'hc708 	:	val_out <= 4'h01e6;
         4'hc709 	:	val_out <= 4'h01e6;
         4'hc70a 	:	val_out <= 4'h01e6;
         4'hc70b 	:	val_out <= 4'h01e6;
         4'hc710 	:	val_out <= 4'h01eb;
         4'hc711 	:	val_out <= 4'h01eb;
         4'hc712 	:	val_out <= 4'h01eb;
         4'hc713 	:	val_out <= 4'h01eb;
         4'hc718 	:	val_out <= 4'h01ef;
         4'hc719 	:	val_out <= 4'h01ef;
         4'hc71a 	:	val_out <= 4'h01ef;
         4'hc71b 	:	val_out <= 4'h01ef;
         4'hc720 	:	val_out <= 4'h01f3;
         4'hc721 	:	val_out <= 4'h01f3;
         4'hc722 	:	val_out <= 4'h01f3;
         4'hc723 	:	val_out <= 4'h01f3;
         4'hc728 	:	val_out <= 4'h01f8;
         4'hc729 	:	val_out <= 4'h01f8;
         4'hc72a 	:	val_out <= 4'h01f8;
         4'hc72b 	:	val_out <= 4'h01f8;
         4'hc730 	:	val_out <= 4'h01fc;
         4'hc731 	:	val_out <= 4'h01fc;
         4'hc732 	:	val_out <= 4'h01fc;
         4'hc733 	:	val_out <= 4'h01fc;
         4'hc738 	:	val_out <= 4'h0200;
         4'hc739 	:	val_out <= 4'h0200;
         4'hc73a 	:	val_out <= 4'h0200;
         4'hc73b 	:	val_out <= 4'h0200;
         4'hc740 	:	val_out <= 4'h0205;
         4'hc741 	:	val_out <= 4'h0205;
         4'hc742 	:	val_out <= 4'h0205;
         4'hc743 	:	val_out <= 4'h0205;
         4'hc748 	:	val_out <= 4'h0209;
         4'hc749 	:	val_out <= 4'h0209;
         4'hc74a 	:	val_out <= 4'h0209;
         4'hc74b 	:	val_out <= 4'h0209;
         4'hc750 	:	val_out <= 4'h020e;
         4'hc751 	:	val_out <= 4'h020e;
         4'hc752 	:	val_out <= 4'h020e;
         4'hc753 	:	val_out <= 4'h020e;
         4'hc758 	:	val_out <= 4'h0212;
         4'hc759 	:	val_out <= 4'h0212;
         4'hc75a 	:	val_out <= 4'h0212;
         4'hc75b 	:	val_out <= 4'h0212;
         4'hc760 	:	val_out <= 4'h0217;
         4'hc761 	:	val_out <= 4'h0217;
         4'hc762 	:	val_out <= 4'h0217;
         4'hc763 	:	val_out <= 4'h0217;
         4'hc768 	:	val_out <= 4'h021b;
         4'hc769 	:	val_out <= 4'h021b;
         4'hc76a 	:	val_out <= 4'h021b;
         4'hc76b 	:	val_out <= 4'h021b;
         4'hc770 	:	val_out <= 4'h0220;
         4'hc771 	:	val_out <= 4'h0220;
         4'hc772 	:	val_out <= 4'h0220;
         4'hc773 	:	val_out <= 4'h0220;
         4'hc778 	:	val_out <= 4'h0225;
         4'hc779 	:	val_out <= 4'h0225;
         4'hc77a 	:	val_out <= 4'h0225;
         4'hc77b 	:	val_out <= 4'h0225;
         4'hc780 	:	val_out <= 4'h0229;
         4'hc781 	:	val_out <= 4'h0229;
         4'hc782 	:	val_out <= 4'h0229;
         4'hc783 	:	val_out <= 4'h0229;
         4'hc788 	:	val_out <= 4'h022e;
         4'hc789 	:	val_out <= 4'h022e;
         4'hc78a 	:	val_out <= 4'h022e;
         4'hc78b 	:	val_out <= 4'h022e;
         4'hc790 	:	val_out <= 4'h0232;
         4'hc791 	:	val_out <= 4'h0232;
         4'hc792 	:	val_out <= 4'h0232;
         4'hc793 	:	val_out <= 4'h0232;
         4'hc798 	:	val_out <= 4'h0237;
         4'hc799 	:	val_out <= 4'h0237;
         4'hc79a 	:	val_out <= 4'h0237;
         4'hc79b 	:	val_out <= 4'h0237;
         4'hc7a0 	:	val_out <= 4'h023c;
         4'hc7a1 	:	val_out <= 4'h023c;
         4'hc7a2 	:	val_out <= 4'h023c;
         4'hc7a3 	:	val_out <= 4'h023c;
         4'hc7a8 	:	val_out <= 4'h0240;
         4'hc7a9 	:	val_out <= 4'h0240;
         4'hc7aa 	:	val_out <= 4'h0240;
         4'hc7ab 	:	val_out <= 4'h0240;
         4'hc7b0 	:	val_out <= 4'h0245;
         4'hc7b1 	:	val_out <= 4'h0245;
         4'hc7b2 	:	val_out <= 4'h0245;
         4'hc7b3 	:	val_out <= 4'h0245;
         4'hc7b8 	:	val_out <= 4'h024a;
         4'hc7b9 	:	val_out <= 4'h024a;
         4'hc7ba 	:	val_out <= 4'h024a;
         4'hc7bb 	:	val_out <= 4'h024a;
         4'hc7c0 	:	val_out <= 4'h024f;
         4'hc7c1 	:	val_out <= 4'h024f;
         4'hc7c2 	:	val_out <= 4'h024f;
         4'hc7c3 	:	val_out <= 4'h024f;
         4'hc7c8 	:	val_out <= 4'h0253;
         4'hc7c9 	:	val_out <= 4'h0253;
         4'hc7ca 	:	val_out <= 4'h0253;
         4'hc7cb 	:	val_out <= 4'h0253;
         4'hc7d0 	:	val_out <= 4'h0258;
         4'hc7d1 	:	val_out <= 4'h0258;
         4'hc7d2 	:	val_out <= 4'h0258;
         4'hc7d3 	:	val_out <= 4'h0258;
         4'hc7d8 	:	val_out <= 4'h025d;
         4'hc7d9 	:	val_out <= 4'h025d;
         4'hc7da 	:	val_out <= 4'h025d;
         4'hc7db 	:	val_out <= 4'h025d;
         4'hc7e0 	:	val_out <= 4'h0262;
         4'hc7e1 	:	val_out <= 4'h0262;
         4'hc7e2 	:	val_out <= 4'h0262;
         4'hc7e3 	:	val_out <= 4'h0262;
         4'hc7e8 	:	val_out <= 4'h0267;
         4'hc7e9 	:	val_out <= 4'h0267;
         4'hc7ea 	:	val_out <= 4'h0267;
         4'hc7eb 	:	val_out <= 4'h0267;
         4'hc7f0 	:	val_out <= 4'h026b;
         4'hc7f1 	:	val_out <= 4'h026b;
         4'hc7f2 	:	val_out <= 4'h026b;
         4'hc7f3 	:	val_out <= 4'h026b;
         4'hc7f8 	:	val_out <= 4'h0270;
         4'hc7f9 	:	val_out <= 4'h0270;
         4'hc7fa 	:	val_out <= 4'h0270;
         4'hc7fb 	:	val_out <= 4'h0270;
         4'hc800 	:	val_out <= 4'h0275;
         4'hc801 	:	val_out <= 4'h0275;
         4'hc802 	:	val_out <= 4'h0275;
         4'hc803 	:	val_out <= 4'h0275;
         4'hc808 	:	val_out <= 4'h027a;
         4'hc809 	:	val_out <= 4'h027a;
         4'hc80a 	:	val_out <= 4'h027a;
         4'hc80b 	:	val_out <= 4'h027a;
         4'hc810 	:	val_out <= 4'h027f;
         4'hc811 	:	val_out <= 4'h027f;
         4'hc812 	:	val_out <= 4'h027f;
         4'hc813 	:	val_out <= 4'h027f;
         4'hc818 	:	val_out <= 4'h0284;
         4'hc819 	:	val_out <= 4'h0284;
         4'hc81a 	:	val_out <= 4'h0284;
         4'hc81b 	:	val_out <= 4'h0284;
         4'hc820 	:	val_out <= 4'h0289;
         4'hc821 	:	val_out <= 4'h0289;
         4'hc822 	:	val_out <= 4'h0289;
         4'hc823 	:	val_out <= 4'h0289;
         4'hc828 	:	val_out <= 4'h028e;
         4'hc829 	:	val_out <= 4'h028e;
         4'hc82a 	:	val_out <= 4'h028e;
         4'hc82b 	:	val_out <= 4'h028e;
         4'hc830 	:	val_out <= 4'h0293;
         4'hc831 	:	val_out <= 4'h0293;
         4'hc832 	:	val_out <= 4'h0293;
         4'hc833 	:	val_out <= 4'h0293;
         4'hc838 	:	val_out <= 4'h0298;
         4'hc839 	:	val_out <= 4'h0298;
         4'hc83a 	:	val_out <= 4'h0298;
         4'hc83b 	:	val_out <= 4'h0298;
         4'hc840 	:	val_out <= 4'h029d;
         4'hc841 	:	val_out <= 4'h029d;
         4'hc842 	:	val_out <= 4'h029d;
         4'hc843 	:	val_out <= 4'h029d;
         4'hc848 	:	val_out <= 4'h02a2;
         4'hc849 	:	val_out <= 4'h02a2;
         4'hc84a 	:	val_out <= 4'h02a2;
         4'hc84b 	:	val_out <= 4'h02a2;
         4'hc850 	:	val_out <= 4'h02a7;
         4'hc851 	:	val_out <= 4'h02a7;
         4'hc852 	:	val_out <= 4'h02a7;
         4'hc853 	:	val_out <= 4'h02a7;
         4'hc858 	:	val_out <= 4'h02ac;
         4'hc859 	:	val_out <= 4'h02ac;
         4'hc85a 	:	val_out <= 4'h02ac;
         4'hc85b 	:	val_out <= 4'h02ac;
         4'hc860 	:	val_out <= 4'h02b1;
         4'hc861 	:	val_out <= 4'h02b1;
         4'hc862 	:	val_out <= 4'h02b1;
         4'hc863 	:	val_out <= 4'h02b1;
         4'hc868 	:	val_out <= 4'h02b6;
         4'hc869 	:	val_out <= 4'h02b6;
         4'hc86a 	:	val_out <= 4'h02b6;
         4'hc86b 	:	val_out <= 4'h02b6;
         4'hc870 	:	val_out <= 4'h02bc;
         4'hc871 	:	val_out <= 4'h02bc;
         4'hc872 	:	val_out <= 4'h02bc;
         4'hc873 	:	val_out <= 4'h02bc;
         4'hc878 	:	val_out <= 4'h02c1;
         4'hc879 	:	val_out <= 4'h02c1;
         4'hc87a 	:	val_out <= 4'h02c1;
         4'hc87b 	:	val_out <= 4'h02c1;
         4'hc880 	:	val_out <= 4'h02c6;
         4'hc881 	:	val_out <= 4'h02c6;
         4'hc882 	:	val_out <= 4'h02c6;
         4'hc883 	:	val_out <= 4'h02c6;
         4'hc888 	:	val_out <= 4'h02cb;
         4'hc889 	:	val_out <= 4'h02cb;
         4'hc88a 	:	val_out <= 4'h02cb;
         4'hc88b 	:	val_out <= 4'h02cb;
         4'hc890 	:	val_out <= 4'h02d0;
         4'hc891 	:	val_out <= 4'h02d0;
         4'hc892 	:	val_out <= 4'h02d0;
         4'hc893 	:	val_out <= 4'h02d0;
         4'hc898 	:	val_out <= 4'h02d6;
         4'hc899 	:	val_out <= 4'h02d6;
         4'hc89a 	:	val_out <= 4'h02d6;
         4'hc89b 	:	val_out <= 4'h02d6;
         4'hc8a0 	:	val_out <= 4'h02db;
         4'hc8a1 	:	val_out <= 4'h02db;
         4'hc8a2 	:	val_out <= 4'h02db;
         4'hc8a3 	:	val_out <= 4'h02db;
         4'hc8a8 	:	val_out <= 4'h02e0;
         4'hc8a9 	:	val_out <= 4'h02e0;
         4'hc8aa 	:	val_out <= 4'h02e0;
         4'hc8ab 	:	val_out <= 4'h02e0;
         4'hc8b0 	:	val_out <= 4'h02e6;
         4'hc8b1 	:	val_out <= 4'h02e6;
         4'hc8b2 	:	val_out <= 4'h02e6;
         4'hc8b3 	:	val_out <= 4'h02e6;
         4'hc8b8 	:	val_out <= 4'h02eb;
         4'hc8b9 	:	val_out <= 4'h02eb;
         4'hc8ba 	:	val_out <= 4'h02eb;
         4'hc8bb 	:	val_out <= 4'h02eb;
         4'hc8c0 	:	val_out <= 4'h02f0;
         4'hc8c1 	:	val_out <= 4'h02f0;
         4'hc8c2 	:	val_out <= 4'h02f0;
         4'hc8c3 	:	val_out <= 4'h02f0;
         4'hc8c8 	:	val_out <= 4'h02f6;
         4'hc8c9 	:	val_out <= 4'h02f6;
         4'hc8ca 	:	val_out <= 4'h02f6;
         4'hc8cb 	:	val_out <= 4'h02f6;
         4'hc8d0 	:	val_out <= 4'h02fb;
         4'hc8d1 	:	val_out <= 4'h02fb;
         4'hc8d2 	:	val_out <= 4'h02fb;
         4'hc8d3 	:	val_out <= 4'h02fb;
         4'hc8d8 	:	val_out <= 4'h0300;
         4'hc8d9 	:	val_out <= 4'h0300;
         4'hc8da 	:	val_out <= 4'h0300;
         4'hc8db 	:	val_out <= 4'h0300;
         4'hc8e0 	:	val_out <= 4'h0306;
         4'hc8e1 	:	val_out <= 4'h0306;
         4'hc8e2 	:	val_out <= 4'h0306;
         4'hc8e3 	:	val_out <= 4'h0306;
         4'hc8e8 	:	val_out <= 4'h030b;
         4'hc8e9 	:	val_out <= 4'h030b;
         4'hc8ea 	:	val_out <= 4'h030b;
         4'hc8eb 	:	val_out <= 4'h030b;
         4'hc8f0 	:	val_out <= 4'h0311;
         4'hc8f1 	:	val_out <= 4'h0311;
         4'hc8f2 	:	val_out <= 4'h0311;
         4'hc8f3 	:	val_out <= 4'h0311;
         4'hc8f8 	:	val_out <= 4'h0316;
         4'hc8f9 	:	val_out <= 4'h0316;
         4'hc8fa 	:	val_out <= 4'h0316;
         4'hc8fb 	:	val_out <= 4'h0316;
         4'hc900 	:	val_out <= 4'h031c;
         4'hc901 	:	val_out <= 4'h031c;
         4'hc902 	:	val_out <= 4'h031c;
         4'hc903 	:	val_out <= 4'h031c;
         4'hc908 	:	val_out <= 4'h0321;
         4'hc909 	:	val_out <= 4'h0321;
         4'hc90a 	:	val_out <= 4'h0321;
         4'hc90b 	:	val_out <= 4'h0321;
         4'hc910 	:	val_out <= 4'h0327;
         4'hc911 	:	val_out <= 4'h0327;
         4'hc912 	:	val_out <= 4'h0327;
         4'hc913 	:	val_out <= 4'h0327;
         4'hc918 	:	val_out <= 4'h032c;
         4'hc919 	:	val_out <= 4'h032c;
         4'hc91a 	:	val_out <= 4'h032c;
         4'hc91b 	:	val_out <= 4'h032c;
         4'hc920 	:	val_out <= 4'h0332;
         4'hc921 	:	val_out <= 4'h0332;
         4'hc922 	:	val_out <= 4'h0332;
         4'hc923 	:	val_out <= 4'h0332;
         4'hc928 	:	val_out <= 4'h0337;
         4'hc929 	:	val_out <= 4'h0337;
         4'hc92a 	:	val_out <= 4'h0337;
         4'hc92b 	:	val_out <= 4'h0337;
         4'hc930 	:	val_out <= 4'h033d;
         4'hc931 	:	val_out <= 4'h033d;
         4'hc932 	:	val_out <= 4'h033d;
         4'hc933 	:	val_out <= 4'h033d;
         4'hc938 	:	val_out <= 4'h0343;
         4'hc939 	:	val_out <= 4'h0343;
         4'hc93a 	:	val_out <= 4'h0343;
         4'hc93b 	:	val_out <= 4'h0343;
         4'hc940 	:	val_out <= 4'h0348;
         4'hc941 	:	val_out <= 4'h0348;
         4'hc942 	:	val_out <= 4'h0348;
         4'hc943 	:	val_out <= 4'h0348;
         4'hc948 	:	val_out <= 4'h034e;
         4'hc949 	:	val_out <= 4'h034e;
         4'hc94a 	:	val_out <= 4'h034e;
         4'hc94b 	:	val_out <= 4'h034e;
         4'hc950 	:	val_out <= 4'h0354;
         4'hc951 	:	val_out <= 4'h0354;
         4'hc952 	:	val_out <= 4'h0354;
         4'hc953 	:	val_out <= 4'h0354;
         4'hc958 	:	val_out <= 4'h0359;
         4'hc959 	:	val_out <= 4'h0359;
         4'hc95a 	:	val_out <= 4'h0359;
         4'hc95b 	:	val_out <= 4'h0359;
         4'hc960 	:	val_out <= 4'h035f;
         4'hc961 	:	val_out <= 4'h035f;
         4'hc962 	:	val_out <= 4'h035f;
         4'hc963 	:	val_out <= 4'h035f;
         4'hc968 	:	val_out <= 4'h0365;
         4'hc969 	:	val_out <= 4'h0365;
         4'hc96a 	:	val_out <= 4'h0365;
         4'hc96b 	:	val_out <= 4'h0365;
         4'hc970 	:	val_out <= 4'h036b;
         4'hc971 	:	val_out <= 4'h036b;
         4'hc972 	:	val_out <= 4'h036b;
         4'hc973 	:	val_out <= 4'h036b;
         4'hc978 	:	val_out <= 4'h0370;
         4'hc979 	:	val_out <= 4'h0370;
         4'hc97a 	:	val_out <= 4'h0370;
         4'hc97b 	:	val_out <= 4'h0370;
         4'hc980 	:	val_out <= 4'h0376;
         4'hc981 	:	val_out <= 4'h0376;
         4'hc982 	:	val_out <= 4'h0376;
         4'hc983 	:	val_out <= 4'h0376;
         4'hc988 	:	val_out <= 4'h037c;
         4'hc989 	:	val_out <= 4'h037c;
         4'hc98a 	:	val_out <= 4'h037c;
         4'hc98b 	:	val_out <= 4'h037c;
         4'hc990 	:	val_out <= 4'h0382;
         4'hc991 	:	val_out <= 4'h0382;
         4'hc992 	:	val_out <= 4'h0382;
         4'hc993 	:	val_out <= 4'h0382;
         4'hc998 	:	val_out <= 4'h0388;
         4'hc999 	:	val_out <= 4'h0388;
         4'hc99a 	:	val_out <= 4'h0388;
         4'hc99b 	:	val_out <= 4'h0388;
         4'hc9a0 	:	val_out <= 4'h038e;
         4'hc9a1 	:	val_out <= 4'h038e;
         4'hc9a2 	:	val_out <= 4'h038e;
         4'hc9a3 	:	val_out <= 4'h038e;
         4'hc9a8 	:	val_out <= 4'h0393;
         4'hc9a9 	:	val_out <= 4'h0393;
         4'hc9aa 	:	val_out <= 4'h0393;
         4'hc9ab 	:	val_out <= 4'h0393;
         4'hc9b0 	:	val_out <= 4'h0399;
         4'hc9b1 	:	val_out <= 4'h0399;
         4'hc9b2 	:	val_out <= 4'h0399;
         4'hc9b3 	:	val_out <= 4'h0399;
         4'hc9b8 	:	val_out <= 4'h039f;
         4'hc9b9 	:	val_out <= 4'h039f;
         4'hc9ba 	:	val_out <= 4'h039f;
         4'hc9bb 	:	val_out <= 4'h039f;
         4'hc9c0 	:	val_out <= 4'h03a5;
         4'hc9c1 	:	val_out <= 4'h03a5;
         4'hc9c2 	:	val_out <= 4'h03a5;
         4'hc9c3 	:	val_out <= 4'h03a5;
         4'hc9c8 	:	val_out <= 4'h03ab;
         4'hc9c9 	:	val_out <= 4'h03ab;
         4'hc9ca 	:	val_out <= 4'h03ab;
         4'hc9cb 	:	val_out <= 4'h03ab;
         4'hc9d0 	:	val_out <= 4'h03b1;
         4'hc9d1 	:	val_out <= 4'h03b1;
         4'hc9d2 	:	val_out <= 4'h03b1;
         4'hc9d3 	:	val_out <= 4'h03b1;
         4'hc9d8 	:	val_out <= 4'h03b7;
         4'hc9d9 	:	val_out <= 4'h03b7;
         4'hc9da 	:	val_out <= 4'h03b7;
         4'hc9db 	:	val_out <= 4'h03b7;
         4'hc9e0 	:	val_out <= 4'h03bd;
         4'hc9e1 	:	val_out <= 4'h03bd;
         4'hc9e2 	:	val_out <= 4'h03bd;
         4'hc9e3 	:	val_out <= 4'h03bd;
         4'hc9e8 	:	val_out <= 4'h03c3;
         4'hc9e9 	:	val_out <= 4'h03c3;
         4'hc9ea 	:	val_out <= 4'h03c3;
         4'hc9eb 	:	val_out <= 4'h03c3;
         4'hc9f0 	:	val_out <= 4'h03c9;
         4'hc9f1 	:	val_out <= 4'h03c9;
         4'hc9f2 	:	val_out <= 4'h03c9;
         4'hc9f3 	:	val_out <= 4'h03c9;
         4'hc9f8 	:	val_out <= 4'h03cf;
         4'hc9f9 	:	val_out <= 4'h03cf;
         4'hc9fa 	:	val_out <= 4'h03cf;
         4'hc9fb 	:	val_out <= 4'h03cf;
         4'hca00 	:	val_out <= 4'h03d6;
         4'hca01 	:	val_out <= 4'h03d6;
         4'hca02 	:	val_out <= 4'h03d6;
         4'hca03 	:	val_out <= 4'h03d6;
         4'hca08 	:	val_out <= 4'h03dc;
         4'hca09 	:	val_out <= 4'h03dc;
         4'hca0a 	:	val_out <= 4'h03dc;
         4'hca0b 	:	val_out <= 4'h03dc;
         4'hca10 	:	val_out <= 4'h03e2;
         4'hca11 	:	val_out <= 4'h03e2;
         4'hca12 	:	val_out <= 4'h03e2;
         4'hca13 	:	val_out <= 4'h03e2;
         4'hca18 	:	val_out <= 4'h03e8;
         4'hca19 	:	val_out <= 4'h03e8;
         4'hca1a 	:	val_out <= 4'h03e8;
         4'hca1b 	:	val_out <= 4'h03e8;
         4'hca20 	:	val_out <= 4'h03ee;
         4'hca21 	:	val_out <= 4'h03ee;
         4'hca22 	:	val_out <= 4'h03ee;
         4'hca23 	:	val_out <= 4'h03ee;
         4'hca28 	:	val_out <= 4'h03f4;
         4'hca29 	:	val_out <= 4'h03f4;
         4'hca2a 	:	val_out <= 4'h03f4;
         4'hca2b 	:	val_out <= 4'h03f4;
         4'hca30 	:	val_out <= 4'h03fa;
         4'hca31 	:	val_out <= 4'h03fa;
         4'hca32 	:	val_out <= 4'h03fa;
         4'hca33 	:	val_out <= 4'h03fa;
         4'hca38 	:	val_out <= 4'h0401;
         4'hca39 	:	val_out <= 4'h0401;
         4'hca3a 	:	val_out <= 4'h0401;
         4'hca3b 	:	val_out <= 4'h0401;
         4'hca40 	:	val_out <= 4'h0407;
         4'hca41 	:	val_out <= 4'h0407;
         4'hca42 	:	val_out <= 4'h0407;
         4'hca43 	:	val_out <= 4'h0407;
         4'hca48 	:	val_out <= 4'h040d;
         4'hca49 	:	val_out <= 4'h040d;
         4'hca4a 	:	val_out <= 4'h040d;
         4'hca4b 	:	val_out <= 4'h040d;
         4'hca50 	:	val_out <= 4'h0414;
         4'hca51 	:	val_out <= 4'h0414;
         4'hca52 	:	val_out <= 4'h0414;
         4'hca53 	:	val_out <= 4'h0414;
         4'hca58 	:	val_out <= 4'h041a;
         4'hca59 	:	val_out <= 4'h041a;
         4'hca5a 	:	val_out <= 4'h041a;
         4'hca5b 	:	val_out <= 4'h041a;
         4'hca60 	:	val_out <= 4'h0420;
         4'hca61 	:	val_out <= 4'h0420;
         4'hca62 	:	val_out <= 4'h0420;
         4'hca63 	:	val_out <= 4'h0420;
         4'hca68 	:	val_out <= 4'h0426;
         4'hca69 	:	val_out <= 4'h0426;
         4'hca6a 	:	val_out <= 4'h0426;
         4'hca6b 	:	val_out <= 4'h0426;
         4'hca70 	:	val_out <= 4'h042d;
         4'hca71 	:	val_out <= 4'h042d;
         4'hca72 	:	val_out <= 4'h042d;
         4'hca73 	:	val_out <= 4'h042d;
         4'hca78 	:	val_out <= 4'h0433;
         4'hca79 	:	val_out <= 4'h0433;
         4'hca7a 	:	val_out <= 4'h0433;
         4'hca7b 	:	val_out <= 4'h0433;
         4'hca80 	:	val_out <= 4'h043a;
         4'hca81 	:	val_out <= 4'h043a;
         4'hca82 	:	val_out <= 4'h043a;
         4'hca83 	:	val_out <= 4'h043a;
         4'hca88 	:	val_out <= 4'h0440;
         4'hca89 	:	val_out <= 4'h0440;
         4'hca8a 	:	val_out <= 4'h0440;
         4'hca8b 	:	val_out <= 4'h0440;
         4'hca90 	:	val_out <= 4'h0446;
         4'hca91 	:	val_out <= 4'h0446;
         4'hca92 	:	val_out <= 4'h0446;
         4'hca93 	:	val_out <= 4'h0446;
         4'hca98 	:	val_out <= 4'h044d;
         4'hca99 	:	val_out <= 4'h044d;
         4'hca9a 	:	val_out <= 4'h044d;
         4'hca9b 	:	val_out <= 4'h044d;
         4'hcaa0 	:	val_out <= 4'h0453;
         4'hcaa1 	:	val_out <= 4'h0453;
         4'hcaa2 	:	val_out <= 4'h0453;
         4'hcaa3 	:	val_out <= 4'h0453;
         4'hcaa8 	:	val_out <= 4'h045a;
         4'hcaa9 	:	val_out <= 4'h045a;
         4'hcaaa 	:	val_out <= 4'h045a;
         4'hcaab 	:	val_out <= 4'h045a;
         4'hcab0 	:	val_out <= 4'h0460;
         4'hcab1 	:	val_out <= 4'h0460;
         4'hcab2 	:	val_out <= 4'h0460;
         4'hcab3 	:	val_out <= 4'h0460;
         4'hcab8 	:	val_out <= 4'h0467;
         4'hcab9 	:	val_out <= 4'h0467;
         4'hcaba 	:	val_out <= 4'h0467;
         4'hcabb 	:	val_out <= 4'h0467;
         4'hcac0 	:	val_out <= 4'h046d;
         4'hcac1 	:	val_out <= 4'h046d;
         4'hcac2 	:	val_out <= 4'h046d;
         4'hcac3 	:	val_out <= 4'h046d;
         4'hcac8 	:	val_out <= 4'h0474;
         4'hcac9 	:	val_out <= 4'h0474;
         4'hcaca 	:	val_out <= 4'h0474;
         4'hcacb 	:	val_out <= 4'h0474;
         4'hcad0 	:	val_out <= 4'h047b;
         4'hcad1 	:	val_out <= 4'h047b;
         4'hcad2 	:	val_out <= 4'h047b;
         4'hcad3 	:	val_out <= 4'h047b;
         4'hcad8 	:	val_out <= 4'h0481;
         4'hcad9 	:	val_out <= 4'h0481;
         4'hcada 	:	val_out <= 4'h0481;
         4'hcadb 	:	val_out <= 4'h0481;
         4'hcae0 	:	val_out <= 4'h0488;
         4'hcae1 	:	val_out <= 4'h0488;
         4'hcae2 	:	val_out <= 4'h0488;
         4'hcae3 	:	val_out <= 4'h0488;
         4'hcae8 	:	val_out <= 4'h048e;
         4'hcae9 	:	val_out <= 4'h048e;
         4'hcaea 	:	val_out <= 4'h048e;
         4'hcaeb 	:	val_out <= 4'h048e;
         4'hcaf0 	:	val_out <= 4'h0495;
         4'hcaf1 	:	val_out <= 4'h0495;
         4'hcaf2 	:	val_out <= 4'h0495;
         4'hcaf3 	:	val_out <= 4'h0495;
         4'hcaf8 	:	val_out <= 4'h049c;
         4'hcaf9 	:	val_out <= 4'h049c;
         4'hcafa 	:	val_out <= 4'h049c;
         4'hcafb 	:	val_out <= 4'h049c;
         4'hcb00 	:	val_out <= 4'h04a2;
         4'hcb01 	:	val_out <= 4'h04a2;
         4'hcb02 	:	val_out <= 4'h04a2;
         4'hcb03 	:	val_out <= 4'h04a2;
         4'hcb08 	:	val_out <= 4'h04a9;
         4'hcb09 	:	val_out <= 4'h04a9;
         4'hcb0a 	:	val_out <= 4'h04a9;
         4'hcb0b 	:	val_out <= 4'h04a9;
         4'hcb10 	:	val_out <= 4'h04b0;
         4'hcb11 	:	val_out <= 4'h04b0;
         4'hcb12 	:	val_out <= 4'h04b0;
         4'hcb13 	:	val_out <= 4'h04b0;
         4'hcb18 	:	val_out <= 4'h04b7;
         4'hcb19 	:	val_out <= 4'h04b7;
         4'hcb1a 	:	val_out <= 4'h04b7;
         4'hcb1b 	:	val_out <= 4'h04b7;
         4'hcb20 	:	val_out <= 4'h04bd;
         4'hcb21 	:	val_out <= 4'h04bd;
         4'hcb22 	:	val_out <= 4'h04bd;
         4'hcb23 	:	val_out <= 4'h04bd;
         4'hcb28 	:	val_out <= 4'h04c4;
         4'hcb29 	:	val_out <= 4'h04c4;
         4'hcb2a 	:	val_out <= 4'h04c4;
         4'hcb2b 	:	val_out <= 4'h04c4;
         4'hcb30 	:	val_out <= 4'h04cb;
         4'hcb31 	:	val_out <= 4'h04cb;
         4'hcb32 	:	val_out <= 4'h04cb;
         4'hcb33 	:	val_out <= 4'h04cb;
         4'hcb38 	:	val_out <= 4'h04d2;
         4'hcb39 	:	val_out <= 4'h04d2;
         4'hcb3a 	:	val_out <= 4'h04d2;
         4'hcb3b 	:	val_out <= 4'h04d2;
         4'hcb40 	:	val_out <= 4'h04d9;
         4'hcb41 	:	val_out <= 4'h04d9;
         4'hcb42 	:	val_out <= 4'h04d9;
         4'hcb43 	:	val_out <= 4'h04d9;
         4'hcb48 	:	val_out <= 4'h04e0;
         4'hcb49 	:	val_out <= 4'h04e0;
         4'hcb4a 	:	val_out <= 4'h04e0;
         4'hcb4b 	:	val_out <= 4'h04e0;
         4'hcb50 	:	val_out <= 4'h04e6;
         4'hcb51 	:	val_out <= 4'h04e6;
         4'hcb52 	:	val_out <= 4'h04e6;
         4'hcb53 	:	val_out <= 4'h04e6;
         4'hcb58 	:	val_out <= 4'h04ed;
         4'hcb59 	:	val_out <= 4'h04ed;
         4'hcb5a 	:	val_out <= 4'h04ed;
         4'hcb5b 	:	val_out <= 4'h04ed;
         4'hcb60 	:	val_out <= 4'h04f4;
         4'hcb61 	:	val_out <= 4'h04f4;
         4'hcb62 	:	val_out <= 4'h04f4;
         4'hcb63 	:	val_out <= 4'h04f4;
         4'hcb68 	:	val_out <= 4'h04fb;
         4'hcb69 	:	val_out <= 4'h04fb;
         4'hcb6a 	:	val_out <= 4'h04fb;
         4'hcb6b 	:	val_out <= 4'h04fb;
         4'hcb70 	:	val_out <= 4'h0502;
         4'hcb71 	:	val_out <= 4'h0502;
         4'hcb72 	:	val_out <= 4'h0502;
         4'hcb73 	:	val_out <= 4'h0502;
         4'hcb78 	:	val_out <= 4'h0509;
         4'hcb79 	:	val_out <= 4'h0509;
         4'hcb7a 	:	val_out <= 4'h0509;
         4'hcb7b 	:	val_out <= 4'h0509;
         4'hcb80 	:	val_out <= 4'h0510;
         4'hcb81 	:	val_out <= 4'h0510;
         4'hcb82 	:	val_out <= 4'h0510;
         4'hcb83 	:	val_out <= 4'h0510;
         4'hcb88 	:	val_out <= 4'h0517;
         4'hcb89 	:	val_out <= 4'h0517;
         4'hcb8a 	:	val_out <= 4'h0517;
         4'hcb8b 	:	val_out <= 4'h0517;
         4'hcb90 	:	val_out <= 4'h051e;
         4'hcb91 	:	val_out <= 4'h051e;
         4'hcb92 	:	val_out <= 4'h051e;
         4'hcb93 	:	val_out <= 4'h051e;
         4'hcb98 	:	val_out <= 4'h0525;
         4'hcb99 	:	val_out <= 4'h0525;
         4'hcb9a 	:	val_out <= 4'h0525;
         4'hcb9b 	:	val_out <= 4'h0525;
         4'hcba0 	:	val_out <= 4'h052c;
         4'hcba1 	:	val_out <= 4'h052c;
         4'hcba2 	:	val_out <= 4'h052c;
         4'hcba3 	:	val_out <= 4'h052c;
         4'hcba8 	:	val_out <= 4'h0533;
         4'hcba9 	:	val_out <= 4'h0533;
         4'hcbaa 	:	val_out <= 4'h0533;
         4'hcbab 	:	val_out <= 4'h0533;
         4'hcbb0 	:	val_out <= 4'h053a;
         4'hcbb1 	:	val_out <= 4'h053a;
         4'hcbb2 	:	val_out <= 4'h053a;
         4'hcbb3 	:	val_out <= 4'h053a;
         4'hcbb8 	:	val_out <= 4'h0542;
         4'hcbb9 	:	val_out <= 4'h0542;
         4'hcbba 	:	val_out <= 4'h0542;
         4'hcbbb 	:	val_out <= 4'h0542;
         4'hcbc0 	:	val_out <= 4'h0549;
         4'hcbc1 	:	val_out <= 4'h0549;
         4'hcbc2 	:	val_out <= 4'h0549;
         4'hcbc3 	:	val_out <= 4'h0549;
         4'hcbc8 	:	val_out <= 4'h0550;
         4'hcbc9 	:	val_out <= 4'h0550;
         4'hcbca 	:	val_out <= 4'h0550;
         4'hcbcb 	:	val_out <= 4'h0550;
         4'hcbd0 	:	val_out <= 4'h0557;
         4'hcbd1 	:	val_out <= 4'h0557;
         4'hcbd2 	:	val_out <= 4'h0557;
         4'hcbd3 	:	val_out <= 4'h0557;
         4'hcbd8 	:	val_out <= 4'h055e;
         4'hcbd9 	:	val_out <= 4'h055e;
         4'hcbda 	:	val_out <= 4'h055e;
         4'hcbdb 	:	val_out <= 4'h055e;
         4'hcbe0 	:	val_out <= 4'h0565;
         4'hcbe1 	:	val_out <= 4'h0565;
         4'hcbe2 	:	val_out <= 4'h0565;
         4'hcbe3 	:	val_out <= 4'h0565;
         4'hcbe8 	:	val_out <= 4'h056d;
         4'hcbe9 	:	val_out <= 4'h056d;
         4'hcbea 	:	val_out <= 4'h056d;
         4'hcbeb 	:	val_out <= 4'h056d;
         4'hcbf0 	:	val_out <= 4'h0574;
         4'hcbf1 	:	val_out <= 4'h0574;
         4'hcbf2 	:	val_out <= 4'h0574;
         4'hcbf3 	:	val_out <= 4'h0574;
         4'hcbf8 	:	val_out <= 4'h057b;
         4'hcbf9 	:	val_out <= 4'h057b;
         4'hcbfa 	:	val_out <= 4'h057b;
         4'hcbfb 	:	val_out <= 4'h057b;
         4'hcc00 	:	val_out <= 4'h0582;
         4'hcc01 	:	val_out <= 4'h0582;
         4'hcc02 	:	val_out <= 4'h0582;
         4'hcc03 	:	val_out <= 4'h0582;
         4'hcc08 	:	val_out <= 4'h058a;
         4'hcc09 	:	val_out <= 4'h058a;
         4'hcc0a 	:	val_out <= 4'h058a;
         4'hcc0b 	:	val_out <= 4'h058a;
         4'hcc10 	:	val_out <= 4'h0591;
         4'hcc11 	:	val_out <= 4'h0591;
         4'hcc12 	:	val_out <= 4'h0591;
         4'hcc13 	:	val_out <= 4'h0591;
         4'hcc18 	:	val_out <= 4'h0598;
         4'hcc19 	:	val_out <= 4'h0598;
         4'hcc1a 	:	val_out <= 4'h0598;
         4'hcc1b 	:	val_out <= 4'h0598;
         4'hcc20 	:	val_out <= 4'h05a0;
         4'hcc21 	:	val_out <= 4'h05a0;
         4'hcc22 	:	val_out <= 4'h05a0;
         4'hcc23 	:	val_out <= 4'h05a0;
         4'hcc28 	:	val_out <= 4'h05a7;
         4'hcc29 	:	val_out <= 4'h05a7;
         4'hcc2a 	:	val_out <= 4'h05a7;
         4'hcc2b 	:	val_out <= 4'h05a7;
         4'hcc30 	:	val_out <= 4'h05af;
         4'hcc31 	:	val_out <= 4'h05af;
         4'hcc32 	:	val_out <= 4'h05af;
         4'hcc33 	:	val_out <= 4'h05af;
         4'hcc38 	:	val_out <= 4'h05b6;
         4'hcc39 	:	val_out <= 4'h05b6;
         4'hcc3a 	:	val_out <= 4'h05b6;
         4'hcc3b 	:	val_out <= 4'h05b6;
         4'hcc40 	:	val_out <= 4'h05bd;
         4'hcc41 	:	val_out <= 4'h05bd;
         4'hcc42 	:	val_out <= 4'h05bd;
         4'hcc43 	:	val_out <= 4'h05bd;
         4'hcc48 	:	val_out <= 4'h05c5;
         4'hcc49 	:	val_out <= 4'h05c5;
         4'hcc4a 	:	val_out <= 4'h05c5;
         4'hcc4b 	:	val_out <= 4'h05c5;
         4'hcc50 	:	val_out <= 4'h05cc;
         4'hcc51 	:	val_out <= 4'h05cc;
         4'hcc52 	:	val_out <= 4'h05cc;
         4'hcc53 	:	val_out <= 4'h05cc;
         4'hcc58 	:	val_out <= 4'h05d4;
         4'hcc59 	:	val_out <= 4'h05d4;
         4'hcc5a 	:	val_out <= 4'h05d4;
         4'hcc5b 	:	val_out <= 4'h05d4;
         4'hcc60 	:	val_out <= 4'h05db;
         4'hcc61 	:	val_out <= 4'h05db;
         4'hcc62 	:	val_out <= 4'h05db;
         4'hcc63 	:	val_out <= 4'h05db;
         4'hcc68 	:	val_out <= 4'h05e3;
         4'hcc69 	:	val_out <= 4'h05e3;
         4'hcc6a 	:	val_out <= 4'h05e3;
         4'hcc6b 	:	val_out <= 4'h05e3;
         4'hcc70 	:	val_out <= 4'h05ea;
         4'hcc71 	:	val_out <= 4'h05ea;
         4'hcc72 	:	val_out <= 4'h05ea;
         4'hcc73 	:	val_out <= 4'h05ea;
         4'hcc78 	:	val_out <= 4'h05f2;
         4'hcc79 	:	val_out <= 4'h05f2;
         4'hcc7a 	:	val_out <= 4'h05f2;
         4'hcc7b 	:	val_out <= 4'h05f2;
         4'hcc80 	:	val_out <= 4'h05fa;
         4'hcc81 	:	val_out <= 4'h05fa;
         4'hcc82 	:	val_out <= 4'h05fa;
         4'hcc83 	:	val_out <= 4'h05fa;
         4'hcc88 	:	val_out <= 4'h0601;
         4'hcc89 	:	val_out <= 4'h0601;
         4'hcc8a 	:	val_out <= 4'h0601;
         4'hcc8b 	:	val_out <= 4'h0601;
         4'hcc90 	:	val_out <= 4'h0609;
         4'hcc91 	:	val_out <= 4'h0609;
         4'hcc92 	:	val_out <= 4'h0609;
         4'hcc93 	:	val_out <= 4'h0609;
         4'hcc98 	:	val_out <= 4'h0610;
         4'hcc99 	:	val_out <= 4'h0610;
         4'hcc9a 	:	val_out <= 4'h0610;
         4'hcc9b 	:	val_out <= 4'h0610;
         4'hcca0 	:	val_out <= 4'h0618;
         4'hcca1 	:	val_out <= 4'h0618;
         4'hcca2 	:	val_out <= 4'h0618;
         4'hcca3 	:	val_out <= 4'h0618;
         4'hcca8 	:	val_out <= 4'h0620;
         4'hcca9 	:	val_out <= 4'h0620;
         4'hccaa 	:	val_out <= 4'h0620;
         4'hccab 	:	val_out <= 4'h0620;
         4'hccb0 	:	val_out <= 4'h0627;
         4'hccb1 	:	val_out <= 4'h0627;
         4'hccb2 	:	val_out <= 4'h0627;
         4'hccb3 	:	val_out <= 4'h0627;
         4'hccb8 	:	val_out <= 4'h062f;
         4'hccb9 	:	val_out <= 4'h062f;
         4'hccba 	:	val_out <= 4'h062f;
         4'hccbb 	:	val_out <= 4'h062f;
         4'hccc0 	:	val_out <= 4'h0637;
         4'hccc1 	:	val_out <= 4'h0637;
         4'hccc2 	:	val_out <= 4'h0637;
         4'hccc3 	:	val_out <= 4'h0637;
         4'hccc8 	:	val_out <= 4'h063f;
         4'hccc9 	:	val_out <= 4'h063f;
         4'hccca 	:	val_out <= 4'h063f;
         4'hcccb 	:	val_out <= 4'h063f;
         4'hccd0 	:	val_out <= 4'h0646;
         4'hccd1 	:	val_out <= 4'h0646;
         4'hccd2 	:	val_out <= 4'h0646;
         4'hccd3 	:	val_out <= 4'h0646;
         4'hccd8 	:	val_out <= 4'h064e;
         4'hccd9 	:	val_out <= 4'h064e;
         4'hccda 	:	val_out <= 4'h064e;
         4'hccdb 	:	val_out <= 4'h064e;
         4'hcce0 	:	val_out <= 4'h0656;
         4'hcce1 	:	val_out <= 4'h0656;
         4'hcce2 	:	val_out <= 4'h0656;
         4'hcce3 	:	val_out <= 4'h0656;
         4'hcce8 	:	val_out <= 4'h065e;
         4'hcce9 	:	val_out <= 4'h065e;
         4'hccea 	:	val_out <= 4'h065e;
         4'hcceb 	:	val_out <= 4'h065e;
         4'hccf0 	:	val_out <= 4'h0666;
         4'hccf1 	:	val_out <= 4'h0666;
         4'hccf2 	:	val_out <= 4'h0666;
         4'hccf3 	:	val_out <= 4'h0666;
         4'hccf8 	:	val_out <= 4'h066d;
         4'hccf9 	:	val_out <= 4'h066d;
         4'hccfa 	:	val_out <= 4'h066d;
         4'hccfb 	:	val_out <= 4'h066d;
         4'hcd00 	:	val_out <= 4'h0675;
         4'hcd01 	:	val_out <= 4'h0675;
         4'hcd02 	:	val_out <= 4'h0675;
         4'hcd03 	:	val_out <= 4'h0675;
         4'hcd08 	:	val_out <= 4'h067d;
         4'hcd09 	:	val_out <= 4'h067d;
         4'hcd0a 	:	val_out <= 4'h067d;
         4'hcd0b 	:	val_out <= 4'h067d;
         4'hcd10 	:	val_out <= 4'h0685;
         4'hcd11 	:	val_out <= 4'h0685;
         4'hcd12 	:	val_out <= 4'h0685;
         4'hcd13 	:	val_out <= 4'h0685;
         4'hcd18 	:	val_out <= 4'h068d;
         4'hcd19 	:	val_out <= 4'h068d;
         4'hcd1a 	:	val_out <= 4'h068d;
         4'hcd1b 	:	val_out <= 4'h068d;
         4'hcd20 	:	val_out <= 4'h0695;
         4'hcd21 	:	val_out <= 4'h0695;
         4'hcd22 	:	val_out <= 4'h0695;
         4'hcd23 	:	val_out <= 4'h0695;
         4'hcd28 	:	val_out <= 4'h069d;
         4'hcd29 	:	val_out <= 4'h069d;
         4'hcd2a 	:	val_out <= 4'h069d;
         4'hcd2b 	:	val_out <= 4'h069d;
         4'hcd30 	:	val_out <= 4'h06a5;
         4'hcd31 	:	val_out <= 4'h06a5;
         4'hcd32 	:	val_out <= 4'h06a5;
         4'hcd33 	:	val_out <= 4'h06a5;
         4'hcd38 	:	val_out <= 4'h06ad;
         4'hcd39 	:	val_out <= 4'h06ad;
         4'hcd3a 	:	val_out <= 4'h06ad;
         4'hcd3b 	:	val_out <= 4'h06ad;
         4'hcd40 	:	val_out <= 4'h06b5;
         4'hcd41 	:	val_out <= 4'h06b5;
         4'hcd42 	:	val_out <= 4'h06b5;
         4'hcd43 	:	val_out <= 4'h06b5;
         4'hcd48 	:	val_out <= 4'h06bd;
         4'hcd49 	:	val_out <= 4'h06bd;
         4'hcd4a 	:	val_out <= 4'h06bd;
         4'hcd4b 	:	val_out <= 4'h06bd;
         4'hcd50 	:	val_out <= 4'h06c5;
         4'hcd51 	:	val_out <= 4'h06c5;
         4'hcd52 	:	val_out <= 4'h06c5;
         4'hcd53 	:	val_out <= 4'h06c5;
         4'hcd58 	:	val_out <= 4'h06cd;
         4'hcd59 	:	val_out <= 4'h06cd;
         4'hcd5a 	:	val_out <= 4'h06cd;
         4'hcd5b 	:	val_out <= 4'h06cd;
         4'hcd60 	:	val_out <= 4'h06d5;
         4'hcd61 	:	val_out <= 4'h06d5;
         4'hcd62 	:	val_out <= 4'h06d5;
         4'hcd63 	:	val_out <= 4'h06d5;
         4'hcd68 	:	val_out <= 4'h06dd;
         4'hcd69 	:	val_out <= 4'h06dd;
         4'hcd6a 	:	val_out <= 4'h06dd;
         4'hcd6b 	:	val_out <= 4'h06dd;
         4'hcd70 	:	val_out <= 4'h06e6;
         4'hcd71 	:	val_out <= 4'h06e6;
         4'hcd72 	:	val_out <= 4'h06e6;
         4'hcd73 	:	val_out <= 4'h06e6;
         4'hcd78 	:	val_out <= 4'h06ee;
         4'hcd79 	:	val_out <= 4'h06ee;
         4'hcd7a 	:	val_out <= 4'h06ee;
         4'hcd7b 	:	val_out <= 4'h06ee;
         4'hcd80 	:	val_out <= 4'h06f6;
         4'hcd81 	:	val_out <= 4'h06f6;
         4'hcd82 	:	val_out <= 4'h06f6;
         4'hcd83 	:	val_out <= 4'h06f6;
         4'hcd88 	:	val_out <= 4'h06fe;
         4'hcd89 	:	val_out <= 4'h06fe;
         4'hcd8a 	:	val_out <= 4'h06fe;
         4'hcd8b 	:	val_out <= 4'h06fe;
         4'hcd90 	:	val_out <= 4'h0706;
         4'hcd91 	:	val_out <= 4'h0706;
         4'hcd92 	:	val_out <= 4'h0706;
         4'hcd93 	:	val_out <= 4'h0706;
         4'hcd98 	:	val_out <= 4'h070e;
         4'hcd99 	:	val_out <= 4'h070e;
         4'hcd9a 	:	val_out <= 4'h070e;
         4'hcd9b 	:	val_out <= 4'h070e;
         4'hcda0 	:	val_out <= 4'h0717;
         4'hcda1 	:	val_out <= 4'h0717;
         4'hcda2 	:	val_out <= 4'h0717;
         4'hcda3 	:	val_out <= 4'h0717;
         4'hcda8 	:	val_out <= 4'h071f;
         4'hcda9 	:	val_out <= 4'h071f;
         4'hcdaa 	:	val_out <= 4'h071f;
         4'hcdab 	:	val_out <= 4'h071f;
         4'hcdb0 	:	val_out <= 4'h0727;
         4'hcdb1 	:	val_out <= 4'h0727;
         4'hcdb2 	:	val_out <= 4'h0727;
         4'hcdb3 	:	val_out <= 4'h0727;
         4'hcdb8 	:	val_out <= 4'h0730;
         4'hcdb9 	:	val_out <= 4'h0730;
         4'hcdba 	:	val_out <= 4'h0730;
         4'hcdbb 	:	val_out <= 4'h0730;
         4'hcdc0 	:	val_out <= 4'h0738;
         4'hcdc1 	:	val_out <= 4'h0738;
         4'hcdc2 	:	val_out <= 4'h0738;
         4'hcdc3 	:	val_out <= 4'h0738;
         4'hcdc8 	:	val_out <= 4'h0740;
         4'hcdc9 	:	val_out <= 4'h0740;
         4'hcdca 	:	val_out <= 4'h0740;
         4'hcdcb 	:	val_out <= 4'h0740;
         4'hcdd0 	:	val_out <= 4'h0749;
         4'hcdd1 	:	val_out <= 4'h0749;
         4'hcdd2 	:	val_out <= 4'h0749;
         4'hcdd3 	:	val_out <= 4'h0749;
         4'hcdd8 	:	val_out <= 4'h0751;
         4'hcdd9 	:	val_out <= 4'h0751;
         4'hcdda 	:	val_out <= 4'h0751;
         4'hcddb 	:	val_out <= 4'h0751;
         4'hcde0 	:	val_out <= 4'h0759;
         4'hcde1 	:	val_out <= 4'h0759;
         4'hcde2 	:	val_out <= 4'h0759;
         4'hcde3 	:	val_out <= 4'h0759;
         4'hcde8 	:	val_out <= 4'h0762;
         4'hcde9 	:	val_out <= 4'h0762;
         4'hcdea 	:	val_out <= 4'h0762;
         4'hcdeb 	:	val_out <= 4'h0762;
         4'hcdf0 	:	val_out <= 4'h076a;
         4'hcdf1 	:	val_out <= 4'h076a;
         4'hcdf2 	:	val_out <= 4'h076a;
         4'hcdf3 	:	val_out <= 4'h076a;
         4'hcdf8 	:	val_out <= 4'h0773;
         4'hcdf9 	:	val_out <= 4'h0773;
         4'hcdfa 	:	val_out <= 4'h0773;
         4'hcdfb 	:	val_out <= 4'h0773;
         4'hce00 	:	val_out <= 4'h077b;
         4'hce01 	:	val_out <= 4'h077b;
         4'hce02 	:	val_out <= 4'h077b;
         4'hce03 	:	val_out <= 4'h077b;
         4'hce08 	:	val_out <= 4'h0783;
         4'hce09 	:	val_out <= 4'h0783;
         4'hce0a 	:	val_out <= 4'h0783;
         4'hce0b 	:	val_out <= 4'h0783;
         4'hce10 	:	val_out <= 4'h078c;
         4'hce11 	:	val_out <= 4'h078c;
         4'hce12 	:	val_out <= 4'h078c;
         4'hce13 	:	val_out <= 4'h078c;
         4'hce18 	:	val_out <= 4'h0794;
         4'hce19 	:	val_out <= 4'h0794;
         4'hce1a 	:	val_out <= 4'h0794;
         4'hce1b 	:	val_out <= 4'h0794;
         4'hce20 	:	val_out <= 4'h079d;
         4'hce21 	:	val_out <= 4'h079d;
         4'hce22 	:	val_out <= 4'h079d;
         4'hce23 	:	val_out <= 4'h079d;
         4'hce28 	:	val_out <= 4'h07a6;
         4'hce29 	:	val_out <= 4'h07a6;
         4'hce2a 	:	val_out <= 4'h07a6;
         4'hce2b 	:	val_out <= 4'h07a6;
         4'hce30 	:	val_out <= 4'h07ae;
         4'hce31 	:	val_out <= 4'h07ae;
         4'hce32 	:	val_out <= 4'h07ae;
         4'hce33 	:	val_out <= 4'h07ae;
         4'hce38 	:	val_out <= 4'h07b7;
         4'hce39 	:	val_out <= 4'h07b7;
         4'hce3a 	:	val_out <= 4'h07b7;
         4'hce3b 	:	val_out <= 4'h07b7;
         4'hce40 	:	val_out <= 4'h07bf;
         4'hce41 	:	val_out <= 4'h07bf;
         4'hce42 	:	val_out <= 4'h07bf;
         4'hce43 	:	val_out <= 4'h07bf;
         4'hce48 	:	val_out <= 4'h07c8;
         4'hce49 	:	val_out <= 4'h07c8;
         4'hce4a 	:	val_out <= 4'h07c8;
         4'hce4b 	:	val_out <= 4'h07c8;
         4'hce50 	:	val_out <= 4'h07d1;
         4'hce51 	:	val_out <= 4'h07d1;
         4'hce52 	:	val_out <= 4'h07d1;
         4'hce53 	:	val_out <= 4'h07d1;
         4'hce58 	:	val_out <= 4'h07d9;
         4'hce59 	:	val_out <= 4'h07d9;
         4'hce5a 	:	val_out <= 4'h07d9;
         4'hce5b 	:	val_out <= 4'h07d9;
         4'hce60 	:	val_out <= 4'h07e2;
         4'hce61 	:	val_out <= 4'h07e2;
         4'hce62 	:	val_out <= 4'h07e2;
         4'hce63 	:	val_out <= 4'h07e2;
         4'hce68 	:	val_out <= 4'h07eb;
         4'hce69 	:	val_out <= 4'h07eb;
         4'hce6a 	:	val_out <= 4'h07eb;
         4'hce6b 	:	val_out <= 4'h07eb;
         4'hce70 	:	val_out <= 4'h07f3;
         4'hce71 	:	val_out <= 4'h07f3;
         4'hce72 	:	val_out <= 4'h07f3;
         4'hce73 	:	val_out <= 4'h07f3;
         4'hce78 	:	val_out <= 4'h07fc;
         4'hce79 	:	val_out <= 4'h07fc;
         4'hce7a 	:	val_out <= 4'h07fc;
         4'hce7b 	:	val_out <= 4'h07fc;
         4'hce80 	:	val_out <= 4'h0805;
         4'hce81 	:	val_out <= 4'h0805;
         4'hce82 	:	val_out <= 4'h0805;
         4'hce83 	:	val_out <= 4'h0805;
         4'hce88 	:	val_out <= 4'h080e;
         4'hce89 	:	val_out <= 4'h080e;
         4'hce8a 	:	val_out <= 4'h080e;
         4'hce8b 	:	val_out <= 4'h080e;
         4'hce90 	:	val_out <= 4'h0816;
         4'hce91 	:	val_out <= 4'h0816;
         4'hce92 	:	val_out <= 4'h0816;
         4'hce93 	:	val_out <= 4'h0816;
         4'hce98 	:	val_out <= 4'h081f;
         4'hce99 	:	val_out <= 4'h081f;
         4'hce9a 	:	val_out <= 4'h081f;
         4'hce9b 	:	val_out <= 4'h081f;
         4'hcea0 	:	val_out <= 4'h0828;
         4'hcea1 	:	val_out <= 4'h0828;
         4'hcea2 	:	val_out <= 4'h0828;
         4'hcea3 	:	val_out <= 4'h0828;
         4'hcea8 	:	val_out <= 4'h0831;
         4'hcea9 	:	val_out <= 4'h0831;
         4'hceaa 	:	val_out <= 4'h0831;
         4'hceab 	:	val_out <= 4'h0831;
         4'hceb0 	:	val_out <= 4'h083a;
         4'hceb1 	:	val_out <= 4'h083a;
         4'hceb2 	:	val_out <= 4'h083a;
         4'hceb3 	:	val_out <= 4'h083a;
         4'hceb8 	:	val_out <= 4'h0843;
         4'hceb9 	:	val_out <= 4'h0843;
         4'hceba 	:	val_out <= 4'h0843;
         4'hcebb 	:	val_out <= 4'h0843;
         4'hcec0 	:	val_out <= 4'h084b;
         4'hcec1 	:	val_out <= 4'h084b;
         4'hcec2 	:	val_out <= 4'h084b;
         4'hcec3 	:	val_out <= 4'h084b;
         4'hcec8 	:	val_out <= 4'h0854;
         4'hcec9 	:	val_out <= 4'h0854;
         4'hceca 	:	val_out <= 4'h0854;
         4'hcecb 	:	val_out <= 4'h0854;
         4'hced0 	:	val_out <= 4'h085d;
         4'hced1 	:	val_out <= 4'h085d;
         4'hced2 	:	val_out <= 4'h085d;
         4'hced3 	:	val_out <= 4'h085d;
         4'hced8 	:	val_out <= 4'h0866;
         4'hced9 	:	val_out <= 4'h0866;
         4'hceda 	:	val_out <= 4'h0866;
         4'hcedb 	:	val_out <= 4'h0866;
         4'hcee0 	:	val_out <= 4'h086f;
         4'hcee1 	:	val_out <= 4'h086f;
         4'hcee2 	:	val_out <= 4'h086f;
         4'hcee3 	:	val_out <= 4'h086f;
         4'hcee8 	:	val_out <= 4'h0878;
         4'hcee9 	:	val_out <= 4'h0878;
         4'hceea 	:	val_out <= 4'h0878;
         4'hceeb 	:	val_out <= 4'h0878;
         4'hcef0 	:	val_out <= 4'h0881;
         4'hcef1 	:	val_out <= 4'h0881;
         4'hcef2 	:	val_out <= 4'h0881;
         4'hcef3 	:	val_out <= 4'h0881;
         4'hcef8 	:	val_out <= 4'h088a;
         4'hcef9 	:	val_out <= 4'h088a;
         4'hcefa 	:	val_out <= 4'h088a;
         4'hcefb 	:	val_out <= 4'h088a;
         4'hcf00 	:	val_out <= 4'h0893;
         4'hcf01 	:	val_out <= 4'h0893;
         4'hcf02 	:	val_out <= 4'h0893;
         4'hcf03 	:	val_out <= 4'h0893;
         4'hcf08 	:	val_out <= 4'h089c;
         4'hcf09 	:	val_out <= 4'h089c;
         4'hcf0a 	:	val_out <= 4'h089c;
         4'hcf0b 	:	val_out <= 4'h089c;
         4'hcf10 	:	val_out <= 4'h08a5;
         4'hcf11 	:	val_out <= 4'h08a5;
         4'hcf12 	:	val_out <= 4'h08a5;
         4'hcf13 	:	val_out <= 4'h08a5;
         4'hcf18 	:	val_out <= 4'h08ae;
         4'hcf19 	:	val_out <= 4'h08ae;
         4'hcf1a 	:	val_out <= 4'h08ae;
         4'hcf1b 	:	val_out <= 4'h08ae;
         4'hcf20 	:	val_out <= 4'h08b8;
         4'hcf21 	:	val_out <= 4'h08b8;
         4'hcf22 	:	val_out <= 4'h08b8;
         4'hcf23 	:	val_out <= 4'h08b8;
         4'hcf28 	:	val_out <= 4'h08c1;
         4'hcf29 	:	val_out <= 4'h08c1;
         4'hcf2a 	:	val_out <= 4'h08c1;
         4'hcf2b 	:	val_out <= 4'h08c1;
         4'hcf30 	:	val_out <= 4'h08ca;
         4'hcf31 	:	val_out <= 4'h08ca;
         4'hcf32 	:	val_out <= 4'h08ca;
         4'hcf33 	:	val_out <= 4'h08ca;
         4'hcf38 	:	val_out <= 4'h08d3;
         4'hcf39 	:	val_out <= 4'h08d3;
         4'hcf3a 	:	val_out <= 4'h08d3;
         4'hcf3b 	:	val_out <= 4'h08d3;
         4'hcf40 	:	val_out <= 4'h08dc;
         4'hcf41 	:	val_out <= 4'h08dc;
         4'hcf42 	:	val_out <= 4'h08dc;
         4'hcf43 	:	val_out <= 4'h08dc;
         4'hcf48 	:	val_out <= 4'h08e5;
         4'hcf49 	:	val_out <= 4'h08e5;
         4'hcf4a 	:	val_out <= 4'h08e5;
         4'hcf4b 	:	val_out <= 4'h08e5;
         4'hcf50 	:	val_out <= 4'h08ef;
         4'hcf51 	:	val_out <= 4'h08ef;
         4'hcf52 	:	val_out <= 4'h08ef;
         4'hcf53 	:	val_out <= 4'h08ef;
         4'hcf58 	:	val_out <= 4'h08f8;
         4'hcf59 	:	val_out <= 4'h08f8;
         4'hcf5a 	:	val_out <= 4'h08f8;
         4'hcf5b 	:	val_out <= 4'h08f8;
         4'hcf60 	:	val_out <= 4'h0901;
         4'hcf61 	:	val_out <= 4'h0901;
         4'hcf62 	:	val_out <= 4'h0901;
         4'hcf63 	:	val_out <= 4'h0901;
         4'hcf68 	:	val_out <= 4'h090a;
         4'hcf69 	:	val_out <= 4'h090a;
         4'hcf6a 	:	val_out <= 4'h090a;
         4'hcf6b 	:	val_out <= 4'h090a;
         4'hcf70 	:	val_out <= 4'h0914;
         4'hcf71 	:	val_out <= 4'h0914;
         4'hcf72 	:	val_out <= 4'h0914;
         4'hcf73 	:	val_out <= 4'h0914;
         4'hcf78 	:	val_out <= 4'h091d;
         4'hcf79 	:	val_out <= 4'h091d;
         4'hcf7a 	:	val_out <= 4'h091d;
         4'hcf7b 	:	val_out <= 4'h091d;
         4'hcf80 	:	val_out <= 4'h0926;
         4'hcf81 	:	val_out <= 4'h0926;
         4'hcf82 	:	val_out <= 4'h0926;
         4'hcf83 	:	val_out <= 4'h0926;
         4'hcf88 	:	val_out <= 4'h0930;
         4'hcf89 	:	val_out <= 4'h0930;
         4'hcf8a 	:	val_out <= 4'h0930;
         4'hcf8b 	:	val_out <= 4'h0930;
         4'hcf90 	:	val_out <= 4'h0939;
         4'hcf91 	:	val_out <= 4'h0939;
         4'hcf92 	:	val_out <= 4'h0939;
         4'hcf93 	:	val_out <= 4'h0939;
         4'hcf98 	:	val_out <= 4'h0942;
         4'hcf99 	:	val_out <= 4'h0942;
         4'hcf9a 	:	val_out <= 4'h0942;
         4'hcf9b 	:	val_out <= 4'h0942;
         4'hcfa0 	:	val_out <= 4'h094c;
         4'hcfa1 	:	val_out <= 4'h094c;
         4'hcfa2 	:	val_out <= 4'h094c;
         4'hcfa3 	:	val_out <= 4'h094c;
         4'hcfa8 	:	val_out <= 4'h0955;
         4'hcfa9 	:	val_out <= 4'h0955;
         4'hcfaa 	:	val_out <= 4'h0955;
         4'hcfab 	:	val_out <= 4'h0955;
         4'hcfb0 	:	val_out <= 4'h095f;
         4'hcfb1 	:	val_out <= 4'h095f;
         4'hcfb2 	:	val_out <= 4'h095f;
         4'hcfb3 	:	val_out <= 4'h095f;
         4'hcfb8 	:	val_out <= 4'h0968;
         4'hcfb9 	:	val_out <= 4'h0968;
         4'hcfba 	:	val_out <= 4'h0968;
         4'hcfbb 	:	val_out <= 4'h0968;
         4'hcfc0 	:	val_out <= 4'h0971;
         4'hcfc1 	:	val_out <= 4'h0971;
         4'hcfc2 	:	val_out <= 4'h0971;
         4'hcfc3 	:	val_out <= 4'h0971;
         4'hcfc8 	:	val_out <= 4'h097b;
         4'hcfc9 	:	val_out <= 4'h097b;
         4'hcfca 	:	val_out <= 4'h097b;
         4'hcfcb 	:	val_out <= 4'h097b;
         4'hcfd0 	:	val_out <= 4'h0984;
         4'hcfd1 	:	val_out <= 4'h0984;
         4'hcfd2 	:	val_out <= 4'h0984;
         4'hcfd3 	:	val_out <= 4'h0984;
         4'hcfd8 	:	val_out <= 4'h098e;
         4'hcfd9 	:	val_out <= 4'h098e;
         4'hcfda 	:	val_out <= 4'h098e;
         4'hcfdb 	:	val_out <= 4'h098e;
         4'hcfe0 	:	val_out <= 4'h0997;
         4'hcfe1 	:	val_out <= 4'h0997;
         4'hcfe2 	:	val_out <= 4'h0997;
         4'hcfe3 	:	val_out <= 4'h0997;
         4'hcfe8 	:	val_out <= 4'h09a1;
         4'hcfe9 	:	val_out <= 4'h09a1;
         4'hcfea 	:	val_out <= 4'h09a1;
         4'hcfeb 	:	val_out <= 4'h09a1;
         4'hcff0 	:	val_out <= 4'h09ab;
         4'hcff1 	:	val_out <= 4'h09ab;
         4'hcff2 	:	val_out <= 4'h09ab;
         4'hcff3 	:	val_out <= 4'h09ab;
         4'hcff8 	:	val_out <= 4'h09b4;
         4'hcff9 	:	val_out <= 4'h09b4;
         4'hcffa 	:	val_out <= 4'h09b4;
         4'hcffb 	:	val_out <= 4'h09b4;
         4'hd000 	:	val_out <= 4'h09be;
         4'hd001 	:	val_out <= 4'h09be;
         4'hd002 	:	val_out <= 4'h09be;
         4'hd003 	:	val_out <= 4'h09be;
         4'hd008 	:	val_out <= 4'h09c7;
         4'hd009 	:	val_out <= 4'h09c7;
         4'hd00a 	:	val_out <= 4'h09c7;
         4'hd00b 	:	val_out <= 4'h09c7;
         4'hd010 	:	val_out <= 4'h09d1;
         4'hd011 	:	val_out <= 4'h09d1;
         4'hd012 	:	val_out <= 4'h09d1;
         4'hd013 	:	val_out <= 4'h09d1;
         4'hd018 	:	val_out <= 4'h09db;
         4'hd019 	:	val_out <= 4'h09db;
         4'hd01a 	:	val_out <= 4'h09db;
         4'hd01b 	:	val_out <= 4'h09db;
         4'hd020 	:	val_out <= 4'h09e4;
         4'hd021 	:	val_out <= 4'h09e4;
         4'hd022 	:	val_out <= 4'h09e4;
         4'hd023 	:	val_out <= 4'h09e4;
         4'hd028 	:	val_out <= 4'h09ee;
         4'hd029 	:	val_out <= 4'h09ee;
         4'hd02a 	:	val_out <= 4'h09ee;
         4'hd02b 	:	val_out <= 4'h09ee;
         4'hd030 	:	val_out <= 4'h09f8;
         4'hd031 	:	val_out <= 4'h09f8;
         4'hd032 	:	val_out <= 4'h09f8;
         4'hd033 	:	val_out <= 4'h09f8;
         4'hd038 	:	val_out <= 4'h0a02;
         4'hd039 	:	val_out <= 4'h0a02;
         4'hd03a 	:	val_out <= 4'h0a02;
         4'hd03b 	:	val_out <= 4'h0a02;
         4'hd040 	:	val_out <= 4'h0a0b;
         4'hd041 	:	val_out <= 4'h0a0b;
         4'hd042 	:	val_out <= 4'h0a0b;
         4'hd043 	:	val_out <= 4'h0a0b;
         4'hd048 	:	val_out <= 4'h0a15;
         4'hd049 	:	val_out <= 4'h0a15;
         4'hd04a 	:	val_out <= 4'h0a15;
         4'hd04b 	:	val_out <= 4'h0a15;
         4'hd050 	:	val_out <= 4'h0a1f;
         4'hd051 	:	val_out <= 4'h0a1f;
         4'hd052 	:	val_out <= 4'h0a1f;
         4'hd053 	:	val_out <= 4'h0a1f;
         4'hd058 	:	val_out <= 4'h0a29;
         4'hd059 	:	val_out <= 4'h0a29;
         4'hd05a 	:	val_out <= 4'h0a29;
         4'hd05b 	:	val_out <= 4'h0a29;
         4'hd060 	:	val_out <= 4'h0a33;
         4'hd061 	:	val_out <= 4'h0a33;
         4'hd062 	:	val_out <= 4'h0a33;
         4'hd063 	:	val_out <= 4'h0a33;
         4'hd068 	:	val_out <= 4'h0a3c;
         4'hd069 	:	val_out <= 4'h0a3c;
         4'hd06a 	:	val_out <= 4'h0a3c;
         4'hd06b 	:	val_out <= 4'h0a3c;
         4'hd070 	:	val_out <= 4'h0a46;
         4'hd071 	:	val_out <= 4'h0a46;
         4'hd072 	:	val_out <= 4'h0a46;
         4'hd073 	:	val_out <= 4'h0a46;
         4'hd078 	:	val_out <= 4'h0a50;
         4'hd079 	:	val_out <= 4'h0a50;
         4'hd07a 	:	val_out <= 4'h0a50;
         4'hd07b 	:	val_out <= 4'h0a50;
         4'hd080 	:	val_out <= 4'h0a5a;
         4'hd081 	:	val_out <= 4'h0a5a;
         4'hd082 	:	val_out <= 4'h0a5a;
         4'hd083 	:	val_out <= 4'h0a5a;
         4'hd088 	:	val_out <= 4'h0a64;
         4'hd089 	:	val_out <= 4'h0a64;
         4'hd08a 	:	val_out <= 4'h0a64;
         4'hd08b 	:	val_out <= 4'h0a64;
         4'hd090 	:	val_out <= 4'h0a6e;
         4'hd091 	:	val_out <= 4'h0a6e;
         4'hd092 	:	val_out <= 4'h0a6e;
         4'hd093 	:	val_out <= 4'h0a6e;
         4'hd098 	:	val_out <= 4'h0a78;
         4'hd099 	:	val_out <= 4'h0a78;
         4'hd09a 	:	val_out <= 4'h0a78;
         4'hd09b 	:	val_out <= 4'h0a78;
         4'hd0a0 	:	val_out <= 4'h0a82;
         4'hd0a1 	:	val_out <= 4'h0a82;
         4'hd0a2 	:	val_out <= 4'h0a82;
         4'hd0a3 	:	val_out <= 4'h0a82;
         4'hd0a8 	:	val_out <= 4'h0a8c;
         4'hd0a9 	:	val_out <= 4'h0a8c;
         4'hd0aa 	:	val_out <= 4'h0a8c;
         4'hd0ab 	:	val_out <= 4'h0a8c;
         4'hd0b0 	:	val_out <= 4'h0a96;
         4'hd0b1 	:	val_out <= 4'h0a96;
         4'hd0b2 	:	val_out <= 4'h0a96;
         4'hd0b3 	:	val_out <= 4'h0a96;
         4'hd0b8 	:	val_out <= 4'h0aa0;
         4'hd0b9 	:	val_out <= 4'h0aa0;
         4'hd0ba 	:	val_out <= 4'h0aa0;
         4'hd0bb 	:	val_out <= 4'h0aa0;
         4'hd0c0 	:	val_out <= 4'h0aaa;
         4'hd0c1 	:	val_out <= 4'h0aaa;
         4'hd0c2 	:	val_out <= 4'h0aaa;
         4'hd0c3 	:	val_out <= 4'h0aaa;
         4'hd0c8 	:	val_out <= 4'h0ab4;
         4'hd0c9 	:	val_out <= 4'h0ab4;
         4'hd0ca 	:	val_out <= 4'h0ab4;
         4'hd0cb 	:	val_out <= 4'h0ab4;
         4'hd0d0 	:	val_out <= 4'h0abe;
         4'hd0d1 	:	val_out <= 4'h0abe;
         4'hd0d2 	:	val_out <= 4'h0abe;
         4'hd0d3 	:	val_out <= 4'h0abe;
         4'hd0d8 	:	val_out <= 4'h0ac8;
         4'hd0d9 	:	val_out <= 4'h0ac8;
         4'hd0da 	:	val_out <= 4'h0ac8;
         4'hd0db 	:	val_out <= 4'h0ac8;
         4'hd0e0 	:	val_out <= 4'h0ad2;
         4'hd0e1 	:	val_out <= 4'h0ad2;
         4'hd0e2 	:	val_out <= 4'h0ad2;
         4'hd0e3 	:	val_out <= 4'h0ad2;
         4'hd0e8 	:	val_out <= 4'h0adc;
         4'hd0e9 	:	val_out <= 4'h0adc;
         4'hd0ea 	:	val_out <= 4'h0adc;
         4'hd0eb 	:	val_out <= 4'h0adc;
         4'hd0f0 	:	val_out <= 4'h0ae6;
         4'hd0f1 	:	val_out <= 4'h0ae6;
         4'hd0f2 	:	val_out <= 4'h0ae6;
         4'hd0f3 	:	val_out <= 4'h0ae6;
         4'hd0f8 	:	val_out <= 4'h0af0;
         4'hd0f9 	:	val_out <= 4'h0af0;
         4'hd0fa 	:	val_out <= 4'h0af0;
         4'hd0fb 	:	val_out <= 4'h0af0;
         4'hd100 	:	val_out <= 4'h0afb;
         4'hd101 	:	val_out <= 4'h0afb;
         4'hd102 	:	val_out <= 4'h0afb;
         4'hd103 	:	val_out <= 4'h0afb;
         4'hd108 	:	val_out <= 4'h0b05;
         4'hd109 	:	val_out <= 4'h0b05;
         4'hd10a 	:	val_out <= 4'h0b05;
         4'hd10b 	:	val_out <= 4'h0b05;
         4'hd110 	:	val_out <= 4'h0b0f;
         4'hd111 	:	val_out <= 4'h0b0f;
         4'hd112 	:	val_out <= 4'h0b0f;
         4'hd113 	:	val_out <= 4'h0b0f;
         4'hd118 	:	val_out <= 4'h0b19;
         4'hd119 	:	val_out <= 4'h0b19;
         4'hd11a 	:	val_out <= 4'h0b19;
         4'hd11b 	:	val_out <= 4'h0b19;
         4'hd120 	:	val_out <= 4'h0b24;
         4'hd121 	:	val_out <= 4'h0b24;
         4'hd122 	:	val_out <= 4'h0b24;
         4'hd123 	:	val_out <= 4'h0b24;
         4'hd128 	:	val_out <= 4'h0b2e;
         4'hd129 	:	val_out <= 4'h0b2e;
         4'hd12a 	:	val_out <= 4'h0b2e;
         4'hd12b 	:	val_out <= 4'h0b2e;
         4'hd130 	:	val_out <= 4'h0b38;
         4'hd131 	:	val_out <= 4'h0b38;
         4'hd132 	:	val_out <= 4'h0b38;
         4'hd133 	:	val_out <= 4'h0b38;
         4'hd138 	:	val_out <= 4'h0b42;
         4'hd139 	:	val_out <= 4'h0b42;
         4'hd13a 	:	val_out <= 4'h0b42;
         4'hd13b 	:	val_out <= 4'h0b42;
         4'hd140 	:	val_out <= 4'h0b4d;
         4'hd141 	:	val_out <= 4'h0b4d;
         4'hd142 	:	val_out <= 4'h0b4d;
         4'hd143 	:	val_out <= 4'h0b4d;
         4'hd148 	:	val_out <= 4'h0b57;
         4'hd149 	:	val_out <= 4'h0b57;
         4'hd14a 	:	val_out <= 4'h0b57;
         4'hd14b 	:	val_out <= 4'h0b57;
         4'hd150 	:	val_out <= 4'h0b61;
         4'hd151 	:	val_out <= 4'h0b61;
         4'hd152 	:	val_out <= 4'h0b61;
         4'hd153 	:	val_out <= 4'h0b61;
         4'hd158 	:	val_out <= 4'h0b6c;
         4'hd159 	:	val_out <= 4'h0b6c;
         4'hd15a 	:	val_out <= 4'h0b6c;
         4'hd15b 	:	val_out <= 4'h0b6c;
         4'hd160 	:	val_out <= 4'h0b76;
         4'hd161 	:	val_out <= 4'h0b76;
         4'hd162 	:	val_out <= 4'h0b76;
         4'hd163 	:	val_out <= 4'h0b76;
         4'hd168 	:	val_out <= 4'h0b81;
         4'hd169 	:	val_out <= 4'h0b81;
         4'hd16a 	:	val_out <= 4'h0b81;
         4'hd16b 	:	val_out <= 4'h0b81;
         4'hd170 	:	val_out <= 4'h0b8b;
         4'hd171 	:	val_out <= 4'h0b8b;
         4'hd172 	:	val_out <= 4'h0b8b;
         4'hd173 	:	val_out <= 4'h0b8b;
         4'hd178 	:	val_out <= 4'h0b95;
         4'hd179 	:	val_out <= 4'h0b95;
         4'hd17a 	:	val_out <= 4'h0b95;
         4'hd17b 	:	val_out <= 4'h0b95;
         4'hd180 	:	val_out <= 4'h0ba0;
         4'hd181 	:	val_out <= 4'h0ba0;
         4'hd182 	:	val_out <= 4'h0ba0;
         4'hd183 	:	val_out <= 4'h0ba0;
         4'hd188 	:	val_out <= 4'h0baa;
         4'hd189 	:	val_out <= 4'h0baa;
         4'hd18a 	:	val_out <= 4'h0baa;
         4'hd18b 	:	val_out <= 4'h0baa;
         4'hd190 	:	val_out <= 4'h0bb5;
         4'hd191 	:	val_out <= 4'h0bb5;
         4'hd192 	:	val_out <= 4'h0bb5;
         4'hd193 	:	val_out <= 4'h0bb5;
         4'hd198 	:	val_out <= 4'h0bbf;
         4'hd199 	:	val_out <= 4'h0bbf;
         4'hd19a 	:	val_out <= 4'h0bbf;
         4'hd19b 	:	val_out <= 4'h0bbf;
         4'hd1a0 	:	val_out <= 4'h0bca;
         4'hd1a1 	:	val_out <= 4'h0bca;
         4'hd1a2 	:	val_out <= 4'h0bca;
         4'hd1a3 	:	val_out <= 4'h0bca;
         4'hd1a8 	:	val_out <= 4'h0bd4;
         4'hd1a9 	:	val_out <= 4'h0bd4;
         4'hd1aa 	:	val_out <= 4'h0bd4;
         4'hd1ab 	:	val_out <= 4'h0bd4;
         4'hd1b0 	:	val_out <= 4'h0bdf;
         4'hd1b1 	:	val_out <= 4'h0bdf;
         4'hd1b2 	:	val_out <= 4'h0bdf;
         4'hd1b3 	:	val_out <= 4'h0bdf;
         4'hd1b8 	:	val_out <= 4'h0bea;
         4'hd1b9 	:	val_out <= 4'h0bea;
         4'hd1ba 	:	val_out <= 4'h0bea;
         4'hd1bb 	:	val_out <= 4'h0bea;
         4'hd1c0 	:	val_out <= 4'h0bf4;
         4'hd1c1 	:	val_out <= 4'h0bf4;
         4'hd1c2 	:	val_out <= 4'h0bf4;
         4'hd1c3 	:	val_out <= 4'h0bf4;
         4'hd1c8 	:	val_out <= 4'h0bff;
         4'hd1c9 	:	val_out <= 4'h0bff;
         4'hd1ca 	:	val_out <= 4'h0bff;
         4'hd1cb 	:	val_out <= 4'h0bff;
         4'hd1d0 	:	val_out <= 4'h0c09;
         4'hd1d1 	:	val_out <= 4'h0c09;
         4'hd1d2 	:	val_out <= 4'h0c09;
         4'hd1d3 	:	val_out <= 4'h0c09;
         4'hd1d8 	:	val_out <= 4'h0c14;
         4'hd1d9 	:	val_out <= 4'h0c14;
         4'hd1da 	:	val_out <= 4'h0c14;
         4'hd1db 	:	val_out <= 4'h0c14;
         4'hd1e0 	:	val_out <= 4'h0c1f;
         4'hd1e1 	:	val_out <= 4'h0c1f;
         4'hd1e2 	:	val_out <= 4'h0c1f;
         4'hd1e3 	:	val_out <= 4'h0c1f;
         4'hd1e8 	:	val_out <= 4'h0c29;
         4'hd1e9 	:	val_out <= 4'h0c29;
         4'hd1ea 	:	val_out <= 4'h0c29;
         4'hd1eb 	:	val_out <= 4'h0c29;
         4'hd1f0 	:	val_out <= 4'h0c34;
         4'hd1f1 	:	val_out <= 4'h0c34;
         4'hd1f2 	:	val_out <= 4'h0c34;
         4'hd1f3 	:	val_out <= 4'h0c34;
         4'hd1f8 	:	val_out <= 4'h0c3f;
         4'hd1f9 	:	val_out <= 4'h0c3f;
         4'hd1fa 	:	val_out <= 4'h0c3f;
         4'hd1fb 	:	val_out <= 4'h0c3f;
         4'hd200 	:	val_out <= 4'h0c4a;
         4'hd201 	:	val_out <= 4'h0c4a;
         4'hd202 	:	val_out <= 4'h0c4a;
         4'hd203 	:	val_out <= 4'h0c4a;
         4'hd208 	:	val_out <= 4'h0c54;
         4'hd209 	:	val_out <= 4'h0c54;
         4'hd20a 	:	val_out <= 4'h0c54;
         4'hd20b 	:	val_out <= 4'h0c54;
         4'hd210 	:	val_out <= 4'h0c5f;
         4'hd211 	:	val_out <= 4'h0c5f;
         4'hd212 	:	val_out <= 4'h0c5f;
         4'hd213 	:	val_out <= 4'h0c5f;
         4'hd218 	:	val_out <= 4'h0c6a;
         4'hd219 	:	val_out <= 4'h0c6a;
         4'hd21a 	:	val_out <= 4'h0c6a;
         4'hd21b 	:	val_out <= 4'h0c6a;
         4'hd220 	:	val_out <= 4'h0c75;
         4'hd221 	:	val_out <= 4'h0c75;
         4'hd222 	:	val_out <= 4'h0c75;
         4'hd223 	:	val_out <= 4'h0c75;
         4'hd228 	:	val_out <= 4'h0c80;
         4'hd229 	:	val_out <= 4'h0c80;
         4'hd22a 	:	val_out <= 4'h0c80;
         4'hd22b 	:	val_out <= 4'h0c80;
         4'hd230 	:	val_out <= 4'h0c8a;
         4'hd231 	:	val_out <= 4'h0c8a;
         4'hd232 	:	val_out <= 4'h0c8a;
         4'hd233 	:	val_out <= 4'h0c8a;
         4'hd238 	:	val_out <= 4'h0c95;
         4'hd239 	:	val_out <= 4'h0c95;
         4'hd23a 	:	val_out <= 4'h0c95;
         4'hd23b 	:	val_out <= 4'h0c95;
         4'hd240 	:	val_out <= 4'h0ca0;
         4'hd241 	:	val_out <= 4'h0ca0;
         4'hd242 	:	val_out <= 4'h0ca0;
         4'hd243 	:	val_out <= 4'h0ca0;
         4'hd248 	:	val_out <= 4'h0cab;
         4'hd249 	:	val_out <= 4'h0cab;
         4'hd24a 	:	val_out <= 4'h0cab;
         4'hd24b 	:	val_out <= 4'h0cab;
         4'hd250 	:	val_out <= 4'h0cb6;
         4'hd251 	:	val_out <= 4'h0cb6;
         4'hd252 	:	val_out <= 4'h0cb6;
         4'hd253 	:	val_out <= 4'h0cb6;
         4'hd258 	:	val_out <= 4'h0cc1;
         4'hd259 	:	val_out <= 4'h0cc1;
         4'hd25a 	:	val_out <= 4'h0cc1;
         4'hd25b 	:	val_out <= 4'h0cc1;
         4'hd260 	:	val_out <= 4'h0ccc;
         4'hd261 	:	val_out <= 4'h0ccc;
         4'hd262 	:	val_out <= 4'h0ccc;
         4'hd263 	:	val_out <= 4'h0ccc;
         4'hd268 	:	val_out <= 4'h0cd7;
         4'hd269 	:	val_out <= 4'h0cd7;
         4'hd26a 	:	val_out <= 4'h0cd7;
         4'hd26b 	:	val_out <= 4'h0cd7;
         4'hd270 	:	val_out <= 4'h0ce2;
         4'hd271 	:	val_out <= 4'h0ce2;
         4'hd272 	:	val_out <= 4'h0ce2;
         4'hd273 	:	val_out <= 4'h0ce2;
         4'hd278 	:	val_out <= 4'h0ced;
         4'hd279 	:	val_out <= 4'h0ced;
         4'hd27a 	:	val_out <= 4'h0ced;
         4'hd27b 	:	val_out <= 4'h0ced;
         4'hd280 	:	val_out <= 4'h0cf8;
         4'hd281 	:	val_out <= 4'h0cf8;
         4'hd282 	:	val_out <= 4'h0cf8;
         4'hd283 	:	val_out <= 4'h0cf8;
         4'hd288 	:	val_out <= 4'h0d03;
         4'hd289 	:	val_out <= 4'h0d03;
         4'hd28a 	:	val_out <= 4'h0d03;
         4'hd28b 	:	val_out <= 4'h0d03;
         4'hd290 	:	val_out <= 4'h0d0e;
         4'hd291 	:	val_out <= 4'h0d0e;
         4'hd292 	:	val_out <= 4'h0d0e;
         4'hd293 	:	val_out <= 4'h0d0e;
         4'hd298 	:	val_out <= 4'h0d19;
         4'hd299 	:	val_out <= 4'h0d19;
         4'hd29a 	:	val_out <= 4'h0d19;
         4'hd29b 	:	val_out <= 4'h0d19;
         4'hd2a0 	:	val_out <= 4'h0d24;
         4'hd2a1 	:	val_out <= 4'h0d24;
         4'hd2a2 	:	val_out <= 4'h0d24;
         4'hd2a3 	:	val_out <= 4'h0d24;
         4'hd2a8 	:	val_out <= 4'h0d2f;
         4'hd2a9 	:	val_out <= 4'h0d2f;
         4'hd2aa 	:	val_out <= 4'h0d2f;
         4'hd2ab 	:	val_out <= 4'h0d2f;
         4'hd2b0 	:	val_out <= 4'h0d3a;
         4'hd2b1 	:	val_out <= 4'h0d3a;
         4'hd2b2 	:	val_out <= 4'h0d3a;
         4'hd2b3 	:	val_out <= 4'h0d3a;
         4'hd2b8 	:	val_out <= 4'h0d45;
         4'hd2b9 	:	val_out <= 4'h0d45;
         4'hd2ba 	:	val_out <= 4'h0d45;
         4'hd2bb 	:	val_out <= 4'h0d45;
         4'hd2c0 	:	val_out <= 4'h0d50;
         4'hd2c1 	:	val_out <= 4'h0d50;
         4'hd2c2 	:	val_out <= 4'h0d50;
         4'hd2c3 	:	val_out <= 4'h0d50;
         4'hd2c8 	:	val_out <= 4'h0d5c;
         4'hd2c9 	:	val_out <= 4'h0d5c;
         4'hd2ca 	:	val_out <= 4'h0d5c;
         4'hd2cb 	:	val_out <= 4'h0d5c;
         4'hd2d0 	:	val_out <= 4'h0d67;
         4'hd2d1 	:	val_out <= 4'h0d67;
         4'hd2d2 	:	val_out <= 4'h0d67;
         4'hd2d3 	:	val_out <= 4'h0d67;
         4'hd2d8 	:	val_out <= 4'h0d72;
         4'hd2d9 	:	val_out <= 4'h0d72;
         4'hd2da 	:	val_out <= 4'h0d72;
         4'hd2db 	:	val_out <= 4'h0d72;
         4'hd2e0 	:	val_out <= 4'h0d7d;
         4'hd2e1 	:	val_out <= 4'h0d7d;
         4'hd2e2 	:	val_out <= 4'h0d7d;
         4'hd2e3 	:	val_out <= 4'h0d7d;
         4'hd2e8 	:	val_out <= 4'h0d89;
         4'hd2e9 	:	val_out <= 4'h0d89;
         4'hd2ea 	:	val_out <= 4'h0d89;
         4'hd2eb 	:	val_out <= 4'h0d89;
         4'hd2f0 	:	val_out <= 4'h0d94;
         4'hd2f1 	:	val_out <= 4'h0d94;
         4'hd2f2 	:	val_out <= 4'h0d94;
         4'hd2f3 	:	val_out <= 4'h0d94;
         4'hd2f8 	:	val_out <= 4'h0d9f;
         4'hd2f9 	:	val_out <= 4'h0d9f;
         4'hd2fa 	:	val_out <= 4'h0d9f;
         4'hd2fb 	:	val_out <= 4'h0d9f;
         4'hd300 	:	val_out <= 4'h0daa;
         4'hd301 	:	val_out <= 4'h0daa;
         4'hd302 	:	val_out <= 4'h0daa;
         4'hd303 	:	val_out <= 4'h0daa;
         4'hd308 	:	val_out <= 4'h0db6;
         4'hd309 	:	val_out <= 4'h0db6;
         4'hd30a 	:	val_out <= 4'h0db6;
         4'hd30b 	:	val_out <= 4'h0db6;
         4'hd310 	:	val_out <= 4'h0dc1;
         4'hd311 	:	val_out <= 4'h0dc1;
         4'hd312 	:	val_out <= 4'h0dc1;
         4'hd313 	:	val_out <= 4'h0dc1;
         4'hd318 	:	val_out <= 4'h0dcc;
         4'hd319 	:	val_out <= 4'h0dcc;
         4'hd31a 	:	val_out <= 4'h0dcc;
         4'hd31b 	:	val_out <= 4'h0dcc;
         4'hd320 	:	val_out <= 4'h0dd8;
         4'hd321 	:	val_out <= 4'h0dd8;
         4'hd322 	:	val_out <= 4'h0dd8;
         4'hd323 	:	val_out <= 4'h0dd8;
         4'hd328 	:	val_out <= 4'h0de3;
         4'hd329 	:	val_out <= 4'h0de3;
         4'hd32a 	:	val_out <= 4'h0de3;
         4'hd32b 	:	val_out <= 4'h0de3;
         4'hd330 	:	val_out <= 4'h0dee;
         4'hd331 	:	val_out <= 4'h0dee;
         4'hd332 	:	val_out <= 4'h0dee;
         4'hd333 	:	val_out <= 4'h0dee;
         4'hd338 	:	val_out <= 4'h0dfa;
         4'hd339 	:	val_out <= 4'h0dfa;
         4'hd33a 	:	val_out <= 4'h0dfa;
         4'hd33b 	:	val_out <= 4'h0dfa;
         4'hd340 	:	val_out <= 4'h0e05;
         4'hd341 	:	val_out <= 4'h0e05;
         4'hd342 	:	val_out <= 4'h0e05;
         4'hd343 	:	val_out <= 4'h0e05;
         4'hd348 	:	val_out <= 4'h0e11;
         4'hd349 	:	val_out <= 4'h0e11;
         4'hd34a 	:	val_out <= 4'h0e11;
         4'hd34b 	:	val_out <= 4'h0e11;
         4'hd350 	:	val_out <= 4'h0e1c;
         4'hd351 	:	val_out <= 4'h0e1c;
         4'hd352 	:	val_out <= 4'h0e1c;
         4'hd353 	:	val_out <= 4'h0e1c;
         4'hd358 	:	val_out <= 4'h0e28;
         4'hd359 	:	val_out <= 4'h0e28;
         4'hd35a 	:	val_out <= 4'h0e28;
         4'hd35b 	:	val_out <= 4'h0e28;
         4'hd360 	:	val_out <= 4'h0e33;
         4'hd361 	:	val_out <= 4'h0e33;
         4'hd362 	:	val_out <= 4'h0e33;
         4'hd363 	:	val_out <= 4'h0e33;
         4'hd368 	:	val_out <= 4'h0e3f;
         4'hd369 	:	val_out <= 4'h0e3f;
         4'hd36a 	:	val_out <= 4'h0e3f;
         4'hd36b 	:	val_out <= 4'h0e3f;
         4'hd370 	:	val_out <= 4'h0e4a;
         4'hd371 	:	val_out <= 4'h0e4a;
         4'hd372 	:	val_out <= 4'h0e4a;
         4'hd373 	:	val_out <= 4'h0e4a;
         4'hd378 	:	val_out <= 4'h0e56;
         4'hd379 	:	val_out <= 4'h0e56;
         4'hd37a 	:	val_out <= 4'h0e56;
         4'hd37b 	:	val_out <= 4'h0e56;
         4'hd380 	:	val_out <= 4'h0e61;
         4'hd381 	:	val_out <= 4'h0e61;
         4'hd382 	:	val_out <= 4'h0e61;
         4'hd383 	:	val_out <= 4'h0e61;
         4'hd388 	:	val_out <= 4'h0e6d;
         4'hd389 	:	val_out <= 4'h0e6d;
         4'hd38a 	:	val_out <= 4'h0e6d;
         4'hd38b 	:	val_out <= 4'h0e6d;
         4'hd390 	:	val_out <= 4'h0e79;
         4'hd391 	:	val_out <= 4'h0e79;
         4'hd392 	:	val_out <= 4'h0e79;
         4'hd393 	:	val_out <= 4'h0e79;
         4'hd398 	:	val_out <= 4'h0e84;
         4'hd399 	:	val_out <= 4'h0e84;
         4'hd39a 	:	val_out <= 4'h0e84;
         4'hd39b 	:	val_out <= 4'h0e84;
         4'hd3a0 	:	val_out <= 4'h0e90;
         4'hd3a1 	:	val_out <= 4'h0e90;
         4'hd3a2 	:	val_out <= 4'h0e90;
         4'hd3a3 	:	val_out <= 4'h0e90;
         4'hd3a8 	:	val_out <= 4'h0e9b;
         4'hd3a9 	:	val_out <= 4'h0e9b;
         4'hd3aa 	:	val_out <= 4'h0e9b;
         4'hd3ab 	:	val_out <= 4'h0e9b;
         4'hd3b0 	:	val_out <= 4'h0ea7;
         4'hd3b1 	:	val_out <= 4'h0ea7;
         4'hd3b2 	:	val_out <= 4'h0ea7;
         4'hd3b3 	:	val_out <= 4'h0ea7;
         4'hd3b8 	:	val_out <= 4'h0eb3;
         4'hd3b9 	:	val_out <= 4'h0eb3;
         4'hd3ba 	:	val_out <= 4'h0eb3;
         4'hd3bb 	:	val_out <= 4'h0eb3;
         4'hd3c0 	:	val_out <= 4'h0ebe;
         4'hd3c1 	:	val_out <= 4'h0ebe;
         4'hd3c2 	:	val_out <= 4'h0ebe;
         4'hd3c3 	:	val_out <= 4'h0ebe;
         4'hd3c8 	:	val_out <= 4'h0eca;
         4'hd3c9 	:	val_out <= 4'h0eca;
         4'hd3ca 	:	val_out <= 4'h0eca;
         4'hd3cb 	:	val_out <= 4'h0eca;
         4'hd3d0 	:	val_out <= 4'h0ed6;
         4'hd3d1 	:	val_out <= 4'h0ed6;
         4'hd3d2 	:	val_out <= 4'h0ed6;
         4'hd3d3 	:	val_out <= 4'h0ed6;
         4'hd3d8 	:	val_out <= 4'h0ee2;
         4'hd3d9 	:	val_out <= 4'h0ee2;
         4'hd3da 	:	val_out <= 4'h0ee2;
         4'hd3db 	:	val_out <= 4'h0ee2;
         4'hd3e0 	:	val_out <= 4'h0eed;
         4'hd3e1 	:	val_out <= 4'h0eed;
         4'hd3e2 	:	val_out <= 4'h0eed;
         4'hd3e3 	:	val_out <= 4'h0eed;
         4'hd3e8 	:	val_out <= 4'h0ef9;
         4'hd3e9 	:	val_out <= 4'h0ef9;
         4'hd3ea 	:	val_out <= 4'h0ef9;
         4'hd3eb 	:	val_out <= 4'h0ef9;
         4'hd3f0 	:	val_out <= 4'h0f05;
         4'hd3f1 	:	val_out <= 4'h0f05;
         4'hd3f2 	:	val_out <= 4'h0f05;
         4'hd3f3 	:	val_out <= 4'h0f05;
         4'hd3f8 	:	val_out <= 4'h0f11;
         4'hd3f9 	:	val_out <= 4'h0f11;
         4'hd3fa 	:	val_out <= 4'h0f11;
         4'hd3fb 	:	val_out <= 4'h0f11;
         4'hd400 	:	val_out <= 4'h0f1d;
         4'hd401 	:	val_out <= 4'h0f1d;
         4'hd402 	:	val_out <= 4'h0f1d;
         4'hd403 	:	val_out <= 4'h0f1d;
         4'hd408 	:	val_out <= 4'h0f29;
         4'hd409 	:	val_out <= 4'h0f29;
         4'hd40a 	:	val_out <= 4'h0f29;
         4'hd40b 	:	val_out <= 4'h0f29;
         4'hd410 	:	val_out <= 4'h0f34;
         4'hd411 	:	val_out <= 4'h0f34;
         4'hd412 	:	val_out <= 4'h0f34;
         4'hd413 	:	val_out <= 4'h0f34;
         4'hd418 	:	val_out <= 4'h0f40;
         4'hd419 	:	val_out <= 4'h0f40;
         4'hd41a 	:	val_out <= 4'h0f40;
         4'hd41b 	:	val_out <= 4'h0f40;
         4'hd420 	:	val_out <= 4'h0f4c;
         4'hd421 	:	val_out <= 4'h0f4c;
         4'hd422 	:	val_out <= 4'h0f4c;
         4'hd423 	:	val_out <= 4'h0f4c;
         4'hd428 	:	val_out <= 4'h0f58;
         4'hd429 	:	val_out <= 4'h0f58;
         4'hd42a 	:	val_out <= 4'h0f58;
         4'hd42b 	:	val_out <= 4'h0f58;
         4'hd430 	:	val_out <= 4'h0f64;
         4'hd431 	:	val_out <= 4'h0f64;
         4'hd432 	:	val_out <= 4'h0f64;
         4'hd433 	:	val_out <= 4'h0f64;
         4'hd438 	:	val_out <= 4'h0f70;
         4'hd439 	:	val_out <= 4'h0f70;
         4'hd43a 	:	val_out <= 4'h0f70;
         4'hd43b 	:	val_out <= 4'h0f70;
         4'hd440 	:	val_out <= 4'h0f7c;
         4'hd441 	:	val_out <= 4'h0f7c;
         4'hd442 	:	val_out <= 4'h0f7c;
         4'hd443 	:	val_out <= 4'h0f7c;
         4'hd448 	:	val_out <= 4'h0f88;
         4'hd449 	:	val_out <= 4'h0f88;
         4'hd44a 	:	val_out <= 4'h0f88;
         4'hd44b 	:	val_out <= 4'h0f88;
         4'hd450 	:	val_out <= 4'h0f94;
         4'hd451 	:	val_out <= 4'h0f94;
         4'hd452 	:	val_out <= 4'h0f94;
         4'hd453 	:	val_out <= 4'h0f94;
         4'hd458 	:	val_out <= 4'h0fa0;
         4'hd459 	:	val_out <= 4'h0fa0;
         4'hd45a 	:	val_out <= 4'h0fa0;
         4'hd45b 	:	val_out <= 4'h0fa0;
         4'hd460 	:	val_out <= 4'h0fac;
         4'hd461 	:	val_out <= 4'h0fac;
         4'hd462 	:	val_out <= 4'h0fac;
         4'hd463 	:	val_out <= 4'h0fac;
         4'hd468 	:	val_out <= 4'h0fb8;
         4'hd469 	:	val_out <= 4'h0fb8;
         4'hd46a 	:	val_out <= 4'h0fb8;
         4'hd46b 	:	val_out <= 4'h0fb8;
         4'hd470 	:	val_out <= 4'h0fc4;
         4'hd471 	:	val_out <= 4'h0fc4;
         4'hd472 	:	val_out <= 4'h0fc4;
         4'hd473 	:	val_out <= 4'h0fc4;
         4'hd478 	:	val_out <= 4'h0fd0;
         4'hd479 	:	val_out <= 4'h0fd0;
         4'hd47a 	:	val_out <= 4'h0fd0;
         4'hd47b 	:	val_out <= 4'h0fd0;
         4'hd480 	:	val_out <= 4'h0fdc;
         4'hd481 	:	val_out <= 4'h0fdc;
         4'hd482 	:	val_out <= 4'h0fdc;
         4'hd483 	:	val_out <= 4'h0fdc;
         4'hd488 	:	val_out <= 4'h0fe9;
         4'hd489 	:	val_out <= 4'h0fe9;
         4'hd48a 	:	val_out <= 4'h0fe9;
         4'hd48b 	:	val_out <= 4'h0fe9;
         4'hd490 	:	val_out <= 4'h0ff5;
         4'hd491 	:	val_out <= 4'h0ff5;
         4'hd492 	:	val_out <= 4'h0ff5;
         4'hd493 	:	val_out <= 4'h0ff5;
         4'hd498 	:	val_out <= 4'h1001;
         4'hd499 	:	val_out <= 4'h1001;
         4'hd49a 	:	val_out <= 4'h1001;
         4'hd49b 	:	val_out <= 4'h1001;
         4'hd4a0 	:	val_out <= 4'h100d;
         4'hd4a1 	:	val_out <= 4'h100d;
         4'hd4a2 	:	val_out <= 4'h100d;
         4'hd4a3 	:	val_out <= 4'h100d;
         4'hd4a8 	:	val_out <= 4'h1019;
         4'hd4a9 	:	val_out <= 4'h1019;
         4'hd4aa 	:	val_out <= 4'h1019;
         4'hd4ab 	:	val_out <= 4'h1019;
         4'hd4b0 	:	val_out <= 4'h1025;
         4'hd4b1 	:	val_out <= 4'h1025;
         4'hd4b2 	:	val_out <= 4'h1025;
         4'hd4b3 	:	val_out <= 4'h1025;
         4'hd4b8 	:	val_out <= 4'h1032;
         4'hd4b9 	:	val_out <= 4'h1032;
         4'hd4ba 	:	val_out <= 4'h1032;
         4'hd4bb 	:	val_out <= 4'h1032;
         4'hd4c0 	:	val_out <= 4'h103e;
         4'hd4c1 	:	val_out <= 4'h103e;
         4'hd4c2 	:	val_out <= 4'h103e;
         4'hd4c3 	:	val_out <= 4'h103e;
         4'hd4c8 	:	val_out <= 4'h104a;
         4'hd4c9 	:	val_out <= 4'h104a;
         4'hd4ca 	:	val_out <= 4'h104a;
         4'hd4cb 	:	val_out <= 4'h104a;
         4'hd4d0 	:	val_out <= 4'h1056;
         4'hd4d1 	:	val_out <= 4'h1056;
         4'hd4d2 	:	val_out <= 4'h1056;
         4'hd4d3 	:	val_out <= 4'h1056;
         4'hd4d8 	:	val_out <= 4'h1063;
         4'hd4d9 	:	val_out <= 4'h1063;
         4'hd4da 	:	val_out <= 4'h1063;
         4'hd4db 	:	val_out <= 4'h1063;
         4'hd4e0 	:	val_out <= 4'h106f;
         4'hd4e1 	:	val_out <= 4'h106f;
         4'hd4e2 	:	val_out <= 4'h106f;
         4'hd4e3 	:	val_out <= 4'h106f;
         4'hd4e8 	:	val_out <= 4'h107b;
         4'hd4e9 	:	val_out <= 4'h107b;
         4'hd4ea 	:	val_out <= 4'h107b;
         4'hd4eb 	:	val_out <= 4'h107b;
         4'hd4f0 	:	val_out <= 4'h1088;
         4'hd4f1 	:	val_out <= 4'h1088;
         4'hd4f2 	:	val_out <= 4'h1088;
         4'hd4f3 	:	val_out <= 4'h1088;
         4'hd4f8 	:	val_out <= 4'h1094;
         4'hd4f9 	:	val_out <= 4'h1094;
         4'hd4fa 	:	val_out <= 4'h1094;
         4'hd4fb 	:	val_out <= 4'h1094;
         4'hd500 	:	val_out <= 4'h10a0;
         4'hd501 	:	val_out <= 4'h10a0;
         4'hd502 	:	val_out <= 4'h10a0;
         4'hd503 	:	val_out <= 4'h10a0;
         4'hd508 	:	val_out <= 4'h10ad;
         4'hd509 	:	val_out <= 4'h10ad;
         4'hd50a 	:	val_out <= 4'h10ad;
         4'hd50b 	:	val_out <= 4'h10ad;
         4'hd510 	:	val_out <= 4'h10b9;
         4'hd511 	:	val_out <= 4'h10b9;
         4'hd512 	:	val_out <= 4'h10b9;
         4'hd513 	:	val_out <= 4'h10b9;
         4'hd518 	:	val_out <= 4'h10c6;
         4'hd519 	:	val_out <= 4'h10c6;
         4'hd51a 	:	val_out <= 4'h10c6;
         4'hd51b 	:	val_out <= 4'h10c6;
         4'hd520 	:	val_out <= 4'h10d2;
         4'hd521 	:	val_out <= 4'h10d2;
         4'hd522 	:	val_out <= 4'h10d2;
         4'hd523 	:	val_out <= 4'h10d2;
         4'hd528 	:	val_out <= 4'h10df;
         4'hd529 	:	val_out <= 4'h10df;
         4'hd52a 	:	val_out <= 4'h10df;
         4'hd52b 	:	val_out <= 4'h10df;
         4'hd530 	:	val_out <= 4'h10eb;
         4'hd531 	:	val_out <= 4'h10eb;
         4'hd532 	:	val_out <= 4'h10eb;
         4'hd533 	:	val_out <= 4'h10eb;
         4'hd538 	:	val_out <= 4'h10f8;
         4'hd539 	:	val_out <= 4'h10f8;
         4'hd53a 	:	val_out <= 4'h10f8;
         4'hd53b 	:	val_out <= 4'h10f8;
         4'hd540 	:	val_out <= 4'h1104;
         4'hd541 	:	val_out <= 4'h1104;
         4'hd542 	:	val_out <= 4'h1104;
         4'hd543 	:	val_out <= 4'h1104;
         4'hd548 	:	val_out <= 4'h1111;
         4'hd549 	:	val_out <= 4'h1111;
         4'hd54a 	:	val_out <= 4'h1111;
         4'hd54b 	:	val_out <= 4'h1111;
         4'hd550 	:	val_out <= 4'h111d;
         4'hd551 	:	val_out <= 4'h111d;
         4'hd552 	:	val_out <= 4'h111d;
         4'hd553 	:	val_out <= 4'h111d;
         4'hd558 	:	val_out <= 4'h112a;
         4'hd559 	:	val_out <= 4'h112a;
         4'hd55a 	:	val_out <= 4'h112a;
         4'hd55b 	:	val_out <= 4'h112a;
         4'hd560 	:	val_out <= 4'h1136;
         4'hd561 	:	val_out <= 4'h1136;
         4'hd562 	:	val_out <= 4'h1136;
         4'hd563 	:	val_out <= 4'h1136;
         4'hd568 	:	val_out <= 4'h1143;
         4'hd569 	:	val_out <= 4'h1143;
         4'hd56a 	:	val_out <= 4'h1143;
         4'hd56b 	:	val_out <= 4'h1143;
         4'hd570 	:	val_out <= 4'h1150;
         4'hd571 	:	val_out <= 4'h1150;
         4'hd572 	:	val_out <= 4'h1150;
         4'hd573 	:	val_out <= 4'h1150;
         4'hd578 	:	val_out <= 4'h115c;
         4'hd579 	:	val_out <= 4'h115c;
         4'hd57a 	:	val_out <= 4'h115c;
         4'hd57b 	:	val_out <= 4'h115c;
         4'hd580 	:	val_out <= 4'h1169;
         4'hd581 	:	val_out <= 4'h1169;
         4'hd582 	:	val_out <= 4'h1169;
         4'hd583 	:	val_out <= 4'h1169;
         4'hd588 	:	val_out <= 4'h1176;
         4'hd589 	:	val_out <= 4'h1176;
         4'hd58a 	:	val_out <= 4'h1176;
         4'hd58b 	:	val_out <= 4'h1176;
         4'hd590 	:	val_out <= 4'h1182;
         4'hd591 	:	val_out <= 4'h1182;
         4'hd592 	:	val_out <= 4'h1182;
         4'hd593 	:	val_out <= 4'h1182;
         4'hd598 	:	val_out <= 4'h118f;
         4'hd599 	:	val_out <= 4'h118f;
         4'hd59a 	:	val_out <= 4'h118f;
         4'hd59b 	:	val_out <= 4'h118f;
         4'hd5a0 	:	val_out <= 4'h119c;
         4'hd5a1 	:	val_out <= 4'h119c;
         4'hd5a2 	:	val_out <= 4'h119c;
         4'hd5a3 	:	val_out <= 4'h119c;
         4'hd5a8 	:	val_out <= 4'h11a8;
         4'hd5a9 	:	val_out <= 4'h11a8;
         4'hd5aa 	:	val_out <= 4'h11a8;
         4'hd5ab 	:	val_out <= 4'h11a8;
         4'hd5b0 	:	val_out <= 4'h11b5;
         4'hd5b1 	:	val_out <= 4'h11b5;
         4'hd5b2 	:	val_out <= 4'h11b5;
         4'hd5b3 	:	val_out <= 4'h11b5;
         4'hd5b8 	:	val_out <= 4'h11c2;
         4'hd5b9 	:	val_out <= 4'h11c2;
         4'hd5ba 	:	val_out <= 4'h11c2;
         4'hd5bb 	:	val_out <= 4'h11c2;
         4'hd5c0 	:	val_out <= 4'h11cf;
         4'hd5c1 	:	val_out <= 4'h11cf;
         4'hd5c2 	:	val_out <= 4'h11cf;
         4'hd5c3 	:	val_out <= 4'h11cf;
         4'hd5c8 	:	val_out <= 4'h11db;
         4'hd5c9 	:	val_out <= 4'h11db;
         4'hd5ca 	:	val_out <= 4'h11db;
         4'hd5cb 	:	val_out <= 4'h11db;
         4'hd5d0 	:	val_out <= 4'h11e8;
         4'hd5d1 	:	val_out <= 4'h11e8;
         4'hd5d2 	:	val_out <= 4'h11e8;
         4'hd5d3 	:	val_out <= 4'h11e8;
         4'hd5d8 	:	val_out <= 4'h11f5;
         4'hd5d9 	:	val_out <= 4'h11f5;
         4'hd5da 	:	val_out <= 4'h11f5;
         4'hd5db 	:	val_out <= 4'h11f5;
         4'hd5e0 	:	val_out <= 4'h1202;
         4'hd5e1 	:	val_out <= 4'h1202;
         4'hd5e2 	:	val_out <= 4'h1202;
         4'hd5e3 	:	val_out <= 4'h1202;
         4'hd5e8 	:	val_out <= 4'h120f;
         4'hd5e9 	:	val_out <= 4'h120f;
         4'hd5ea 	:	val_out <= 4'h120f;
         4'hd5eb 	:	val_out <= 4'h120f;
         4'hd5f0 	:	val_out <= 4'h121c;
         4'hd5f1 	:	val_out <= 4'h121c;
         4'hd5f2 	:	val_out <= 4'h121c;
         4'hd5f3 	:	val_out <= 4'h121c;
         4'hd5f8 	:	val_out <= 4'h1229;
         4'hd5f9 	:	val_out <= 4'h1229;
         4'hd5fa 	:	val_out <= 4'h1229;
         4'hd5fb 	:	val_out <= 4'h1229;
         4'hd600 	:	val_out <= 4'h1235;
         4'hd601 	:	val_out <= 4'h1235;
         4'hd602 	:	val_out <= 4'h1235;
         4'hd603 	:	val_out <= 4'h1235;
         4'hd608 	:	val_out <= 4'h1242;
         4'hd609 	:	val_out <= 4'h1242;
         4'hd60a 	:	val_out <= 4'h1242;
         4'hd60b 	:	val_out <= 4'h1242;
         4'hd610 	:	val_out <= 4'h124f;
         4'hd611 	:	val_out <= 4'h124f;
         4'hd612 	:	val_out <= 4'h124f;
         4'hd613 	:	val_out <= 4'h124f;
         4'hd618 	:	val_out <= 4'h125c;
         4'hd619 	:	val_out <= 4'h125c;
         4'hd61a 	:	val_out <= 4'h125c;
         4'hd61b 	:	val_out <= 4'h125c;
         4'hd620 	:	val_out <= 4'h1269;
         4'hd621 	:	val_out <= 4'h1269;
         4'hd622 	:	val_out <= 4'h1269;
         4'hd623 	:	val_out <= 4'h1269;
         4'hd628 	:	val_out <= 4'h1276;
         4'hd629 	:	val_out <= 4'h1276;
         4'hd62a 	:	val_out <= 4'h1276;
         4'hd62b 	:	val_out <= 4'h1276;
         4'hd630 	:	val_out <= 4'h1283;
         4'hd631 	:	val_out <= 4'h1283;
         4'hd632 	:	val_out <= 4'h1283;
         4'hd633 	:	val_out <= 4'h1283;
         4'hd638 	:	val_out <= 4'h1290;
         4'hd639 	:	val_out <= 4'h1290;
         4'hd63a 	:	val_out <= 4'h1290;
         4'hd63b 	:	val_out <= 4'h1290;
         4'hd640 	:	val_out <= 4'h129d;
         4'hd641 	:	val_out <= 4'h129d;
         4'hd642 	:	val_out <= 4'h129d;
         4'hd643 	:	val_out <= 4'h129d;
         4'hd648 	:	val_out <= 4'h12aa;
         4'hd649 	:	val_out <= 4'h12aa;
         4'hd64a 	:	val_out <= 4'h12aa;
         4'hd64b 	:	val_out <= 4'h12aa;
         4'hd650 	:	val_out <= 4'h12b7;
         4'hd651 	:	val_out <= 4'h12b7;
         4'hd652 	:	val_out <= 4'h12b7;
         4'hd653 	:	val_out <= 4'h12b7;
         4'hd658 	:	val_out <= 4'h12c5;
         4'hd659 	:	val_out <= 4'h12c5;
         4'hd65a 	:	val_out <= 4'h12c5;
         4'hd65b 	:	val_out <= 4'h12c5;
         4'hd660 	:	val_out <= 4'h12d2;
         4'hd661 	:	val_out <= 4'h12d2;
         4'hd662 	:	val_out <= 4'h12d2;
         4'hd663 	:	val_out <= 4'h12d2;
         4'hd668 	:	val_out <= 4'h12df;
         4'hd669 	:	val_out <= 4'h12df;
         4'hd66a 	:	val_out <= 4'h12df;
         4'hd66b 	:	val_out <= 4'h12df;
         4'hd670 	:	val_out <= 4'h12ec;
         4'hd671 	:	val_out <= 4'h12ec;
         4'hd672 	:	val_out <= 4'h12ec;
         4'hd673 	:	val_out <= 4'h12ec;
         4'hd678 	:	val_out <= 4'h12f9;
         4'hd679 	:	val_out <= 4'h12f9;
         4'hd67a 	:	val_out <= 4'h12f9;
         4'hd67b 	:	val_out <= 4'h12f9;
         4'hd680 	:	val_out <= 4'h1306;
         4'hd681 	:	val_out <= 4'h1306;
         4'hd682 	:	val_out <= 4'h1306;
         4'hd683 	:	val_out <= 4'h1306;
         4'hd688 	:	val_out <= 4'h1313;
         4'hd689 	:	val_out <= 4'h1313;
         4'hd68a 	:	val_out <= 4'h1313;
         4'hd68b 	:	val_out <= 4'h1313;
         4'hd690 	:	val_out <= 4'h1321;
         4'hd691 	:	val_out <= 4'h1321;
         4'hd692 	:	val_out <= 4'h1321;
         4'hd693 	:	val_out <= 4'h1321;
         4'hd698 	:	val_out <= 4'h132e;
         4'hd699 	:	val_out <= 4'h132e;
         4'hd69a 	:	val_out <= 4'h132e;
         4'hd69b 	:	val_out <= 4'h132e;
         4'hd6a0 	:	val_out <= 4'h133b;
         4'hd6a1 	:	val_out <= 4'h133b;
         4'hd6a2 	:	val_out <= 4'h133b;
         4'hd6a3 	:	val_out <= 4'h133b;
         4'hd6a8 	:	val_out <= 4'h1348;
         4'hd6a9 	:	val_out <= 4'h1348;
         4'hd6aa 	:	val_out <= 4'h1348;
         4'hd6ab 	:	val_out <= 4'h1348;
         4'hd6b0 	:	val_out <= 4'h1356;
         4'hd6b1 	:	val_out <= 4'h1356;
         4'hd6b2 	:	val_out <= 4'h1356;
         4'hd6b3 	:	val_out <= 4'h1356;
         4'hd6b8 	:	val_out <= 4'h1363;
         4'hd6b9 	:	val_out <= 4'h1363;
         4'hd6ba 	:	val_out <= 4'h1363;
         4'hd6bb 	:	val_out <= 4'h1363;
         4'hd6c0 	:	val_out <= 4'h1370;
         4'hd6c1 	:	val_out <= 4'h1370;
         4'hd6c2 	:	val_out <= 4'h1370;
         4'hd6c3 	:	val_out <= 4'h1370;
         4'hd6c8 	:	val_out <= 4'h137e;
         4'hd6c9 	:	val_out <= 4'h137e;
         4'hd6ca 	:	val_out <= 4'h137e;
         4'hd6cb 	:	val_out <= 4'h137e;
         4'hd6d0 	:	val_out <= 4'h138b;
         4'hd6d1 	:	val_out <= 4'h138b;
         4'hd6d2 	:	val_out <= 4'h138b;
         4'hd6d3 	:	val_out <= 4'h138b;
         4'hd6d8 	:	val_out <= 4'h1398;
         4'hd6d9 	:	val_out <= 4'h1398;
         4'hd6da 	:	val_out <= 4'h1398;
         4'hd6db 	:	val_out <= 4'h1398;
         4'hd6e0 	:	val_out <= 4'h13a6;
         4'hd6e1 	:	val_out <= 4'h13a6;
         4'hd6e2 	:	val_out <= 4'h13a6;
         4'hd6e3 	:	val_out <= 4'h13a6;
         4'hd6e8 	:	val_out <= 4'h13b3;
         4'hd6e9 	:	val_out <= 4'h13b3;
         4'hd6ea 	:	val_out <= 4'h13b3;
         4'hd6eb 	:	val_out <= 4'h13b3;
         4'hd6f0 	:	val_out <= 4'h13c0;
         4'hd6f1 	:	val_out <= 4'h13c0;
         4'hd6f2 	:	val_out <= 4'h13c0;
         4'hd6f3 	:	val_out <= 4'h13c0;
         4'hd6f8 	:	val_out <= 4'h13ce;
         4'hd6f9 	:	val_out <= 4'h13ce;
         4'hd6fa 	:	val_out <= 4'h13ce;
         4'hd6fb 	:	val_out <= 4'h13ce;
         4'hd700 	:	val_out <= 4'h13db;
         4'hd701 	:	val_out <= 4'h13db;
         4'hd702 	:	val_out <= 4'h13db;
         4'hd703 	:	val_out <= 4'h13db;
         4'hd708 	:	val_out <= 4'h13e9;
         4'hd709 	:	val_out <= 4'h13e9;
         4'hd70a 	:	val_out <= 4'h13e9;
         4'hd70b 	:	val_out <= 4'h13e9;
         4'hd710 	:	val_out <= 4'h13f6;
         4'hd711 	:	val_out <= 4'h13f6;
         4'hd712 	:	val_out <= 4'h13f6;
         4'hd713 	:	val_out <= 4'h13f6;
         4'hd718 	:	val_out <= 4'h1404;
         4'hd719 	:	val_out <= 4'h1404;
         4'hd71a 	:	val_out <= 4'h1404;
         4'hd71b 	:	val_out <= 4'h1404;
         4'hd720 	:	val_out <= 4'h1411;
         4'hd721 	:	val_out <= 4'h1411;
         4'hd722 	:	val_out <= 4'h1411;
         4'hd723 	:	val_out <= 4'h1411;
         4'hd728 	:	val_out <= 4'h141f;
         4'hd729 	:	val_out <= 4'h141f;
         4'hd72a 	:	val_out <= 4'h141f;
         4'hd72b 	:	val_out <= 4'h141f;
         4'hd730 	:	val_out <= 4'h142c;
         4'hd731 	:	val_out <= 4'h142c;
         4'hd732 	:	val_out <= 4'h142c;
         4'hd733 	:	val_out <= 4'h142c;
         4'hd738 	:	val_out <= 4'h143a;
         4'hd739 	:	val_out <= 4'h143a;
         4'hd73a 	:	val_out <= 4'h143a;
         4'hd73b 	:	val_out <= 4'h143a;
         4'hd740 	:	val_out <= 4'h1447;
         4'hd741 	:	val_out <= 4'h1447;
         4'hd742 	:	val_out <= 4'h1447;
         4'hd743 	:	val_out <= 4'h1447;
         4'hd748 	:	val_out <= 4'h1455;
         4'hd749 	:	val_out <= 4'h1455;
         4'hd74a 	:	val_out <= 4'h1455;
         4'hd74b 	:	val_out <= 4'h1455;
         4'hd750 	:	val_out <= 4'h1463;
         4'hd751 	:	val_out <= 4'h1463;
         4'hd752 	:	val_out <= 4'h1463;
         4'hd753 	:	val_out <= 4'h1463;
         4'hd758 	:	val_out <= 4'h1470;
         4'hd759 	:	val_out <= 4'h1470;
         4'hd75a 	:	val_out <= 4'h1470;
         4'hd75b 	:	val_out <= 4'h1470;
         4'hd760 	:	val_out <= 4'h147e;
         4'hd761 	:	val_out <= 4'h147e;
         4'hd762 	:	val_out <= 4'h147e;
         4'hd763 	:	val_out <= 4'h147e;
         4'hd768 	:	val_out <= 4'h148c;
         4'hd769 	:	val_out <= 4'h148c;
         4'hd76a 	:	val_out <= 4'h148c;
         4'hd76b 	:	val_out <= 4'h148c;
         4'hd770 	:	val_out <= 4'h1499;
         4'hd771 	:	val_out <= 4'h1499;
         4'hd772 	:	val_out <= 4'h1499;
         4'hd773 	:	val_out <= 4'h1499;
         4'hd778 	:	val_out <= 4'h14a7;
         4'hd779 	:	val_out <= 4'h14a7;
         4'hd77a 	:	val_out <= 4'h14a7;
         4'hd77b 	:	val_out <= 4'h14a7;
         4'hd780 	:	val_out <= 4'h14b5;
         4'hd781 	:	val_out <= 4'h14b5;
         4'hd782 	:	val_out <= 4'h14b5;
         4'hd783 	:	val_out <= 4'h14b5;
         4'hd788 	:	val_out <= 4'h14c2;
         4'hd789 	:	val_out <= 4'h14c2;
         4'hd78a 	:	val_out <= 4'h14c2;
         4'hd78b 	:	val_out <= 4'h14c2;
         4'hd790 	:	val_out <= 4'h14d0;
         4'hd791 	:	val_out <= 4'h14d0;
         4'hd792 	:	val_out <= 4'h14d0;
         4'hd793 	:	val_out <= 4'h14d0;
         4'hd798 	:	val_out <= 4'h14de;
         4'hd799 	:	val_out <= 4'h14de;
         4'hd79a 	:	val_out <= 4'h14de;
         4'hd79b 	:	val_out <= 4'h14de;
         4'hd7a0 	:	val_out <= 4'h14ec;
         4'hd7a1 	:	val_out <= 4'h14ec;
         4'hd7a2 	:	val_out <= 4'h14ec;
         4'hd7a3 	:	val_out <= 4'h14ec;
         4'hd7a8 	:	val_out <= 4'h14f9;
         4'hd7a9 	:	val_out <= 4'h14f9;
         4'hd7aa 	:	val_out <= 4'h14f9;
         4'hd7ab 	:	val_out <= 4'h14f9;
         4'hd7b0 	:	val_out <= 4'h1507;
         4'hd7b1 	:	val_out <= 4'h1507;
         4'hd7b2 	:	val_out <= 4'h1507;
         4'hd7b3 	:	val_out <= 4'h1507;
         4'hd7b8 	:	val_out <= 4'h1515;
         4'hd7b9 	:	val_out <= 4'h1515;
         4'hd7ba 	:	val_out <= 4'h1515;
         4'hd7bb 	:	val_out <= 4'h1515;
         4'hd7c0 	:	val_out <= 4'h1523;
         4'hd7c1 	:	val_out <= 4'h1523;
         4'hd7c2 	:	val_out <= 4'h1523;
         4'hd7c3 	:	val_out <= 4'h1523;
         4'hd7c8 	:	val_out <= 4'h1531;
         4'hd7c9 	:	val_out <= 4'h1531;
         4'hd7ca 	:	val_out <= 4'h1531;
         4'hd7cb 	:	val_out <= 4'h1531;
         4'hd7d0 	:	val_out <= 4'h153e;
         4'hd7d1 	:	val_out <= 4'h153e;
         4'hd7d2 	:	val_out <= 4'h153e;
         4'hd7d3 	:	val_out <= 4'h153e;
         4'hd7d8 	:	val_out <= 4'h154c;
         4'hd7d9 	:	val_out <= 4'h154c;
         4'hd7da 	:	val_out <= 4'h154c;
         4'hd7db 	:	val_out <= 4'h154c;
         4'hd7e0 	:	val_out <= 4'h155a;
         4'hd7e1 	:	val_out <= 4'h155a;
         4'hd7e2 	:	val_out <= 4'h155a;
         4'hd7e3 	:	val_out <= 4'h155a;
         4'hd7e8 	:	val_out <= 4'h1568;
         4'hd7e9 	:	val_out <= 4'h1568;
         4'hd7ea 	:	val_out <= 4'h1568;
         4'hd7eb 	:	val_out <= 4'h1568;
         4'hd7f0 	:	val_out <= 4'h1576;
         4'hd7f1 	:	val_out <= 4'h1576;
         4'hd7f2 	:	val_out <= 4'h1576;
         4'hd7f3 	:	val_out <= 4'h1576;
         4'hd7f8 	:	val_out <= 4'h1584;
         4'hd7f9 	:	val_out <= 4'h1584;
         4'hd7fa 	:	val_out <= 4'h1584;
         4'hd7fb 	:	val_out <= 4'h1584;
         4'hd800 	:	val_out <= 4'h1592;
         4'hd801 	:	val_out <= 4'h1592;
         4'hd802 	:	val_out <= 4'h1592;
         4'hd803 	:	val_out <= 4'h1592;
         4'hd808 	:	val_out <= 4'h15a0;
         4'hd809 	:	val_out <= 4'h15a0;
         4'hd80a 	:	val_out <= 4'h15a0;
         4'hd80b 	:	val_out <= 4'h15a0;
         4'hd810 	:	val_out <= 4'h15ae;
         4'hd811 	:	val_out <= 4'h15ae;
         4'hd812 	:	val_out <= 4'h15ae;
         4'hd813 	:	val_out <= 4'h15ae;
         4'hd818 	:	val_out <= 4'h15bc;
         4'hd819 	:	val_out <= 4'h15bc;
         4'hd81a 	:	val_out <= 4'h15bc;
         4'hd81b 	:	val_out <= 4'h15bc;
         4'hd820 	:	val_out <= 4'h15ca;
         4'hd821 	:	val_out <= 4'h15ca;
         4'hd822 	:	val_out <= 4'h15ca;
         4'hd823 	:	val_out <= 4'h15ca;
         4'hd828 	:	val_out <= 4'h15d8;
         4'hd829 	:	val_out <= 4'h15d8;
         4'hd82a 	:	val_out <= 4'h15d8;
         4'hd82b 	:	val_out <= 4'h15d8;
         4'hd830 	:	val_out <= 4'h15e6;
         4'hd831 	:	val_out <= 4'h15e6;
         4'hd832 	:	val_out <= 4'h15e6;
         4'hd833 	:	val_out <= 4'h15e6;
         4'hd838 	:	val_out <= 4'h15f4;
         4'hd839 	:	val_out <= 4'h15f4;
         4'hd83a 	:	val_out <= 4'h15f4;
         4'hd83b 	:	val_out <= 4'h15f4;
         4'hd840 	:	val_out <= 4'h1602;
         4'hd841 	:	val_out <= 4'h1602;
         4'hd842 	:	val_out <= 4'h1602;
         4'hd843 	:	val_out <= 4'h1602;
         4'hd848 	:	val_out <= 4'h1610;
         4'hd849 	:	val_out <= 4'h1610;
         4'hd84a 	:	val_out <= 4'h1610;
         4'hd84b 	:	val_out <= 4'h1610;
         4'hd850 	:	val_out <= 4'h161e;
         4'hd851 	:	val_out <= 4'h161e;
         4'hd852 	:	val_out <= 4'h161e;
         4'hd853 	:	val_out <= 4'h161e;
         4'hd858 	:	val_out <= 4'h162c;
         4'hd859 	:	val_out <= 4'h162c;
         4'hd85a 	:	val_out <= 4'h162c;
         4'hd85b 	:	val_out <= 4'h162c;
         4'hd860 	:	val_out <= 4'h163b;
         4'hd861 	:	val_out <= 4'h163b;
         4'hd862 	:	val_out <= 4'h163b;
         4'hd863 	:	val_out <= 4'h163b;
         4'hd868 	:	val_out <= 4'h1649;
         4'hd869 	:	val_out <= 4'h1649;
         4'hd86a 	:	val_out <= 4'h1649;
         4'hd86b 	:	val_out <= 4'h1649;
         4'hd870 	:	val_out <= 4'h1657;
         4'hd871 	:	val_out <= 4'h1657;
         4'hd872 	:	val_out <= 4'h1657;
         4'hd873 	:	val_out <= 4'h1657;
         4'hd878 	:	val_out <= 4'h1665;
         4'hd879 	:	val_out <= 4'h1665;
         4'hd87a 	:	val_out <= 4'h1665;
         4'hd87b 	:	val_out <= 4'h1665;
         4'hd880 	:	val_out <= 4'h1673;
         4'hd881 	:	val_out <= 4'h1673;
         4'hd882 	:	val_out <= 4'h1673;
         4'hd883 	:	val_out <= 4'h1673;
         4'hd888 	:	val_out <= 4'h1682;
         4'hd889 	:	val_out <= 4'h1682;
         4'hd88a 	:	val_out <= 4'h1682;
         4'hd88b 	:	val_out <= 4'h1682;
         4'hd890 	:	val_out <= 4'h1690;
         4'hd891 	:	val_out <= 4'h1690;
         4'hd892 	:	val_out <= 4'h1690;
         4'hd893 	:	val_out <= 4'h1690;
         4'hd898 	:	val_out <= 4'h169e;
         4'hd899 	:	val_out <= 4'h169e;
         4'hd89a 	:	val_out <= 4'h169e;
         4'hd89b 	:	val_out <= 4'h169e;
         4'hd8a0 	:	val_out <= 4'h16ac;
         4'hd8a1 	:	val_out <= 4'h16ac;
         4'hd8a2 	:	val_out <= 4'h16ac;
         4'hd8a3 	:	val_out <= 4'h16ac;
         4'hd8a8 	:	val_out <= 4'h16bb;
         4'hd8a9 	:	val_out <= 4'h16bb;
         4'hd8aa 	:	val_out <= 4'h16bb;
         4'hd8ab 	:	val_out <= 4'h16bb;
         4'hd8b0 	:	val_out <= 4'h16c9;
         4'hd8b1 	:	val_out <= 4'h16c9;
         4'hd8b2 	:	val_out <= 4'h16c9;
         4'hd8b3 	:	val_out <= 4'h16c9;
         4'hd8b8 	:	val_out <= 4'h16d7;
         4'hd8b9 	:	val_out <= 4'h16d7;
         4'hd8ba 	:	val_out <= 4'h16d7;
         4'hd8bb 	:	val_out <= 4'h16d7;
         4'hd8c0 	:	val_out <= 4'h16e6;
         4'hd8c1 	:	val_out <= 4'h16e6;
         4'hd8c2 	:	val_out <= 4'h16e6;
         4'hd8c3 	:	val_out <= 4'h16e6;
         4'hd8c8 	:	val_out <= 4'h16f4;
         4'hd8c9 	:	val_out <= 4'h16f4;
         4'hd8ca 	:	val_out <= 4'h16f4;
         4'hd8cb 	:	val_out <= 4'h16f4;
         4'hd8d0 	:	val_out <= 4'h1702;
         4'hd8d1 	:	val_out <= 4'h1702;
         4'hd8d2 	:	val_out <= 4'h1702;
         4'hd8d3 	:	val_out <= 4'h1702;
         4'hd8d8 	:	val_out <= 4'h1711;
         4'hd8d9 	:	val_out <= 4'h1711;
         4'hd8da 	:	val_out <= 4'h1711;
         4'hd8db 	:	val_out <= 4'h1711;
         4'hd8e0 	:	val_out <= 4'h171f;
         4'hd8e1 	:	val_out <= 4'h171f;
         4'hd8e2 	:	val_out <= 4'h171f;
         4'hd8e3 	:	val_out <= 4'h171f;
         4'hd8e8 	:	val_out <= 4'h172e;
         4'hd8e9 	:	val_out <= 4'h172e;
         4'hd8ea 	:	val_out <= 4'h172e;
         4'hd8eb 	:	val_out <= 4'h172e;
         4'hd8f0 	:	val_out <= 4'h173c;
         4'hd8f1 	:	val_out <= 4'h173c;
         4'hd8f2 	:	val_out <= 4'h173c;
         4'hd8f3 	:	val_out <= 4'h173c;
         4'hd8f8 	:	val_out <= 4'h174a;
         4'hd8f9 	:	val_out <= 4'h174a;
         4'hd8fa 	:	val_out <= 4'h174a;
         4'hd8fb 	:	val_out <= 4'h174a;
         4'hd900 	:	val_out <= 4'h1759;
         4'hd901 	:	val_out <= 4'h1759;
         4'hd902 	:	val_out <= 4'h1759;
         4'hd903 	:	val_out <= 4'h1759;
         4'hd908 	:	val_out <= 4'h1767;
         4'hd909 	:	val_out <= 4'h1767;
         4'hd90a 	:	val_out <= 4'h1767;
         4'hd90b 	:	val_out <= 4'h1767;
         4'hd910 	:	val_out <= 4'h1776;
         4'hd911 	:	val_out <= 4'h1776;
         4'hd912 	:	val_out <= 4'h1776;
         4'hd913 	:	val_out <= 4'h1776;
         4'hd918 	:	val_out <= 4'h1784;
         4'hd919 	:	val_out <= 4'h1784;
         4'hd91a 	:	val_out <= 4'h1784;
         4'hd91b 	:	val_out <= 4'h1784;
         4'hd920 	:	val_out <= 4'h1793;
         4'hd921 	:	val_out <= 4'h1793;
         4'hd922 	:	val_out <= 4'h1793;
         4'hd923 	:	val_out <= 4'h1793;
         4'hd928 	:	val_out <= 4'h17a1;
         4'hd929 	:	val_out <= 4'h17a1;
         4'hd92a 	:	val_out <= 4'h17a1;
         4'hd92b 	:	val_out <= 4'h17a1;
         4'hd930 	:	val_out <= 4'h17b0;
         4'hd931 	:	val_out <= 4'h17b0;
         4'hd932 	:	val_out <= 4'h17b0;
         4'hd933 	:	val_out <= 4'h17b0;
         4'hd938 	:	val_out <= 4'h17bf;
         4'hd939 	:	val_out <= 4'h17bf;
         4'hd93a 	:	val_out <= 4'h17bf;
         4'hd93b 	:	val_out <= 4'h17bf;
         4'hd940 	:	val_out <= 4'h17cd;
         4'hd941 	:	val_out <= 4'h17cd;
         4'hd942 	:	val_out <= 4'h17cd;
         4'hd943 	:	val_out <= 4'h17cd;
         4'hd948 	:	val_out <= 4'h17dc;
         4'hd949 	:	val_out <= 4'h17dc;
         4'hd94a 	:	val_out <= 4'h17dc;
         4'hd94b 	:	val_out <= 4'h17dc;
         4'hd950 	:	val_out <= 4'h17ea;
         4'hd951 	:	val_out <= 4'h17ea;
         4'hd952 	:	val_out <= 4'h17ea;
         4'hd953 	:	val_out <= 4'h17ea;
         4'hd958 	:	val_out <= 4'h17f9;
         4'hd959 	:	val_out <= 4'h17f9;
         4'hd95a 	:	val_out <= 4'h17f9;
         4'hd95b 	:	val_out <= 4'h17f9;
         4'hd960 	:	val_out <= 4'h1808;
         4'hd961 	:	val_out <= 4'h1808;
         4'hd962 	:	val_out <= 4'h1808;
         4'hd963 	:	val_out <= 4'h1808;
         4'hd968 	:	val_out <= 4'h1816;
         4'hd969 	:	val_out <= 4'h1816;
         4'hd96a 	:	val_out <= 4'h1816;
         4'hd96b 	:	val_out <= 4'h1816;
         4'hd970 	:	val_out <= 4'h1825;
         4'hd971 	:	val_out <= 4'h1825;
         4'hd972 	:	val_out <= 4'h1825;
         4'hd973 	:	val_out <= 4'h1825;
         4'hd978 	:	val_out <= 4'h1834;
         4'hd979 	:	val_out <= 4'h1834;
         4'hd97a 	:	val_out <= 4'h1834;
         4'hd97b 	:	val_out <= 4'h1834;
         4'hd980 	:	val_out <= 4'h1842;
         4'hd981 	:	val_out <= 4'h1842;
         4'hd982 	:	val_out <= 4'h1842;
         4'hd983 	:	val_out <= 4'h1842;
         4'hd988 	:	val_out <= 4'h1851;
         4'hd989 	:	val_out <= 4'h1851;
         4'hd98a 	:	val_out <= 4'h1851;
         4'hd98b 	:	val_out <= 4'h1851;
         4'hd990 	:	val_out <= 4'h1860;
         4'hd991 	:	val_out <= 4'h1860;
         4'hd992 	:	val_out <= 4'h1860;
         4'hd993 	:	val_out <= 4'h1860;
         4'hd998 	:	val_out <= 4'h186f;
         4'hd999 	:	val_out <= 4'h186f;
         4'hd99a 	:	val_out <= 4'h186f;
         4'hd99b 	:	val_out <= 4'h186f;
         4'hd9a0 	:	val_out <= 4'h187d;
         4'hd9a1 	:	val_out <= 4'h187d;
         4'hd9a2 	:	val_out <= 4'h187d;
         4'hd9a3 	:	val_out <= 4'h187d;
         4'hd9a8 	:	val_out <= 4'h188c;
         4'hd9a9 	:	val_out <= 4'h188c;
         4'hd9aa 	:	val_out <= 4'h188c;
         4'hd9ab 	:	val_out <= 4'h188c;
         4'hd9b0 	:	val_out <= 4'h189b;
         4'hd9b1 	:	val_out <= 4'h189b;
         4'hd9b2 	:	val_out <= 4'h189b;
         4'hd9b3 	:	val_out <= 4'h189b;
         4'hd9b8 	:	val_out <= 4'h18aa;
         4'hd9b9 	:	val_out <= 4'h18aa;
         4'hd9ba 	:	val_out <= 4'h18aa;
         4'hd9bb 	:	val_out <= 4'h18aa;
         4'hd9c0 	:	val_out <= 4'h18b9;
         4'hd9c1 	:	val_out <= 4'h18b9;
         4'hd9c2 	:	val_out <= 4'h18b9;
         4'hd9c3 	:	val_out <= 4'h18b9;
         4'hd9c8 	:	val_out <= 4'h18c8;
         4'hd9c9 	:	val_out <= 4'h18c8;
         4'hd9ca 	:	val_out <= 4'h18c8;
         4'hd9cb 	:	val_out <= 4'h18c8;
         4'hd9d0 	:	val_out <= 4'h18d6;
         4'hd9d1 	:	val_out <= 4'h18d6;
         4'hd9d2 	:	val_out <= 4'h18d6;
         4'hd9d3 	:	val_out <= 4'h18d6;
         4'hd9d8 	:	val_out <= 4'h18e5;
         4'hd9d9 	:	val_out <= 4'h18e5;
         4'hd9da 	:	val_out <= 4'h18e5;
         4'hd9db 	:	val_out <= 4'h18e5;
         4'hd9e0 	:	val_out <= 4'h18f4;
         4'hd9e1 	:	val_out <= 4'h18f4;
         4'hd9e2 	:	val_out <= 4'h18f4;
         4'hd9e3 	:	val_out <= 4'h18f4;
         4'hd9e8 	:	val_out <= 4'h1903;
         4'hd9e9 	:	val_out <= 4'h1903;
         4'hd9ea 	:	val_out <= 4'h1903;
         4'hd9eb 	:	val_out <= 4'h1903;
         4'hd9f0 	:	val_out <= 4'h1912;
         4'hd9f1 	:	val_out <= 4'h1912;
         4'hd9f2 	:	val_out <= 4'h1912;
         4'hd9f3 	:	val_out <= 4'h1912;
         4'hd9f8 	:	val_out <= 4'h1921;
         4'hd9f9 	:	val_out <= 4'h1921;
         4'hd9fa 	:	val_out <= 4'h1921;
         4'hd9fb 	:	val_out <= 4'h1921;
         4'hda00 	:	val_out <= 4'h1930;
         4'hda01 	:	val_out <= 4'h1930;
         4'hda02 	:	val_out <= 4'h1930;
         4'hda03 	:	val_out <= 4'h1930;
         4'hda08 	:	val_out <= 4'h193f;
         4'hda09 	:	val_out <= 4'h193f;
         4'hda0a 	:	val_out <= 4'h193f;
         4'hda0b 	:	val_out <= 4'h193f;
         4'hda10 	:	val_out <= 4'h194e;
         4'hda11 	:	val_out <= 4'h194e;
         4'hda12 	:	val_out <= 4'h194e;
         4'hda13 	:	val_out <= 4'h194e;
         4'hda18 	:	val_out <= 4'h195d;
         4'hda19 	:	val_out <= 4'h195d;
         4'hda1a 	:	val_out <= 4'h195d;
         4'hda1b 	:	val_out <= 4'h195d;
         4'hda20 	:	val_out <= 4'h196c;
         4'hda21 	:	val_out <= 4'h196c;
         4'hda22 	:	val_out <= 4'h196c;
         4'hda23 	:	val_out <= 4'h196c;
         4'hda28 	:	val_out <= 4'h197b;
         4'hda29 	:	val_out <= 4'h197b;
         4'hda2a 	:	val_out <= 4'h197b;
         4'hda2b 	:	val_out <= 4'h197b;
         4'hda30 	:	val_out <= 4'h198a;
         4'hda31 	:	val_out <= 4'h198a;
         4'hda32 	:	val_out <= 4'h198a;
         4'hda33 	:	val_out <= 4'h198a;
         4'hda38 	:	val_out <= 4'h1999;
         4'hda39 	:	val_out <= 4'h1999;
         4'hda3a 	:	val_out <= 4'h1999;
         4'hda3b 	:	val_out <= 4'h1999;
         4'hda40 	:	val_out <= 4'h19a8;
         4'hda41 	:	val_out <= 4'h19a8;
         4'hda42 	:	val_out <= 4'h19a8;
         4'hda43 	:	val_out <= 4'h19a8;
         4'hda48 	:	val_out <= 4'h19b7;
         4'hda49 	:	val_out <= 4'h19b7;
         4'hda4a 	:	val_out <= 4'h19b7;
         4'hda4b 	:	val_out <= 4'h19b7;
         4'hda50 	:	val_out <= 4'h19c6;
         4'hda51 	:	val_out <= 4'h19c6;
         4'hda52 	:	val_out <= 4'h19c6;
         4'hda53 	:	val_out <= 4'h19c6;
         4'hda58 	:	val_out <= 4'h19d6;
         4'hda59 	:	val_out <= 4'h19d6;
         4'hda5a 	:	val_out <= 4'h19d6;
         4'hda5b 	:	val_out <= 4'h19d6;
         4'hda60 	:	val_out <= 4'h19e5;
         4'hda61 	:	val_out <= 4'h19e5;
         4'hda62 	:	val_out <= 4'h19e5;
         4'hda63 	:	val_out <= 4'h19e5;
         4'hda68 	:	val_out <= 4'h19f4;
         4'hda69 	:	val_out <= 4'h19f4;
         4'hda6a 	:	val_out <= 4'h19f4;
         4'hda6b 	:	val_out <= 4'h19f4;
         4'hda70 	:	val_out <= 4'h1a03;
         4'hda71 	:	val_out <= 4'h1a03;
         4'hda72 	:	val_out <= 4'h1a03;
         4'hda73 	:	val_out <= 4'h1a03;
         4'hda78 	:	val_out <= 4'h1a12;
         4'hda79 	:	val_out <= 4'h1a12;
         4'hda7a 	:	val_out <= 4'h1a12;
         4'hda7b 	:	val_out <= 4'h1a12;
         4'hda80 	:	val_out <= 4'h1a22;
         4'hda81 	:	val_out <= 4'h1a22;
         4'hda82 	:	val_out <= 4'h1a22;
         4'hda83 	:	val_out <= 4'h1a22;
         4'hda88 	:	val_out <= 4'h1a31;
         4'hda89 	:	val_out <= 4'h1a31;
         4'hda8a 	:	val_out <= 4'h1a31;
         4'hda8b 	:	val_out <= 4'h1a31;
         4'hda90 	:	val_out <= 4'h1a40;
         4'hda91 	:	val_out <= 4'h1a40;
         4'hda92 	:	val_out <= 4'h1a40;
         4'hda93 	:	val_out <= 4'h1a40;
         4'hda98 	:	val_out <= 4'h1a4f;
         4'hda99 	:	val_out <= 4'h1a4f;
         4'hda9a 	:	val_out <= 4'h1a4f;
         4'hda9b 	:	val_out <= 4'h1a4f;
         4'hdaa0 	:	val_out <= 4'h1a5f;
         4'hdaa1 	:	val_out <= 4'h1a5f;
         4'hdaa2 	:	val_out <= 4'h1a5f;
         4'hdaa3 	:	val_out <= 4'h1a5f;
         4'hdaa8 	:	val_out <= 4'h1a6e;
         4'hdaa9 	:	val_out <= 4'h1a6e;
         4'hdaaa 	:	val_out <= 4'h1a6e;
         4'hdaab 	:	val_out <= 4'h1a6e;
         4'hdab0 	:	val_out <= 4'h1a7d;
         4'hdab1 	:	val_out <= 4'h1a7d;
         4'hdab2 	:	val_out <= 4'h1a7d;
         4'hdab3 	:	val_out <= 4'h1a7d;
         4'hdab8 	:	val_out <= 4'h1a8c;
         4'hdab9 	:	val_out <= 4'h1a8c;
         4'hdaba 	:	val_out <= 4'h1a8c;
         4'hdabb 	:	val_out <= 4'h1a8c;
         4'hdac0 	:	val_out <= 4'h1a9c;
         4'hdac1 	:	val_out <= 4'h1a9c;
         4'hdac2 	:	val_out <= 4'h1a9c;
         4'hdac3 	:	val_out <= 4'h1a9c;
         4'hdac8 	:	val_out <= 4'h1aab;
         4'hdac9 	:	val_out <= 4'h1aab;
         4'hdaca 	:	val_out <= 4'h1aab;
         4'hdacb 	:	val_out <= 4'h1aab;
         4'hdad0 	:	val_out <= 4'h1aba;
         4'hdad1 	:	val_out <= 4'h1aba;
         4'hdad2 	:	val_out <= 4'h1aba;
         4'hdad3 	:	val_out <= 4'h1aba;
         4'hdad8 	:	val_out <= 4'h1aca;
         4'hdad9 	:	val_out <= 4'h1aca;
         4'hdada 	:	val_out <= 4'h1aca;
         4'hdadb 	:	val_out <= 4'h1aca;
         4'hdae0 	:	val_out <= 4'h1ad9;
         4'hdae1 	:	val_out <= 4'h1ad9;
         4'hdae2 	:	val_out <= 4'h1ad9;
         4'hdae3 	:	val_out <= 4'h1ad9;
         4'hdae8 	:	val_out <= 4'h1ae9;
         4'hdae9 	:	val_out <= 4'h1ae9;
         4'hdaea 	:	val_out <= 4'h1ae9;
         4'hdaeb 	:	val_out <= 4'h1ae9;
         4'hdaf0 	:	val_out <= 4'h1af8;
         4'hdaf1 	:	val_out <= 4'h1af8;
         4'hdaf2 	:	val_out <= 4'h1af8;
         4'hdaf3 	:	val_out <= 4'h1af8;
         4'hdaf8 	:	val_out <= 4'h1b08;
         4'hdaf9 	:	val_out <= 4'h1b08;
         4'hdafa 	:	val_out <= 4'h1b08;
         4'hdafb 	:	val_out <= 4'h1b08;
         4'hdb00 	:	val_out <= 4'h1b17;
         4'hdb01 	:	val_out <= 4'h1b17;
         4'hdb02 	:	val_out <= 4'h1b17;
         4'hdb03 	:	val_out <= 4'h1b17;
         4'hdb08 	:	val_out <= 4'h1b26;
         4'hdb09 	:	val_out <= 4'h1b26;
         4'hdb0a 	:	val_out <= 4'h1b26;
         4'hdb0b 	:	val_out <= 4'h1b26;
         4'hdb10 	:	val_out <= 4'h1b36;
         4'hdb11 	:	val_out <= 4'h1b36;
         4'hdb12 	:	val_out <= 4'h1b36;
         4'hdb13 	:	val_out <= 4'h1b36;
         4'hdb18 	:	val_out <= 4'h1b45;
         4'hdb19 	:	val_out <= 4'h1b45;
         4'hdb1a 	:	val_out <= 4'h1b45;
         4'hdb1b 	:	val_out <= 4'h1b45;
         4'hdb20 	:	val_out <= 4'h1b55;
         4'hdb21 	:	val_out <= 4'h1b55;
         4'hdb22 	:	val_out <= 4'h1b55;
         4'hdb23 	:	val_out <= 4'h1b55;
         4'hdb28 	:	val_out <= 4'h1b64;
         4'hdb29 	:	val_out <= 4'h1b64;
         4'hdb2a 	:	val_out <= 4'h1b64;
         4'hdb2b 	:	val_out <= 4'h1b64;
         4'hdb30 	:	val_out <= 4'h1b74;
         4'hdb31 	:	val_out <= 4'h1b74;
         4'hdb32 	:	val_out <= 4'h1b74;
         4'hdb33 	:	val_out <= 4'h1b74;
         4'hdb38 	:	val_out <= 4'h1b84;
         4'hdb39 	:	val_out <= 4'h1b84;
         4'hdb3a 	:	val_out <= 4'h1b84;
         4'hdb3b 	:	val_out <= 4'h1b84;
         4'hdb40 	:	val_out <= 4'h1b93;
         4'hdb41 	:	val_out <= 4'h1b93;
         4'hdb42 	:	val_out <= 4'h1b93;
         4'hdb43 	:	val_out <= 4'h1b93;
         4'hdb48 	:	val_out <= 4'h1ba3;
         4'hdb49 	:	val_out <= 4'h1ba3;
         4'hdb4a 	:	val_out <= 4'h1ba3;
         4'hdb4b 	:	val_out <= 4'h1ba3;
         4'hdb50 	:	val_out <= 4'h1bb2;
         4'hdb51 	:	val_out <= 4'h1bb2;
         4'hdb52 	:	val_out <= 4'h1bb2;
         4'hdb53 	:	val_out <= 4'h1bb2;
         4'hdb58 	:	val_out <= 4'h1bc2;
         4'hdb59 	:	val_out <= 4'h1bc2;
         4'hdb5a 	:	val_out <= 4'h1bc2;
         4'hdb5b 	:	val_out <= 4'h1bc2;
         4'hdb60 	:	val_out <= 4'h1bd2;
         4'hdb61 	:	val_out <= 4'h1bd2;
         4'hdb62 	:	val_out <= 4'h1bd2;
         4'hdb63 	:	val_out <= 4'h1bd2;
         4'hdb68 	:	val_out <= 4'h1be1;
         4'hdb69 	:	val_out <= 4'h1be1;
         4'hdb6a 	:	val_out <= 4'h1be1;
         4'hdb6b 	:	val_out <= 4'h1be1;
         4'hdb70 	:	val_out <= 4'h1bf1;
         4'hdb71 	:	val_out <= 4'h1bf1;
         4'hdb72 	:	val_out <= 4'h1bf1;
         4'hdb73 	:	val_out <= 4'h1bf1;
         4'hdb78 	:	val_out <= 4'h1c01;
         4'hdb79 	:	val_out <= 4'h1c01;
         4'hdb7a 	:	val_out <= 4'h1c01;
         4'hdb7b 	:	val_out <= 4'h1c01;
         4'hdb80 	:	val_out <= 4'h1c10;
         4'hdb81 	:	val_out <= 4'h1c10;
         4'hdb82 	:	val_out <= 4'h1c10;
         4'hdb83 	:	val_out <= 4'h1c10;
         4'hdb88 	:	val_out <= 4'h1c20;
         4'hdb89 	:	val_out <= 4'h1c20;
         4'hdb8a 	:	val_out <= 4'h1c20;
         4'hdb8b 	:	val_out <= 4'h1c20;
         4'hdb90 	:	val_out <= 4'h1c30;
         4'hdb91 	:	val_out <= 4'h1c30;
         4'hdb92 	:	val_out <= 4'h1c30;
         4'hdb93 	:	val_out <= 4'h1c30;
         4'hdb98 	:	val_out <= 4'h1c3f;
         4'hdb99 	:	val_out <= 4'h1c3f;
         4'hdb9a 	:	val_out <= 4'h1c3f;
         4'hdb9b 	:	val_out <= 4'h1c3f;
         4'hdba0 	:	val_out <= 4'h1c4f;
         4'hdba1 	:	val_out <= 4'h1c4f;
         4'hdba2 	:	val_out <= 4'h1c4f;
         4'hdba3 	:	val_out <= 4'h1c4f;
         4'hdba8 	:	val_out <= 4'h1c5f;
         4'hdba9 	:	val_out <= 4'h1c5f;
         4'hdbaa 	:	val_out <= 4'h1c5f;
         4'hdbab 	:	val_out <= 4'h1c5f;
         4'hdbb0 	:	val_out <= 4'h1c6f;
         4'hdbb1 	:	val_out <= 4'h1c6f;
         4'hdbb2 	:	val_out <= 4'h1c6f;
         4'hdbb3 	:	val_out <= 4'h1c6f;
         4'hdbb8 	:	val_out <= 4'h1c7f;
         4'hdbb9 	:	val_out <= 4'h1c7f;
         4'hdbba 	:	val_out <= 4'h1c7f;
         4'hdbbb 	:	val_out <= 4'h1c7f;
         4'hdbc0 	:	val_out <= 4'h1c8e;
         4'hdbc1 	:	val_out <= 4'h1c8e;
         4'hdbc2 	:	val_out <= 4'h1c8e;
         4'hdbc3 	:	val_out <= 4'h1c8e;
         4'hdbc8 	:	val_out <= 4'h1c9e;
         4'hdbc9 	:	val_out <= 4'h1c9e;
         4'hdbca 	:	val_out <= 4'h1c9e;
         4'hdbcb 	:	val_out <= 4'h1c9e;
         4'hdbd0 	:	val_out <= 4'h1cae;
         4'hdbd1 	:	val_out <= 4'h1cae;
         4'hdbd2 	:	val_out <= 4'h1cae;
         4'hdbd3 	:	val_out <= 4'h1cae;
         4'hdbd8 	:	val_out <= 4'h1cbe;
         4'hdbd9 	:	val_out <= 4'h1cbe;
         4'hdbda 	:	val_out <= 4'h1cbe;
         4'hdbdb 	:	val_out <= 4'h1cbe;
         4'hdbe0 	:	val_out <= 4'h1cce;
         4'hdbe1 	:	val_out <= 4'h1cce;
         4'hdbe2 	:	val_out <= 4'h1cce;
         4'hdbe3 	:	val_out <= 4'h1cce;
         4'hdbe8 	:	val_out <= 4'h1cde;
         4'hdbe9 	:	val_out <= 4'h1cde;
         4'hdbea 	:	val_out <= 4'h1cde;
         4'hdbeb 	:	val_out <= 4'h1cde;
         4'hdbf0 	:	val_out <= 4'h1cee;
         4'hdbf1 	:	val_out <= 4'h1cee;
         4'hdbf2 	:	val_out <= 4'h1cee;
         4'hdbf3 	:	val_out <= 4'h1cee;
         4'hdbf8 	:	val_out <= 4'h1cfe;
         4'hdbf9 	:	val_out <= 4'h1cfe;
         4'hdbfa 	:	val_out <= 4'h1cfe;
         4'hdbfb 	:	val_out <= 4'h1cfe;
         4'hdc00 	:	val_out <= 4'h1d0d;
         4'hdc01 	:	val_out <= 4'h1d0d;
         4'hdc02 	:	val_out <= 4'h1d0d;
         4'hdc03 	:	val_out <= 4'h1d0d;
         4'hdc08 	:	val_out <= 4'h1d1d;
         4'hdc09 	:	val_out <= 4'h1d1d;
         4'hdc0a 	:	val_out <= 4'h1d1d;
         4'hdc0b 	:	val_out <= 4'h1d1d;
         4'hdc10 	:	val_out <= 4'h1d2d;
         4'hdc11 	:	val_out <= 4'h1d2d;
         4'hdc12 	:	val_out <= 4'h1d2d;
         4'hdc13 	:	val_out <= 4'h1d2d;
         4'hdc18 	:	val_out <= 4'h1d3d;
         4'hdc19 	:	val_out <= 4'h1d3d;
         4'hdc1a 	:	val_out <= 4'h1d3d;
         4'hdc1b 	:	val_out <= 4'h1d3d;
         4'hdc20 	:	val_out <= 4'h1d4d;
         4'hdc21 	:	val_out <= 4'h1d4d;
         4'hdc22 	:	val_out <= 4'h1d4d;
         4'hdc23 	:	val_out <= 4'h1d4d;
         4'hdc28 	:	val_out <= 4'h1d5d;
         4'hdc29 	:	val_out <= 4'h1d5d;
         4'hdc2a 	:	val_out <= 4'h1d5d;
         4'hdc2b 	:	val_out <= 4'h1d5d;
         4'hdc30 	:	val_out <= 4'h1d6d;
         4'hdc31 	:	val_out <= 4'h1d6d;
         4'hdc32 	:	val_out <= 4'h1d6d;
         4'hdc33 	:	val_out <= 4'h1d6d;
         4'hdc38 	:	val_out <= 4'h1d7d;
         4'hdc39 	:	val_out <= 4'h1d7d;
         4'hdc3a 	:	val_out <= 4'h1d7d;
         4'hdc3b 	:	val_out <= 4'h1d7d;
         4'hdc40 	:	val_out <= 4'h1d8e;
         4'hdc41 	:	val_out <= 4'h1d8e;
         4'hdc42 	:	val_out <= 4'h1d8e;
         4'hdc43 	:	val_out <= 4'h1d8e;
         4'hdc48 	:	val_out <= 4'h1d9e;
         4'hdc49 	:	val_out <= 4'h1d9e;
         4'hdc4a 	:	val_out <= 4'h1d9e;
         4'hdc4b 	:	val_out <= 4'h1d9e;
         4'hdc50 	:	val_out <= 4'h1dae;
         4'hdc51 	:	val_out <= 4'h1dae;
         4'hdc52 	:	val_out <= 4'h1dae;
         4'hdc53 	:	val_out <= 4'h1dae;
         4'hdc58 	:	val_out <= 4'h1dbe;
         4'hdc59 	:	val_out <= 4'h1dbe;
         4'hdc5a 	:	val_out <= 4'h1dbe;
         4'hdc5b 	:	val_out <= 4'h1dbe;
         4'hdc60 	:	val_out <= 4'h1dce;
         4'hdc61 	:	val_out <= 4'h1dce;
         4'hdc62 	:	val_out <= 4'h1dce;
         4'hdc63 	:	val_out <= 4'h1dce;
         4'hdc68 	:	val_out <= 4'h1dde;
         4'hdc69 	:	val_out <= 4'h1dde;
         4'hdc6a 	:	val_out <= 4'h1dde;
         4'hdc6b 	:	val_out <= 4'h1dde;
         4'hdc70 	:	val_out <= 4'h1dee;
         4'hdc71 	:	val_out <= 4'h1dee;
         4'hdc72 	:	val_out <= 4'h1dee;
         4'hdc73 	:	val_out <= 4'h1dee;
         4'hdc78 	:	val_out <= 4'h1dfe;
         4'hdc79 	:	val_out <= 4'h1dfe;
         4'hdc7a 	:	val_out <= 4'h1dfe;
         4'hdc7b 	:	val_out <= 4'h1dfe;
         4'hdc80 	:	val_out <= 4'h1e0e;
         4'hdc81 	:	val_out <= 4'h1e0e;
         4'hdc82 	:	val_out <= 4'h1e0e;
         4'hdc83 	:	val_out <= 4'h1e0e;
         4'hdc88 	:	val_out <= 4'h1e1f;
         4'hdc89 	:	val_out <= 4'h1e1f;
         4'hdc8a 	:	val_out <= 4'h1e1f;
         4'hdc8b 	:	val_out <= 4'h1e1f;
         4'hdc90 	:	val_out <= 4'h1e2f;
         4'hdc91 	:	val_out <= 4'h1e2f;
         4'hdc92 	:	val_out <= 4'h1e2f;
         4'hdc93 	:	val_out <= 4'h1e2f;
         4'hdc98 	:	val_out <= 4'h1e3f;
         4'hdc99 	:	val_out <= 4'h1e3f;
         4'hdc9a 	:	val_out <= 4'h1e3f;
         4'hdc9b 	:	val_out <= 4'h1e3f;
         4'hdca0 	:	val_out <= 4'h1e4f;
         4'hdca1 	:	val_out <= 4'h1e4f;
         4'hdca2 	:	val_out <= 4'h1e4f;
         4'hdca3 	:	val_out <= 4'h1e4f;
         4'hdca8 	:	val_out <= 4'h1e60;
         4'hdca9 	:	val_out <= 4'h1e60;
         4'hdcaa 	:	val_out <= 4'h1e60;
         4'hdcab 	:	val_out <= 4'h1e60;
         4'hdcb0 	:	val_out <= 4'h1e70;
         4'hdcb1 	:	val_out <= 4'h1e70;
         4'hdcb2 	:	val_out <= 4'h1e70;
         4'hdcb3 	:	val_out <= 4'h1e70;
         4'hdcb8 	:	val_out <= 4'h1e80;
         4'hdcb9 	:	val_out <= 4'h1e80;
         4'hdcba 	:	val_out <= 4'h1e80;
         4'hdcbb 	:	val_out <= 4'h1e80;
         4'hdcc0 	:	val_out <= 4'h1e90;
         4'hdcc1 	:	val_out <= 4'h1e90;
         4'hdcc2 	:	val_out <= 4'h1e90;
         4'hdcc3 	:	val_out <= 4'h1e90;
         4'hdcc8 	:	val_out <= 4'h1ea1;
         4'hdcc9 	:	val_out <= 4'h1ea1;
         4'hdcca 	:	val_out <= 4'h1ea1;
         4'hdccb 	:	val_out <= 4'h1ea1;
         4'hdcd0 	:	val_out <= 4'h1eb1;
         4'hdcd1 	:	val_out <= 4'h1eb1;
         4'hdcd2 	:	val_out <= 4'h1eb1;
         4'hdcd3 	:	val_out <= 4'h1eb1;
         4'hdcd8 	:	val_out <= 4'h1ec1;
         4'hdcd9 	:	val_out <= 4'h1ec1;
         4'hdcda 	:	val_out <= 4'h1ec1;
         4'hdcdb 	:	val_out <= 4'h1ec1;
         4'hdce0 	:	val_out <= 4'h1ed2;
         4'hdce1 	:	val_out <= 4'h1ed2;
         4'hdce2 	:	val_out <= 4'h1ed2;
         4'hdce3 	:	val_out <= 4'h1ed2;
         4'hdce8 	:	val_out <= 4'h1ee2;
         4'hdce9 	:	val_out <= 4'h1ee2;
         4'hdcea 	:	val_out <= 4'h1ee2;
         4'hdceb 	:	val_out <= 4'h1ee2;
         4'hdcf0 	:	val_out <= 4'h1ef2;
         4'hdcf1 	:	val_out <= 4'h1ef2;
         4'hdcf2 	:	val_out <= 4'h1ef2;
         4'hdcf3 	:	val_out <= 4'h1ef2;
         4'hdcf8 	:	val_out <= 4'h1f03;
         4'hdcf9 	:	val_out <= 4'h1f03;
         4'hdcfa 	:	val_out <= 4'h1f03;
         4'hdcfb 	:	val_out <= 4'h1f03;
         4'hdd00 	:	val_out <= 4'h1f13;
         4'hdd01 	:	val_out <= 4'h1f13;
         4'hdd02 	:	val_out <= 4'h1f13;
         4'hdd03 	:	val_out <= 4'h1f13;
         4'hdd08 	:	val_out <= 4'h1f24;
         4'hdd09 	:	val_out <= 4'h1f24;
         4'hdd0a 	:	val_out <= 4'h1f24;
         4'hdd0b 	:	val_out <= 4'h1f24;
         4'hdd10 	:	val_out <= 4'h1f34;
         4'hdd11 	:	val_out <= 4'h1f34;
         4'hdd12 	:	val_out <= 4'h1f34;
         4'hdd13 	:	val_out <= 4'h1f34;
         4'hdd18 	:	val_out <= 4'h1f45;
         4'hdd19 	:	val_out <= 4'h1f45;
         4'hdd1a 	:	val_out <= 4'h1f45;
         4'hdd1b 	:	val_out <= 4'h1f45;
         4'hdd20 	:	val_out <= 4'h1f55;
         4'hdd21 	:	val_out <= 4'h1f55;
         4'hdd22 	:	val_out <= 4'h1f55;
         4'hdd23 	:	val_out <= 4'h1f55;
         4'hdd28 	:	val_out <= 4'h1f66;
         4'hdd29 	:	val_out <= 4'h1f66;
         4'hdd2a 	:	val_out <= 4'h1f66;
         4'hdd2b 	:	val_out <= 4'h1f66;
         4'hdd30 	:	val_out <= 4'h1f76;
         4'hdd31 	:	val_out <= 4'h1f76;
         4'hdd32 	:	val_out <= 4'h1f76;
         4'hdd33 	:	val_out <= 4'h1f76;
         4'hdd38 	:	val_out <= 4'h1f87;
         4'hdd39 	:	val_out <= 4'h1f87;
         4'hdd3a 	:	val_out <= 4'h1f87;
         4'hdd3b 	:	val_out <= 4'h1f87;
         4'hdd40 	:	val_out <= 4'h1f97;
         4'hdd41 	:	val_out <= 4'h1f97;
         4'hdd42 	:	val_out <= 4'h1f97;
         4'hdd43 	:	val_out <= 4'h1f97;
         4'hdd48 	:	val_out <= 4'h1fa8;
         4'hdd49 	:	val_out <= 4'h1fa8;
         4'hdd4a 	:	val_out <= 4'h1fa8;
         4'hdd4b 	:	val_out <= 4'h1fa8;
         4'hdd50 	:	val_out <= 4'h1fb8;
         4'hdd51 	:	val_out <= 4'h1fb8;
         4'hdd52 	:	val_out <= 4'h1fb8;
         4'hdd53 	:	val_out <= 4'h1fb8;
         4'hdd58 	:	val_out <= 4'h1fc9;
         4'hdd59 	:	val_out <= 4'h1fc9;
         4'hdd5a 	:	val_out <= 4'h1fc9;
         4'hdd5b 	:	val_out <= 4'h1fc9;
         4'hdd60 	:	val_out <= 4'h1fd9;
         4'hdd61 	:	val_out <= 4'h1fd9;
         4'hdd62 	:	val_out <= 4'h1fd9;
         4'hdd63 	:	val_out <= 4'h1fd9;
         4'hdd68 	:	val_out <= 4'h1fea;
         4'hdd69 	:	val_out <= 4'h1fea;
         4'hdd6a 	:	val_out <= 4'h1fea;
         4'hdd6b 	:	val_out <= 4'h1fea;
         4'hdd70 	:	val_out <= 4'h1ffb;
         4'hdd71 	:	val_out <= 4'h1ffb;
         4'hdd72 	:	val_out <= 4'h1ffb;
         4'hdd73 	:	val_out <= 4'h1ffb;
         4'hdd78 	:	val_out <= 4'h200b;
         4'hdd79 	:	val_out <= 4'h200b;
         4'hdd7a 	:	val_out <= 4'h200b;
         4'hdd7b 	:	val_out <= 4'h200b;
         4'hdd80 	:	val_out <= 4'h201c;
         4'hdd81 	:	val_out <= 4'h201c;
         4'hdd82 	:	val_out <= 4'h201c;
         4'hdd83 	:	val_out <= 4'h201c;
         4'hdd88 	:	val_out <= 4'h202c;
         4'hdd89 	:	val_out <= 4'h202c;
         4'hdd8a 	:	val_out <= 4'h202c;
         4'hdd8b 	:	val_out <= 4'h202c;
         4'hdd90 	:	val_out <= 4'h203d;
         4'hdd91 	:	val_out <= 4'h203d;
         4'hdd92 	:	val_out <= 4'h203d;
         4'hdd93 	:	val_out <= 4'h203d;
         4'hdd98 	:	val_out <= 4'h204e;
         4'hdd99 	:	val_out <= 4'h204e;
         4'hdd9a 	:	val_out <= 4'h204e;
         4'hdd9b 	:	val_out <= 4'h204e;
         4'hdda0 	:	val_out <= 4'h205f;
         4'hdda1 	:	val_out <= 4'h205f;
         4'hdda2 	:	val_out <= 4'h205f;
         4'hdda3 	:	val_out <= 4'h205f;
         4'hdda8 	:	val_out <= 4'h206f;
         4'hdda9 	:	val_out <= 4'h206f;
         4'hddaa 	:	val_out <= 4'h206f;
         4'hddab 	:	val_out <= 4'h206f;
         4'hddb0 	:	val_out <= 4'h2080;
         4'hddb1 	:	val_out <= 4'h2080;
         4'hddb2 	:	val_out <= 4'h2080;
         4'hddb3 	:	val_out <= 4'h2080;
         4'hddb8 	:	val_out <= 4'h2091;
         4'hddb9 	:	val_out <= 4'h2091;
         4'hddba 	:	val_out <= 4'h2091;
         4'hddbb 	:	val_out <= 4'h2091;
         4'hddc0 	:	val_out <= 4'h20a1;
         4'hddc1 	:	val_out <= 4'h20a1;
         4'hddc2 	:	val_out <= 4'h20a1;
         4'hddc3 	:	val_out <= 4'h20a1;
         4'hddc8 	:	val_out <= 4'h20b2;
         4'hddc9 	:	val_out <= 4'h20b2;
         4'hddca 	:	val_out <= 4'h20b2;
         4'hddcb 	:	val_out <= 4'h20b2;
         4'hddd0 	:	val_out <= 4'h20c3;
         4'hddd1 	:	val_out <= 4'h20c3;
         4'hddd2 	:	val_out <= 4'h20c3;
         4'hddd3 	:	val_out <= 4'h20c3;
         4'hddd8 	:	val_out <= 4'h20d4;
         4'hddd9 	:	val_out <= 4'h20d4;
         4'hddda 	:	val_out <= 4'h20d4;
         4'hdddb 	:	val_out <= 4'h20d4;
         4'hdde0 	:	val_out <= 4'h20e5;
         4'hdde1 	:	val_out <= 4'h20e5;
         4'hdde2 	:	val_out <= 4'h20e5;
         4'hdde3 	:	val_out <= 4'h20e5;
         4'hdde8 	:	val_out <= 4'h20f5;
         4'hdde9 	:	val_out <= 4'h20f5;
         4'hddea 	:	val_out <= 4'h20f5;
         4'hddeb 	:	val_out <= 4'h20f5;
         4'hddf0 	:	val_out <= 4'h2106;
         4'hddf1 	:	val_out <= 4'h2106;
         4'hddf2 	:	val_out <= 4'h2106;
         4'hddf3 	:	val_out <= 4'h2106;
         4'hddf8 	:	val_out <= 4'h2117;
         4'hddf9 	:	val_out <= 4'h2117;
         4'hddfa 	:	val_out <= 4'h2117;
         4'hddfb 	:	val_out <= 4'h2117;
         4'hde00 	:	val_out <= 4'h2128;
         4'hde01 	:	val_out <= 4'h2128;
         4'hde02 	:	val_out <= 4'h2128;
         4'hde03 	:	val_out <= 4'h2128;
         4'hde08 	:	val_out <= 4'h2139;
         4'hde09 	:	val_out <= 4'h2139;
         4'hde0a 	:	val_out <= 4'h2139;
         4'hde0b 	:	val_out <= 4'h2139;
         4'hde10 	:	val_out <= 4'h214a;
         4'hde11 	:	val_out <= 4'h214a;
         4'hde12 	:	val_out <= 4'h214a;
         4'hde13 	:	val_out <= 4'h214a;
         4'hde18 	:	val_out <= 4'h215b;
         4'hde19 	:	val_out <= 4'h215b;
         4'hde1a 	:	val_out <= 4'h215b;
         4'hde1b 	:	val_out <= 4'h215b;
         4'hde20 	:	val_out <= 4'h216c;
         4'hde21 	:	val_out <= 4'h216c;
         4'hde22 	:	val_out <= 4'h216c;
         4'hde23 	:	val_out <= 4'h216c;
         4'hde28 	:	val_out <= 4'h217d;
         4'hde29 	:	val_out <= 4'h217d;
         4'hde2a 	:	val_out <= 4'h217d;
         4'hde2b 	:	val_out <= 4'h217d;
         4'hde30 	:	val_out <= 4'h218e;
         4'hde31 	:	val_out <= 4'h218e;
         4'hde32 	:	val_out <= 4'h218e;
         4'hde33 	:	val_out <= 4'h218e;
         4'hde38 	:	val_out <= 4'h219f;
         4'hde39 	:	val_out <= 4'h219f;
         4'hde3a 	:	val_out <= 4'h219f;
         4'hde3b 	:	val_out <= 4'h219f;
         4'hde40 	:	val_out <= 4'h21af;
         4'hde41 	:	val_out <= 4'h21af;
         4'hde42 	:	val_out <= 4'h21af;
         4'hde43 	:	val_out <= 4'h21af;
         4'hde48 	:	val_out <= 4'h21c0;
         4'hde49 	:	val_out <= 4'h21c0;
         4'hde4a 	:	val_out <= 4'h21c0;
         4'hde4b 	:	val_out <= 4'h21c0;
         4'hde50 	:	val_out <= 4'h21d2;
         4'hde51 	:	val_out <= 4'h21d2;
         4'hde52 	:	val_out <= 4'h21d2;
         4'hde53 	:	val_out <= 4'h21d2;
         4'hde58 	:	val_out <= 4'h21e3;
         4'hde59 	:	val_out <= 4'h21e3;
         4'hde5a 	:	val_out <= 4'h21e3;
         4'hde5b 	:	val_out <= 4'h21e3;
         4'hde60 	:	val_out <= 4'h21f4;
         4'hde61 	:	val_out <= 4'h21f4;
         4'hde62 	:	val_out <= 4'h21f4;
         4'hde63 	:	val_out <= 4'h21f4;
         4'hde68 	:	val_out <= 4'h2205;
         4'hde69 	:	val_out <= 4'h2205;
         4'hde6a 	:	val_out <= 4'h2205;
         4'hde6b 	:	val_out <= 4'h2205;
         4'hde70 	:	val_out <= 4'h2216;
         4'hde71 	:	val_out <= 4'h2216;
         4'hde72 	:	val_out <= 4'h2216;
         4'hde73 	:	val_out <= 4'h2216;
         4'hde78 	:	val_out <= 4'h2227;
         4'hde79 	:	val_out <= 4'h2227;
         4'hde7a 	:	val_out <= 4'h2227;
         4'hde7b 	:	val_out <= 4'h2227;
         4'hde80 	:	val_out <= 4'h2238;
         4'hde81 	:	val_out <= 4'h2238;
         4'hde82 	:	val_out <= 4'h2238;
         4'hde83 	:	val_out <= 4'h2238;
         4'hde88 	:	val_out <= 4'h2249;
         4'hde89 	:	val_out <= 4'h2249;
         4'hde8a 	:	val_out <= 4'h2249;
         4'hde8b 	:	val_out <= 4'h2249;
         4'hde90 	:	val_out <= 4'h225a;
         4'hde91 	:	val_out <= 4'h225a;
         4'hde92 	:	val_out <= 4'h225a;
         4'hde93 	:	val_out <= 4'h225a;
         4'hde98 	:	val_out <= 4'h226b;
         4'hde99 	:	val_out <= 4'h226b;
         4'hde9a 	:	val_out <= 4'h226b;
         4'hde9b 	:	val_out <= 4'h226b;
         4'hdea0 	:	val_out <= 4'h227c;
         4'hdea1 	:	val_out <= 4'h227c;
         4'hdea2 	:	val_out <= 4'h227c;
         4'hdea3 	:	val_out <= 4'h227c;
         4'hdea8 	:	val_out <= 4'h228e;
         4'hdea9 	:	val_out <= 4'h228e;
         4'hdeaa 	:	val_out <= 4'h228e;
         4'hdeab 	:	val_out <= 4'h228e;
         4'hdeb0 	:	val_out <= 4'h229f;
         4'hdeb1 	:	val_out <= 4'h229f;
         4'hdeb2 	:	val_out <= 4'h229f;
         4'hdeb3 	:	val_out <= 4'h229f;
         4'hdeb8 	:	val_out <= 4'h22b0;
         4'hdeb9 	:	val_out <= 4'h22b0;
         4'hdeba 	:	val_out <= 4'h22b0;
         4'hdebb 	:	val_out <= 4'h22b0;
         4'hdec0 	:	val_out <= 4'h22c1;
         4'hdec1 	:	val_out <= 4'h22c1;
         4'hdec2 	:	val_out <= 4'h22c1;
         4'hdec3 	:	val_out <= 4'h22c1;
         4'hdec8 	:	val_out <= 4'h22d2;
         4'hdec9 	:	val_out <= 4'h22d2;
         4'hdeca 	:	val_out <= 4'h22d2;
         4'hdecb 	:	val_out <= 4'h22d2;
         4'hded0 	:	val_out <= 4'h22e4;
         4'hded1 	:	val_out <= 4'h22e4;
         4'hded2 	:	val_out <= 4'h22e4;
         4'hded3 	:	val_out <= 4'h22e4;
         4'hded8 	:	val_out <= 4'h22f5;
         4'hded9 	:	val_out <= 4'h22f5;
         4'hdeda 	:	val_out <= 4'h22f5;
         4'hdedb 	:	val_out <= 4'h22f5;
         4'hdee0 	:	val_out <= 4'h2306;
         4'hdee1 	:	val_out <= 4'h2306;
         4'hdee2 	:	val_out <= 4'h2306;
         4'hdee3 	:	val_out <= 4'h2306;
         4'hdee8 	:	val_out <= 4'h2317;
         4'hdee9 	:	val_out <= 4'h2317;
         4'hdeea 	:	val_out <= 4'h2317;
         4'hdeeb 	:	val_out <= 4'h2317;
         4'hdef0 	:	val_out <= 4'h2329;
         4'hdef1 	:	val_out <= 4'h2329;
         4'hdef2 	:	val_out <= 4'h2329;
         4'hdef3 	:	val_out <= 4'h2329;
         4'hdef8 	:	val_out <= 4'h233a;
         4'hdef9 	:	val_out <= 4'h233a;
         4'hdefa 	:	val_out <= 4'h233a;
         4'hdefb 	:	val_out <= 4'h233a;
         4'hdf00 	:	val_out <= 4'h234b;
         4'hdf01 	:	val_out <= 4'h234b;
         4'hdf02 	:	val_out <= 4'h234b;
         4'hdf03 	:	val_out <= 4'h234b;
         4'hdf08 	:	val_out <= 4'h235d;
         4'hdf09 	:	val_out <= 4'h235d;
         4'hdf0a 	:	val_out <= 4'h235d;
         4'hdf0b 	:	val_out <= 4'h235d;
         4'hdf10 	:	val_out <= 4'h236e;
         4'hdf11 	:	val_out <= 4'h236e;
         4'hdf12 	:	val_out <= 4'h236e;
         4'hdf13 	:	val_out <= 4'h236e;
         4'hdf18 	:	val_out <= 4'h237f;
         4'hdf19 	:	val_out <= 4'h237f;
         4'hdf1a 	:	val_out <= 4'h237f;
         4'hdf1b 	:	val_out <= 4'h237f;
         4'hdf20 	:	val_out <= 4'h2391;
         4'hdf21 	:	val_out <= 4'h2391;
         4'hdf22 	:	val_out <= 4'h2391;
         4'hdf23 	:	val_out <= 4'h2391;
         4'hdf28 	:	val_out <= 4'h23a2;
         4'hdf29 	:	val_out <= 4'h23a2;
         4'hdf2a 	:	val_out <= 4'h23a2;
         4'hdf2b 	:	val_out <= 4'h23a2;
         4'hdf30 	:	val_out <= 4'h23b4;
         4'hdf31 	:	val_out <= 4'h23b4;
         4'hdf32 	:	val_out <= 4'h23b4;
         4'hdf33 	:	val_out <= 4'h23b4;
         4'hdf38 	:	val_out <= 4'h23c5;
         4'hdf39 	:	val_out <= 4'h23c5;
         4'hdf3a 	:	val_out <= 4'h23c5;
         4'hdf3b 	:	val_out <= 4'h23c5;
         4'hdf40 	:	val_out <= 4'h23d6;
         4'hdf41 	:	val_out <= 4'h23d6;
         4'hdf42 	:	val_out <= 4'h23d6;
         4'hdf43 	:	val_out <= 4'h23d6;
         4'hdf48 	:	val_out <= 4'h23e8;
         4'hdf49 	:	val_out <= 4'h23e8;
         4'hdf4a 	:	val_out <= 4'h23e8;
         4'hdf4b 	:	val_out <= 4'h23e8;
         4'hdf50 	:	val_out <= 4'h23f9;
         4'hdf51 	:	val_out <= 4'h23f9;
         4'hdf52 	:	val_out <= 4'h23f9;
         4'hdf53 	:	val_out <= 4'h23f9;
         4'hdf58 	:	val_out <= 4'h240b;
         4'hdf59 	:	val_out <= 4'h240b;
         4'hdf5a 	:	val_out <= 4'h240b;
         4'hdf5b 	:	val_out <= 4'h240b;
         4'hdf60 	:	val_out <= 4'h241c;
         4'hdf61 	:	val_out <= 4'h241c;
         4'hdf62 	:	val_out <= 4'h241c;
         4'hdf63 	:	val_out <= 4'h241c;
         4'hdf68 	:	val_out <= 4'h242e;
         4'hdf69 	:	val_out <= 4'h242e;
         4'hdf6a 	:	val_out <= 4'h242e;
         4'hdf6b 	:	val_out <= 4'h242e;
         4'hdf70 	:	val_out <= 4'h243f;
         4'hdf71 	:	val_out <= 4'h243f;
         4'hdf72 	:	val_out <= 4'h243f;
         4'hdf73 	:	val_out <= 4'h243f;
         4'hdf78 	:	val_out <= 4'h2451;
         4'hdf79 	:	val_out <= 4'h2451;
         4'hdf7a 	:	val_out <= 4'h2451;
         4'hdf7b 	:	val_out <= 4'h2451;
         4'hdf80 	:	val_out <= 4'h2462;
         4'hdf81 	:	val_out <= 4'h2462;
         4'hdf82 	:	val_out <= 4'h2462;
         4'hdf83 	:	val_out <= 4'h2462;
         4'hdf88 	:	val_out <= 4'h2474;
         4'hdf89 	:	val_out <= 4'h2474;
         4'hdf8a 	:	val_out <= 4'h2474;
         4'hdf8b 	:	val_out <= 4'h2474;
         4'hdf90 	:	val_out <= 4'h2486;
         4'hdf91 	:	val_out <= 4'h2486;
         4'hdf92 	:	val_out <= 4'h2486;
         4'hdf93 	:	val_out <= 4'h2486;
         4'hdf98 	:	val_out <= 4'h2497;
         4'hdf99 	:	val_out <= 4'h2497;
         4'hdf9a 	:	val_out <= 4'h2497;
         4'hdf9b 	:	val_out <= 4'h2497;
         4'hdfa0 	:	val_out <= 4'h24a9;
         4'hdfa1 	:	val_out <= 4'h24a9;
         4'hdfa2 	:	val_out <= 4'h24a9;
         4'hdfa3 	:	val_out <= 4'h24a9;
         4'hdfa8 	:	val_out <= 4'h24ba;
         4'hdfa9 	:	val_out <= 4'h24ba;
         4'hdfaa 	:	val_out <= 4'h24ba;
         4'hdfab 	:	val_out <= 4'h24ba;
         4'hdfb0 	:	val_out <= 4'h24cc;
         4'hdfb1 	:	val_out <= 4'h24cc;
         4'hdfb2 	:	val_out <= 4'h24cc;
         4'hdfb3 	:	val_out <= 4'h24cc;
         4'hdfb8 	:	val_out <= 4'h24de;
         4'hdfb9 	:	val_out <= 4'h24de;
         4'hdfba 	:	val_out <= 4'h24de;
         4'hdfbb 	:	val_out <= 4'h24de;
         4'hdfc0 	:	val_out <= 4'h24ef;
         4'hdfc1 	:	val_out <= 4'h24ef;
         4'hdfc2 	:	val_out <= 4'h24ef;
         4'hdfc3 	:	val_out <= 4'h24ef;
         4'hdfc8 	:	val_out <= 4'h2501;
         4'hdfc9 	:	val_out <= 4'h2501;
         4'hdfca 	:	val_out <= 4'h2501;
         4'hdfcb 	:	val_out <= 4'h2501;
         4'hdfd0 	:	val_out <= 4'h2513;
         4'hdfd1 	:	val_out <= 4'h2513;
         4'hdfd2 	:	val_out <= 4'h2513;
         4'hdfd3 	:	val_out <= 4'h2513;
         4'hdfd8 	:	val_out <= 4'h2524;
         4'hdfd9 	:	val_out <= 4'h2524;
         4'hdfda 	:	val_out <= 4'h2524;
         4'hdfdb 	:	val_out <= 4'h2524;
         4'hdfe0 	:	val_out <= 4'h2536;
         4'hdfe1 	:	val_out <= 4'h2536;
         4'hdfe2 	:	val_out <= 4'h2536;
         4'hdfe3 	:	val_out <= 4'h2536;
         4'hdfe8 	:	val_out <= 4'h2548;
         4'hdfe9 	:	val_out <= 4'h2548;
         4'hdfea 	:	val_out <= 4'h2548;
         4'hdfeb 	:	val_out <= 4'h2548;
         4'hdff0 	:	val_out <= 4'h255a;
         4'hdff1 	:	val_out <= 4'h255a;
         4'hdff2 	:	val_out <= 4'h255a;
         4'hdff3 	:	val_out <= 4'h255a;
         4'hdff8 	:	val_out <= 4'h256b;
         4'hdff9 	:	val_out <= 4'h256b;
         4'hdffa 	:	val_out <= 4'h256b;
         4'hdffb 	:	val_out <= 4'h256b;
         4'he000 	:	val_out <= 4'h257d;
         4'he001 	:	val_out <= 4'h257d;
         4'he002 	:	val_out <= 4'h257d;
         4'he003 	:	val_out <= 4'h257d;
         4'he008 	:	val_out <= 4'h258f;
         4'he009 	:	val_out <= 4'h258f;
         4'he00a 	:	val_out <= 4'h258f;
         4'he00b 	:	val_out <= 4'h258f;
         4'he010 	:	val_out <= 4'h25a1;
         4'he011 	:	val_out <= 4'h25a1;
         4'he012 	:	val_out <= 4'h25a1;
         4'he013 	:	val_out <= 4'h25a1;
         4'he018 	:	val_out <= 4'h25b2;
         4'he019 	:	val_out <= 4'h25b2;
         4'he01a 	:	val_out <= 4'h25b2;
         4'he01b 	:	val_out <= 4'h25b2;
         4'he020 	:	val_out <= 4'h25c4;
         4'he021 	:	val_out <= 4'h25c4;
         4'he022 	:	val_out <= 4'h25c4;
         4'he023 	:	val_out <= 4'h25c4;
         4'he028 	:	val_out <= 4'h25d6;
         4'he029 	:	val_out <= 4'h25d6;
         4'he02a 	:	val_out <= 4'h25d6;
         4'he02b 	:	val_out <= 4'h25d6;
         4'he030 	:	val_out <= 4'h25e8;
         4'he031 	:	val_out <= 4'h25e8;
         4'he032 	:	val_out <= 4'h25e8;
         4'he033 	:	val_out <= 4'h25e8;
         4'he038 	:	val_out <= 4'h25fa;
         4'he039 	:	val_out <= 4'h25fa;
         4'he03a 	:	val_out <= 4'h25fa;
         4'he03b 	:	val_out <= 4'h25fa;
         4'he040 	:	val_out <= 4'h260c;
         4'he041 	:	val_out <= 4'h260c;
         4'he042 	:	val_out <= 4'h260c;
         4'he043 	:	val_out <= 4'h260c;
         4'he048 	:	val_out <= 4'h261e;
         4'he049 	:	val_out <= 4'h261e;
         4'he04a 	:	val_out <= 4'h261e;
         4'he04b 	:	val_out <= 4'h261e;
         4'he050 	:	val_out <= 4'h262f;
         4'he051 	:	val_out <= 4'h262f;
         4'he052 	:	val_out <= 4'h262f;
         4'he053 	:	val_out <= 4'h262f;
         4'he058 	:	val_out <= 4'h2641;
         4'he059 	:	val_out <= 4'h2641;
         4'he05a 	:	val_out <= 4'h2641;
         4'he05b 	:	val_out <= 4'h2641;
         4'he060 	:	val_out <= 4'h2653;
         4'he061 	:	val_out <= 4'h2653;
         4'he062 	:	val_out <= 4'h2653;
         4'he063 	:	val_out <= 4'h2653;
         4'he068 	:	val_out <= 4'h2665;
         4'he069 	:	val_out <= 4'h2665;
         4'he06a 	:	val_out <= 4'h2665;
         4'he06b 	:	val_out <= 4'h2665;
         4'he070 	:	val_out <= 4'h2677;
         4'he071 	:	val_out <= 4'h2677;
         4'he072 	:	val_out <= 4'h2677;
         4'he073 	:	val_out <= 4'h2677;
         4'he078 	:	val_out <= 4'h2689;
         4'he079 	:	val_out <= 4'h2689;
         4'he07a 	:	val_out <= 4'h2689;
         4'he07b 	:	val_out <= 4'h2689;
         4'he080 	:	val_out <= 4'h269b;
         4'he081 	:	val_out <= 4'h269b;
         4'he082 	:	val_out <= 4'h269b;
         4'he083 	:	val_out <= 4'h269b;
         4'he088 	:	val_out <= 4'h26ad;
         4'he089 	:	val_out <= 4'h26ad;
         4'he08a 	:	val_out <= 4'h26ad;
         4'he08b 	:	val_out <= 4'h26ad;
         4'he090 	:	val_out <= 4'h26bf;
         4'he091 	:	val_out <= 4'h26bf;
         4'he092 	:	val_out <= 4'h26bf;
         4'he093 	:	val_out <= 4'h26bf;
         4'he098 	:	val_out <= 4'h26d1;
         4'he099 	:	val_out <= 4'h26d1;
         4'he09a 	:	val_out <= 4'h26d1;
         4'he09b 	:	val_out <= 4'h26d1;
         4'he0a0 	:	val_out <= 4'h26e3;
         4'he0a1 	:	val_out <= 4'h26e3;
         4'he0a2 	:	val_out <= 4'h26e3;
         4'he0a3 	:	val_out <= 4'h26e3;
         4'he0a8 	:	val_out <= 4'h26f5;
         4'he0a9 	:	val_out <= 4'h26f5;
         4'he0aa 	:	val_out <= 4'h26f5;
         4'he0ab 	:	val_out <= 4'h26f5;
         4'he0b0 	:	val_out <= 4'h2707;
         4'he0b1 	:	val_out <= 4'h2707;
         4'he0b2 	:	val_out <= 4'h2707;
         4'he0b3 	:	val_out <= 4'h2707;
         4'he0b8 	:	val_out <= 4'h2719;
         4'he0b9 	:	val_out <= 4'h2719;
         4'he0ba 	:	val_out <= 4'h2719;
         4'he0bb 	:	val_out <= 4'h2719;
         4'he0c0 	:	val_out <= 4'h272b;
         4'he0c1 	:	val_out <= 4'h272b;
         4'he0c2 	:	val_out <= 4'h272b;
         4'he0c3 	:	val_out <= 4'h272b;
         4'he0c8 	:	val_out <= 4'h273e;
         4'he0c9 	:	val_out <= 4'h273e;
         4'he0ca 	:	val_out <= 4'h273e;
         4'he0cb 	:	val_out <= 4'h273e;
         4'he0d0 	:	val_out <= 4'h2750;
         4'he0d1 	:	val_out <= 4'h2750;
         4'he0d2 	:	val_out <= 4'h2750;
         4'he0d3 	:	val_out <= 4'h2750;
         4'he0d8 	:	val_out <= 4'h2762;
         4'he0d9 	:	val_out <= 4'h2762;
         4'he0da 	:	val_out <= 4'h2762;
         4'he0db 	:	val_out <= 4'h2762;
         4'he0e0 	:	val_out <= 4'h2774;
         4'he0e1 	:	val_out <= 4'h2774;
         4'he0e2 	:	val_out <= 4'h2774;
         4'he0e3 	:	val_out <= 4'h2774;
         4'he0e8 	:	val_out <= 4'h2786;
         4'he0e9 	:	val_out <= 4'h2786;
         4'he0ea 	:	val_out <= 4'h2786;
         4'he0eb 	:	val_out <= 4'h2786;
         4'he0f0 	:	val_out <= 4'h2798;
         4'he0f1 	:	val_out <= 4'h2798;
         4'he0f2 	:	val_out <= 4'h2798;
         4'he0f3 	:	val_out <= 4'h2798;
         4'he0f8 	:	val_out <= 4'h27aa;
         4'he0f9 	:	val_out <= 4'h27aa;
         4'he0fa 	:	val_out <= 4'h27aa;
         4'he0fb 	:	val_out <= 4'h27aa;
         4'he100 	:	val_out <= 4'h27bd;
         4'he101 	:	val_out <= 4'h27bd;
         4'he102 	:	val_out <= 4'h27bd;
         4'he103 	:	val_out <= 4'h27bd;
         4'he108 	:	val_out <= 4'h27cf;
         4'he109 	:	val_out <= 4'h27cf;
         4'he10a 	:	val_out <= 4'h27cf;
         4'he10b 	:	val_out <= 4'h27cf;
         4'he110 	:	val_out <= 4'h27e1;
         4'he111 	:	val_out <= 4'h27e1;
         4'he112 	:	val_out <= 4'h27e1;
         4'he113 	:	val_out <= 4'h27e1;
         4'he118 	:	val_out <= 4'h27f3;
         4'he119 	:	val_out <= 4'h27f3;
         4'he11a 	:	val_out <= 4'h27f3;
         4'he11b 	:	val_out <= 4'h27f3;
         4'he120 	:	val_out <= 4'h2806;
         4'he121 	:	val_out <= 4'h2806;
         4'he122 	:	val_out <= 4'h2806;
         4'he123 	:	val_out <= 4'h2806;
         4'he128 	:	val_out <= 4'h2818;
         4'he129 	:	val_out <= 4'h2818;
         4'he12a 	:	val_out <= 4'h2818;
         4'he12b 	:	val_out <= 4'h2818;
         4'he130 	:	val_out <= 4'h282a;
         4'he131 	:	val_out <= 4'h282a;
         4'he132 	:	val_out <= 4'h282a;
         4'he133 	:	val_out <= 4'h282a;
         4'he138 	:	val_out <= 4'h283c;
         4'he139 	:	val_out <= 4'h283c;
         4'he13a 	:	val_out <= 4'h283c;
         4'he13b 	:	val_out <= 4'h283c;
         4'he140 	:	val_out <= 4'h284f;
         4'he141 	:	val_out <= 4'h284f;
         4'he142 	:	val_out <= 4'h284f;
         4'he143 	:	val_out <= 4'h284f;
         4'he148 	:	val_out <= 4'h2861;
         4'he149 	:	val_out <= 4'h2861;
         4'he14a 	:	val_out <= 4'h2861;
         4'he14b 	:	val_out <= 4'h2861;
         4'he150 	:	val_out <= 4'h2873;
         4'he151 	:	val_out <= 4'h2873;
         4'he152 	:	val_out <= 4'h2873;
         4'he153 	:	val_out <= 4'h2873;
         4'he158 	:	val_out <= 4'h2886;
         4'he159 	:	val_out <= 4'h2886;
         4'he15a 	:	val_out <= 4'h2886;
         4'he15b 	:	val_out <= 4'h2886;
         4'he160 	:	val_out <= 4'h2898;
         4'he161 	:	val_out <= 4'h2898;
         4'he162 	:	val_out <= 4'h2898;
         4'he163 	:	val_out <= 4'h2898;
         4'he168 	:	val_out <= 4'h28aa;
         4'he169 	:	val_out <= 4'h28aa;
         4'he16a 	:	val_out <= 4'h28aa;
         4'he16b 	:	val_out <= 4'h28aa;
         4'he170 	:	val_out <= 4'h28bd;
         4'he171 	:	val_out <= 4'h28bd;
         4'he172 	:	val_out <= 4'h28bd;
         4'he173 	:	val_out <= 4'h28bd;
         4'he178 	:	val_out <= 4'h28cf;
         4'he179 	:	val_out <= 4'h28cf;
         4'he17a 	:	val_out <= 4'h28cf;
         4'he17b 	:	val_out <= 4'h28cf;
         4'he180 	:	val_out <= 4'h28e2;
         4'he181 	:	val_out <= 4'h28e2;
         4'he182 	:	val_out <= 4'h28e2;
         4'he183 	:	val_out <= 4'h28e2;
         4'he188 	:	val_out <= 4'h28f4;
         4'he189 	:	val_out <= 4'h28f4;
         4'he18a 	:	val_out <= 4'h28f4;
         4'he18b 	:	val_out <= 4'h28f4;
         4'he190 	:	val_out <= 4'h2906;
         4'he191 	:	val_out <= 4'h2906;
         4'he192 	:	val_out <= 4'h2906;
         4'he193 	:	val_out <= 4'h2906;
         4'he198 	:	val_out <= 4'h2919;
         4'he199 	:	val_out <= 4'h2919;
         4'he19a 	:	val_out <= 4'h2919;
         4'he19b 	:	val_out <= 4'h2919;
         4'he1a0 	:	val_out <= 4'h292b;
         4'he1a1 	:	val_out <= 4'h292b;
         4'he1a2 	:	val_out <= 4'h292b;
         4'he1a3 	:	val_out <= 4'h292b;
         4'he1a8 	:	val_out <= 4'h293e;
         4'he1a9 	:	val_out <= 4'h293e;
         4'he1aa 	:	val_out <= 4'h293e;
         4'he1ab 	:	val_out <= 4'h293e;
         4'he1b0 	:	val_out <= 4'h2950;
         4'he1b1 	:	val_out <= 4'h2950;
         4'he1b2 	:	val_out <= 4'h2950;
         4'he1b3 	:	val_out <= 4'h2950;
         4'he1b8 	:	val_out <= 4'h2963;
         4'he1b9 	:	val_out <= 4'h2963;
         4'he1ba 	:	val_out <= 4'h2963;
         4'he1bb 	:	val_out <= 4'h2963;
         4'he1c0 	:	val_out <= 4'h2975;
         4'he1c1 	:	val_out <= 4'h2975;
         4'he1c2 	:	val_out <= 4'h2975;
         4'he1c3 	:	val_out <= 4'h2975;
         4'he1c8 	:	val_out <= 4'h2988;
         4'he1c9 	:	val_out <= 4'h2988;
         4'he1ca 	:	val_out <= 4'h2988;
         4'he1cb 	:	val_out <= 4'h2988;
         4'he1d0 	:	val_out <= 4'h299a;
         4'he1d1 	:	val_out <= 4'h299a;
         4'he1d2 	:	val_out <= 4'h299a;
         4'he1d3 	:	val_out <= 4'h299a;
         4'he1d8 	:	val_out <= 4'h29ad;
         4'he1d9 	:	val_out <= 4'h29ad;
         4'he1da 	:	val_out <= 4'h29ad;
         4'he1db 	:	val_out <= 4'h29ad;
         4'he1e0 	:	val_out <= 4'h29bf;
         4'he1e1 	:	val_out <= 4'h29bf;
         4'he1e2 	:	val_out <= 4'h29bf;
         4'he1e3 	:	val_out <= 4'h29bf;
         4'he1e8 	:	val_out <= 4'h29d2;
         4'he1e9 	:	val_out <= 4'h29d2;
         4'he1ea 	:	val_out <= 4'h29d2;
         4'he1eb 	:	val_out <= 4'h29d2;
         4'he1f0 	:	val_out <= 4'h29e5;
         4'he1f1 	:	val_out <= 4'h29e5;
         4'he1f2 	:	val_out <= 4'h29e5;
         4'he1f3 	:	val_out <= 4'h29e5;
         4'he1f8 	:	val_out <= 4'h29f7;
         4'he1f9 	:	val_out <= 4'h29f7;
         4'he1fa 	:	val_out <= 4'h29f7;
         4'he1fb 	:	val_out <= 4'h29f7;
         4'he200 	:	val_out <= 4'h2a0a;
         4'he201 	:	val_out <= 4'h2a0a;
         4'he202 	:	val_out <= 4'h2a0a;
         4'he203 	:	val_out <= 4'h2a0a;
         4'he208 	:	val_out <= 4'h2a1c;
         4'he209 	:	val_out <= 4'h2a1c;
         4'he20a 	:	val_out <= 4'h2a1c;
         4'he20b 	:	val_out <= 4'h2a1c;
         4'he210 	:	val_out <= 4'h2a2f;
         4'he211 	:	val_out <= 4'h2a2f;
         4'he212 	:	val_out <= 4'h2a2f;
         4'he213 	:	val_out <= 4'h2a2f;
         4'he218 	:	val_out <= 4'h2a42;
         4'he219 	:	val_out <= 4'h2a42;
         4'he21a 	:	val_out <= 4'h2a42;
         4'he21b 	:	val_out <= 4'h2a42;
         4'he220 	:	val_out <= 4'h2a54;
         4'he221 	:	val_out <= 4'h2a54;
         4'he222 	:	val_out <= 4'h2a54;
         4'he223 	:	val_out <= 4'h2a54;
         4'he228 	:	val_out <= 4'h2a67;
         4'he229 	:	val_out <= 4'h2a67;
         4'he22a 	:	val_out <= 4'h2a67;
         4'he22b 	:	val_out <= 4'h2a67;
         4'he230 	:	val_out <= 4'h2a7a;
         4'he231 	:	val_out <= 4'h2a7a;
         4'he232 	:	val_out <= 4'h2a7a;
         4'he233 	:	val_out <= 4'h2a7a;
         4'he238 	:	val_out <= 4'h2a8d;
         4'he239 	:	val_out <= 4'h2a8d;
         4'he23a 	:	val_out <= 4'h2a8d;
         4'he23b 	:	val_out <= 4'h2a8d;
         4'he240 	:	val_out <= 4'h2a9f;
         4'he241 	:	val_out <= 4'h2a9f;
         4'he242 	:	val_out <= 4'h2a9f;
         4'he243 	:	val_out <= 4'h2a9f;
         4'he248 	:	val_out <= 4'h2ab2;
         4'he249 	:	val_out <= 4'h2ab2;
         4'he24a 	:	val_out <= 4'h2ab2;
         4'he24b 	:	val_out <= 4'h2ab2;
         4'he250 	:	val_out <= 4'h2ac5;
         4'he251 	:	val_out <= 4'h2ac5;
         4'he252 	:	val_out <= 4'h2ac5;
         4'he253 	:	val_out <= 4'h2ac5;
         4'he258 	:	val_out <= 4'h2ad7;
         4'he259 	:	val_out <= 4'h2ad7;
         4'he25a 	:	val_out <= 4'h2ad7;
         4'he25b 	:	val_out <= 4'h2ad7;
         4'he260 	:	val_out <= 4'h2aea;
         4'he261 	:	val_out <= 4'h2aea;
         4'he262 	:	val_out <= 4'h2aea;
         4'he263 	:	val_out <= 4'h2aea;
         4'he268 	:	val_out <= 4'h2afd;
         4'he269 	:	val_out <= 4'h2afd;
         4'he26a 	:	val_out <= 4'h2afd;
         4'he26b 	:	val_out <= 4'h2afd;
         4'he270 	:	val_out <= 4'h2b10;
         4'he271 	:	val_out <= 4'h2b10;
         4'he272 	:	val_out <= 4'h2b10;
         4'he273 	:	val_out <= 4'h2b10;
         4'he278 	:	val_out <= 4'h2b23;
         4'he279 	:	val_out <= 4'h2b23;
         4'he27a 	:	val_out <= 4'h2b23;
         4'he27b 	:	val_out <= 4'h2b23;
         4'he280 	:	val_out <= 4'h2b35;
         4'he281 	:	val_out <= 4'h2b35;
         4'he282 	:	val_out <= 4'h2b35;
         4'he283 	:	val_out <= 4'h2b35;
         4'he288 	:	val_out <= 4'h2b48;
         4'he289 	:	val_out <= 4'h2b48;
         4'he28a 	:	val_out <= 4'h2b48;
         4'he28b 	:	val_out <= 4'h2b48;
         4'he290 	:	val_out <= 4'h2b5b;
         4'he291 	:	val_out <= 4'h2b5b;
         4'he292 	:	val_out <= 4'h2b5b;
         4'he293 	:	val_out <= 4'h2b5b;
         4'he298 	:	val_out <= 4'h2b6e;
         4'he299 	:	val_out <= 4'h2b6e;
         4'he29a 	:	val_out <= 4'h2b6e;
         4'he29b 	:	val_out <= 4'h2b6e;
         4'he2a0 	:	val_out <= 4'h2b81;
         4'he2a1 	:	val_out <= 4'h2b81;
         4'he2a2 	:	val_out <= 4'h2b81;
         4'he2a3 	:	val_out <= 4'h2b81;
         4'he2a8 	:	val_out <= 4'h2b94;
         4'he2a9 	:	val_out <= 4'h2b94;
         4'he2aa 	:	val_out <= 4'h2b94;
         4'he2ab 	:	val_out <= 4'h2b94;
         4'he2b0 	:	val_out <= 4'h2ba7;
         4'he2b1 	:	val_out <= 4'h2ba7;
         4'he2b2 	:	val_out <= 4'h2ba7;
         4'he2b3 	:	val_out <= 4'h2ba7;
         4'he2b8 	:	val_out <= 4'h2bba;
         4'he2b9 	:	val_out <= 4'h2bba;
         4'he2ba 	:	val_out <= 4'h2bba;
         4'he2bb 	:	val_out <= 4'h2bba;
         4'he2c0 	:	val_out <= 4'h2bcc;
         4'he2c1 	:	val_out <= 4'h2bcc;
         4'he2c2 	:	val_out <= 4'h2bcc;
         4'he2c3 	:	val_out <= 4'h2bcc;
         4'he2c8 	:	val_out <= 4'h2bdf;
         4'he2c9 	:	val_out <= 4'h2bdf;
         4'he2ca 	:	val_out <= 4'h2bdf;
         4'he2cb 	:	val_out <= 4'h2bdf;
         4'he2d0 	:	val_out <= 4'h2bf2;
         4'he2d1 	:	val_out <= 4'h2bf2;
         4'he2d2 	:	val_out <= 4'h2bf2;
         4'he2d3 	:	val_out <= 4'h2bf2;
         4'he2d8 	:	val_out <= 4'h2c05;
         4'he2d9 	:	val_out <= 4'h2c05;
         4'he2da 	:	val_out <= 4'h2c05;
         4'he2db 	:	val_out <= 4'h2c05;
         4'he2e0 	:	val_out <= 4'h2c18;
         4'he2e1 	:	val_out <= 4'h2c18;
         4'he2e2 	:	val_out <= 4'h2c18;
         4'he2e3 	:	val_out <= 4'h2c18;
         4'he2e8 	:	val_out <= 4'h2c2b;
         4'he2e9 	:	val_out <= 4'h2c2b;
         4'he2ea 	:	val_out <= 4'h2c2b;
         4'he2eb 	:	val_out <= 4'h2c2b;
         4'he2f0 	:	val_out <= 4'h2c3e;
         4'he2f1 	:	val_out <= 4'h2c3e;
         4'he2f2 	:	val_out <= 4'h2c3e;
         4'he2f3 	:	val_out <= 4'h2c3e;
         4'he2f8 	:	val_out <= 4'h2c51;
         4'he2f9 	:	val_out <= 4'h2c51;
         4'he2fa 	:	val_out <= 4'h2c51;
         4'he2fb 	:	val_out <= 4'h2c51;
         4'he300 	:	val_out <= 4'h2c64;
         4'he301 	:	val_out <= 4'h2c64;
         4'he302 	:	val_out <= 4'h2c64;
         4'he303 	:	val_out <= 4'h2c64;
         4'he308 	:	val_out <= 4'h2c77;
         4'he309 	:	val_out <= 4'h2c77;
         4'he30a 	:	val_out <= 4'h2c77;
         4'he30b 	:	val_out <= 4'h2c77;
         4'he310 	:	val_out <= 4'h2c8a;
         4'he311 	:	val_out <= 4'h2c8a;
         4'he312 	:	val_out <= 4'h2c8a;
         4'he313 	:	val_out <= 4'h2c8a;
         4'he318 	:	val_out <= 4'h2c9d;
         4'he319 	:	val_out <= 4'h2c9d;
         4'he31a 	:	val_out <= 4'h2c9d;
         4'he31b 	:	val_out <= 4'h2c9d;
         4'he320 	:	val_out <= 4'h2cb1;
         4'he321 	:	val_out <= 4'h2cb1;
         4'he322 	:	val_out <= 4'h2cb1;
         4'he323 	:	val_out <= 4'h2cb1;
         4'he328 	:	val_out <= 4'h2cc4;
         4'he329 	:	val_out <= 4'h2cc4;
         4'he32a 	:	val_out <= 4'h2cc4;
         4'he32b 	:	val_out <= 4'h2cc4;
         4'he330 	:	val_out <= 4'h2cd7;
         4'he331 	:	val_out <= 4'h2cd7;
         4'he332 	:	val_out <= 4'h2cd7;
         4'he333 	:	val_out <= 4'h2cd7;
         4'he338 	:	val_out <= 4'h2cea;
         4'he339 	:	val_out <= 4'h2cea;
         4'he33a 	:	val_out <= 4'h2cea;
         4'he33b 	:	val_out <= 4'h2cea;
         4'he340 	:	val_out <= 4'h2cfd;
         4'he341 	:	val_out <= 4'h2cfd;
         4'he342 	:	val_out <= 4'h2cfd;
         4'he343 	:	val_out <= 4'h2cfd;
         4'he348 	:	val_out <= 4'h2d10;
         4'he349 	:	val_out <= 4'h2d10;
         4'he34a 	:	val_out <= 4'h2d10;
         4'he34b 	:	val_out <= 4'h2d10;
         4'he350 	:	val_out <= 4'h2d23;
         4'he351 	:	val_out <= 4'h2d23;
         4'he352 	:	val_out <= 4'h2d23;
         4'he353 	:	val_out <= 4'h2d23;
         4'he358 	:	val_out <= 4'h2d36;
         4'he359 	:	val_out <= 4'h2d36;
         4'he35a 	:	val_out <= 4'h2d36;
         4'he35b 	:	val_out <= 4'h2d36;
         4'he360 	:	val_out <= 4'h2d4a;
         4'he361 	:	val_out <= 4'h2d4a;
         4'he362 	:	val_out <= 4'h2d4a;
         4'he363 	:	val_out <= 4'h2d4a;
         4'he368 	:	val_out <= 4'h2d5d;
         4'he369 	:	val_out <= 4'h2d5d;
         4'he36a 	:	val_out <= 4'h2d5d;
         4'he36b 	:	val_out <= 4'h2d5d;
         4'he370 	:	val_out <= 4'h2d70;
         4'he371 	:	val_out <= 4'h2d70;
         4'he372 	:	val_out <= 4'h2d70;
         4'he373 	:	val_out <= 4'h2d70;
         4'he378 	:	val_out <= 4'h2d83;
         4'he379 	:	val_out <= 4'h2d83;
         4'he37a 	:	val_out <= 4'h2d83;
         4'he37b 	:	val_out <= 4'h2d83;
         4'he380 	:	val_out <= 4'h2d96;
         4'he381 	:	val_out <= 4'h2d96;
         4'he382 	:	val_out <= 4'h2d96;
         4'he383 	:	val_out <= 4'h2d96;
         4'he388 	:	val_out <= 4'h2daa;
         4'he389 	:	val_out <= 4'h2daa;
         4'he38a 	:	val_out <= 4'h2daa;
         4'he38b 	:	val_out <= 4'h2daa;
         4'he390 	:	val_out <= 4'h2dbd;
         4'he391 	:	val_out <= 4'h2dbd;
         4'he392 	:	val_out <= 4'h2dbd;
         4'he393 	:	val_out <= 4'h2dbd;
         4'he398 	:	val_out <= 4'h2dd0;
         4'he399 	:	val_out <= 4'h2dd0;
         4'he39a 	:	val_out <= 4'h2dd0;
         4'he39b 	:	val_out <= 4'h2dd0;
         4'he3a0 	:	val_out <= 4'h2de3;
         4'he3a1 	:	val_out <= 4'h2de3;
         4'he3a2 	:	val_out <= 4'h2de3;
         4'he3a3 	:	val_out <= 4'h2de3;
         4'he3a8 	:	val_out <= 4'h2df7;
         4'he3a9 	:	val_out <= 4'h2df7;
         4'he3aa 	:	val_out <= 4'h2df7;
         4'he3ab 	:	val_out <= 4'h2df7;
         4'he3b0 	:	val_out <= 4'h2e0a;
         4'he3b1 	:	val_out <= 4'h2e0a;
         4'he3b2 	:	val_out <= 4'h2e0a;
         4'he3b3 	:	val_out <= 4'h2e0a;
         4'he3b8 	:	val_out <= 4'h2e1d;
         4'he3b9 	:	val_out <= 4'h2e1d;
         4'he3ba 	:	val_out <= 4'h2e1d;
         4'he3bb 	:	val_out <= 4'h2e1d;
         4'he3c0 	:	val_out <= 4'h2e31;
         4'he3c1 	:	val_out <= 4'h2e31;
         4'he3c2 	:	val_out <= 4'h2e31;
         4'he3c3 	:	val_out <= 4'h2e31;
         4'he3c8 	:	val_out <= 4'h2e44;
         4'he3c9 	:	val_out <= 4'h2e44;
         4'he3ca 	:	val_out <= 4'h2e44;
         4'he3cb 	:	val_out <= 4'h2e44;
         4'he3d0 	:	val_out <= 4'h2e57;
         4'he3d1 	:	val_out <= 4'h2e57;
         4'he3d2 	:	val_out <= 4'h2e57;
         4'he3d3 	:	val_out <= 4'h2e57;
         4'he3d8 	:	val_out <= 4'h2e6b;
         4'he3d9 	:	val_out <= 4'h2e6b;
         4'he3da 	:	val_out <= 4'h2e6b;
         4'he3db 	:	val_out <= 4'h2e6b;
         4'he3e0 	:	val_out <= 4'h2e7e;
         4'he3e1 	:	val_out <= 4'h2e7e;
         4'he3e2 	:	val_out <= 4'h2e7e;
         4'he3e3 	:	val_out <= 4'h2e7e;
         4'he3e8 	:	val_out <= 4'h2e91;
         4'he3e9 	:	val_out <= 4'h2e91;
         4'he3ea 	:	val_out <= 4'h2e91;
         4'he3eb 	:	val_out <= 4'h2e91;
         4'he3f0 	:	val_out <= 4'h2ea5;
         4'he3f1 	:	val_out <= 4'h2ea5;
         4'he3f2 	:	val_out <= 4'h2ea5;
         4'he3f3 	:	val_out <= 4'h2ea5;
         4'he3f8 	:	val_out <= 4'h2eb8;
         4'he3f9 	:	val_out <= 4'h2eb8;
         4'he3fa 	:	val_out <= 4'h2eb8;
         4'he3fb 	:	val_out <= 4'h2eb8;
         4'he400 	:	val_out <= 4'h2ecc;
         4'he401 	:	val_out <= 4'h2ecc;
         4'he402 	:	val_out <= 4'h2ecc;
         4'he403 	:	val_out <= 4'h2ecc;
         4'he408 	:	val_out <= 4'h2edf;
         4'he409 	:	val_out <= 4'h2edf;
         4'he40a 	:	val_out <= 4'h2edf;
         4'he40b 	:	val_out <= 4'h2edf;
         4'he410 	:	val_out <= 4'h2ef3;
         4'he411 	:	val_out <= 4'h2ef3;
         4'he412 	:	val_out <= 4'h2ef3;
         4'he413 	:	val_out <= 4'h2ef3;
         4'he418 	:	val_out <= 4'h2f06;
         4'he419 	:	val_out <= 4'h2f06;
         4'he41a 	:	val_out <= 4'h2f06;
         4'he41b 	:	val_out <= 4'h2f06;
         4'he420 	:	val_out <= 4'h2f1a;
         4'he421 	:	val_out <= 4'h2f1a;
         4'he422 	:	val_out <= 4'h2f1a;
         4'he423 	:	val_out <= 4'h2f1a;
         4'he428 	:	val_out <= 4'h2f2d;
         4'he429 	:	val_out <= 4'h2f2d;
         4'he42a 	:	val_out <= 4'h2f2d;
         4'he42b 	:	val_out <= 4'h2f2d;
         4'he430 	:	val_out <= 4'h2f40;
         4'he431 	:	val_out <= 4'h2f40;
         4'he432 	:	val_out <= 4'h2f40;
         4'he433 	:	val_out <= 4'h2f40;
         4'he438 	:	val_out <= 4'h2f54;
         4'he439 	:	val_out <= 4'h2f54;
         4'he43a 	:	val_out <= 4'h2f54;
         4'he43b 	:	val_out <= 4'h2f54;
         4'he440 	:	val_out <= 4'h2f68;
         4'he441 	:	val_out <= 4'h2f68;
         4'he442 	:	val_out <= 4'h2f68;
         4'he443 	:	val_out <= 4'h2f68;
         4'he448 	:	val_out <= 4'h2f7b;
         4'he449 	:	val_out <= 4'h2f7b;
         4'he44a 	:	val_out <= 4'h2f7b;
         4'he44b 	:	val_out <= 4'h2f7b;
         4'he450 	:	val_out <= 4'h2f8f;
         4'he451 	:	val_out <= 4'h2f8f;
         4'he452 	:	val_out <= 4'h2f8f;
         4'he453 	:	val_out <= 4'h2f8f;
         4'he458 	:	val_out <= 4'h2fa2;
         4'he459 	:	val_out <= 4'h2fa2;
         4'he45a 	:	val_out <= 4'h2fa2;
         4'he45b 	:	val_out <= 4'h2fa2;
         4'he460 	:	val_out <= 4'h2fb6;
         4'he461 	:	val_out <= 4'h2fb6;
         4'he462 	:	val_out <= 4'h2fb6;
         4'he463 	:	val_out <= 4'h2fb6;
         4'he468 	:	val_out <= 4'h2fc9;
         4'he469 	:	val_out <= 4'h2fc9;
         4'he46a 	:	val_out <= 4'h2fc9;
         4'he46b 	:	val_out <= 4'h2fc9;
         4'he470 	:	val_out <= 4'h2fdd;
         4'he471 	:	val_out <= 4'h2fdd;
         4'he472 	:	val_out <= 4'h2fdd;
         4'he473 	:	val_out <= 4'h2fdd;
         4'he478 	:	val_out <= 4'h2ff0;
         4'he479 	:	val_out <= 4'h2ff0;
         4'he47a 	:	val_out <= 4'h2ff0;
         4'he47b 	:	val_out <= 4'h2ff0;
         4'he480 	:	val_out <= 4'h3004;
         4'he481 	:	val_out <= 4'h3004;
         4'he482 	:	val_out <= 4'h3004;
         4'he483 	:	val_out <= 4'h3004;
         4'he488 	:	val_out <= 4'h3018;
         4'he489 	:	val_out <= 4'h3018;
         4'he48a 	:	val_out <= 4'h3018;
         4'he48b 	:	val_out <= 4'h3018;
         4'he490 	:	val_out <= 4'h302b;
         4'he491 	:	val_out <= 4'h302b;
         4'he492 	:	val_out <= 4'h302b;
         4'he493 	:	val_out <= 4'h302b;
         4'he498 	:	val_out <= 4'h303f;
         4'he499 	:	val_out <= 4'h303f;
         4'he49a 	:	val_out <= 4'h303f;
         4'he49b 	:	val_out <= 4'h303f;
         4'he4a0 	:	val_out <= 4'h3053;
         4'he4a1 	:	val_out <= 4'h3053;
         4'he4a2 	:	val_out <= 4'h3053;
         4'he4a3 	:	val_out <= 4'h3053;
         4'he4a8 	:	val_out <= 4'h3066;
         4'he4a9 	:	val_out <= 4'h3066;
         4'he4aa 	:	val_out <= 4'h3066;
         4'he4ab 	:	val_out <= 4'h3066;
         4'he4b0 	:	val_out <= 4'h307a;
         4'he4b1 	:	val_out <= 4'h307a;
         4'he4b2 	:	val_out <= 4'h307a;
         4'he4b3 	:	val_out <= 4'h307a;
         4'he4b8 	:	val_out <= 4'h308e;
         4'he4b9 	:	val_out <= 4'h308e;
         4'he4ba 	:	val_out <= 4'h308e;
         4'he4bb 	:	val_out <= 4'h308e;
         4'he4c0 	:	val_out <= 4'h30a1;
         4'he4c1 	:	val_out <= 4'h30a1;
         4'he4c2 	:	val_out <= 4'h30a1;
         4'he4c3 	:	val_out <= 4'h30a1;
         4'he4c8 	:	val_out <= 4'h30b5;
         4'he4c9 	:	val_out <= 4'h30b5;
         4'he4ca 	:	val_out <= 4'h30b5;
         4'he4cb 	:	val_out <= 4'h30b5;
         4'he4d0 	:	val_out <= 4'h30c9;
         4'he4d1 	:	val_out <= 4'h30c9;
         4'he4d2 	:	val_out <= 4'h30c9;
         4'he4d3 	:	val_out <= 4'h30c9;
         4'he4d8 	:	val_out <= 4'h30dd;
         4'he4d9 	:	val_out <= 4'h30dd;
         4'he4da 	:	val_out <= 4'h30dd;
         4'he4db 	:	val_out <= 4'h30dd;
         4'he4e0 	:	val_out <= 4'h30f0;
         4'he4e1 	:	val_out <= 4'h30f0;
         4'he4e2 	:	val_out <= 4'h30f0;
         4'he4e3 	:	val_out <= 4'h30f0;
         4'he4e8 	:	val_out <= 4'h3104;
         4'he4e9 	:	val_out <= 4'h3104;
         4'he4ea 	:	val_out <= 4'h3104;
         4'he4eb 	:	val_out <= 4'h3104;
         4'he4f0 	:	val_out <= 4'h3118;
         4'he4f1 	:	val_out <= 4'h3118;
         4'he4f2 	:	val_out <= 4'h3118;
         4'he4f3 	:	val_out <= 4'h3118;
         4'he4f8 	:	val_out <= 4'h312c;
         4'he4f9 	:	val_out <= 4'h312c;
         4'he4fa 	:	val_out <= 4'h312c;
         4'he4fb 	:	val_out <= 4'h312c;
         4'he500 	:	val_out <= 4'h3140;
         4'he501 	:	val_out <= 4'h3140;
         4'he502 	:	val_out <= 4'h3140;
         4'he503 	:	val_out <= 4'h3140;
         4'he508 	:	val_out <= 4'h3153;
         4'he509 	:	val_out <= 4'h3153;
         4'he50a 	:	val_out <= 4'h3153;
         4'he50b 	:	val_out <= 4'h3153;
         4'he510 	:	val_out <= 4'h3167;
         4'he511 	:	val_out <= 4'h3167;
         4'he512 	:	val_out <= 4'h3167;
         4'he513 	:	val_out <= 4'h3167;
         4'he518 	:	val_out <= 4'h317b;
         4'he519 	:	val_out <= 4'h317b;
         4'he51a 	:	val_out <= 4'h317b;
         4'he51b 	:	val_out <= 4'h317b;
         4'he520 	:	val_out <= 4'h318f;
         4'he521 	:	val_out <= 4'h318f;
         4'he522 	:	val_out <= 4'h318f;
         4'he523 	:	val_out <= 4'h318f;
         4'he528 	:	val_out <= 4'h31a3;
         4'he529 	:	val_out <= 4'h31a3;
         4'he52a 	:	val_out <= 4'h31a3;
         4'he52b 	:	val_out <= 4'h31a3;
         4'he530 	:	val_out <= 4'h31b7;
         4'he531 	:	val_out <= 4'h31b7;
         4'he532 	:	val_out <= 4'h31b7;
         4'he533 	:	val_out <= 4'h31b7;
         4'he538 	:	val_out <= 4'h31cb;
         4'he539 	:	val_out <= 4'h31cb;
         4'he53a 	:	val_out <= 4'h31cb;
         4'he53b 	:	val_out <= 4'h31cb;
         4'he540 	:	val_out <= 4'h31de;
         4'he541 	:	val_out <= 4'h31de;
         4'he542 	:	val_out <= 4'h31de;
         4'he543 	:	val_out <= 4'h31de;
         4'he548 	:	val_out <= 4'h31f2;
         4'he549 	:	val_out <= 4'h31f2;
         4'he54a 	:	val_out <= 4'h31f2;
         4'he54b 	:	val_out <= 4'h31f2;
         4'he550 	:	val_out <= 4'h3206;
         4'he551 	:	val_out <= 4'h3206;
         4'he552 	:	val_out <= 4'h3206;
         4'he553 	:	val_out <= 4'h3206;
         4'he558 	:	val_out <= 4'h321a;
         4'he559 	:	val_out <= 4'h321a;
         4'he55a 	:	val_out <= 4'h321a;
         4'he55b 	:	val_out <= 4'h321a;
         4'he560 	:	val_out <= 4'h322e;
         4'he561 	:	val_out <= 4'h322e;
         4'he562 	:	val_out <= 4'h322e;
         4'he563 	:	val_out <= 4'h322e;
         4'he568 	:	val_out <= 4'h3242;
         4'he569 	:	val_out <= 4'h3242;
         4'he56a 	:	val_out <= 4'h3242;
         4'he56b 	:	val_out <= 4'h3242;
         4'he570 	:	val_out <= 4'h3256;
         4'he571 	:	val_out <= 4'h3256;
         4'he572 	:	val_out <= 4'h3256;
         4'he573 	:	val_out <= 4'h3256;
         4'he578 	:	val_out <= 4'h326a;
         4'he579 	:	val_out <= 4'h326a;
         4'he57a 	:	val_out <= 4'h326a;
         4'he57b 	:	val_out <= 4'h326a;
         4'he580 	:	val_out <= 4'h327e;
         4'he581 	:	val_out <= 4'h327e;
         4'he582 	:	val_out <= 4'h327e;
         4'he583 	:	val_out <= 4'h327e;
         4'he588 	:	val_out <= 4'h3292;
         4'he589 	:	val_out <= 4'h3292;
         4'he58a 	:	val_out <= 4'h3292;
         4'he58b 	:	val_out <= 4'h3292;
         4'he590 	:	val_out <= 4'h32a6;
         4'he591 	:	val_out <= 4'h32a6;
         4'he592 	:	val_out <= 4'h32a6;
         4'he593 	:	val_out <= 4'h32a6;
         4'he598 	:	val_out <= 4'h32ba;
         4'he599 	:	val_out <= 4'h32ba;
         4'he59a 	:	val_out <= 4'h32ba;
         4'he59b 	:	val_out <= 4'h32ba;
         4'he5a0 	:	val_out <= 4'h32ce;
         4'he5a1 	:	val_out <= 4'h32ce;
         4'he5a2 	:	val_out <= 4'h32ce;
         4'he5a3 	:	val_out <= 4'h32ce;
         4'he5a8 	:	val_out <= 4'h32e2;
         4'he5a9 	:	val_out <= 4'h32e2;
         4'he5aa 	:	val_out <= 4'h32e2;
         4'he5ab 	:	val_out <= 4'h32e2;
         4'he5b0 	:	val_out <= 4'h32f6;
         4'he5b1 	:	val_out <= 4'h32f6;
         4'he5b2 	:	val_out <= 4'h32f6;
         4'he5b3 	:	val_out <= 4'h32f6;
         4'he5b8 	:	val_out <= 4'h330a;
         4'he5b9 	:	val_out <= 4'h330a;
         4'he5ba 	:	val_out <= 4'h330a;
         4'he5bb 	:	val_out <= 4'h330a;
         4'he5c0 	:	val_out <= 4'h331e;
         4'he5c1 	:	val_out <= 4'h331e;
         4'he5c2 	:	val_out <= 4'h331e;
         4'he5c3 	:	val_out <= 4'h331e;
         4'he5c8 	:	val_out <= 4'h3333;
         4'he5c9 	:	val_out <= 4'h3333;
         4'he5ca 	:	val_out <= 4'h3333;
         4'he5cb 	:	val_out <= 4'h3333;
         4'he5d0 	:	val_out <= 4'h3347;
         4'he5d1 	:	val_out <= 4'h3347;
         4'he5d2 	:	val_out <= 4'h3347;
         4'he5d3 	:	val_out <= 4'h3347;
         4'he5d8 	:	val_out <= 4'h335b;
         4'he5d9 	:	val_out <= 4'h335b;
         4'he5da 	:	val_out <= 4'h335b;
         4'he5db 	:	val_out <= 4'h335b;
         4'he5e0 	:	val_out <= 4'h336f;
         4'he5e1 	:	val_out <= 4'h336f;
         4'he5e2 	:	val_out <= 4'h336f;
         4'he5e3 	:	val_out <= 4'h336f;
         4'he5e8 	:	val_out <= 4'h3383;
         4'he5e9 	:	val_out <= 4'h3383;
         4'he5ea 	:	val_out <= 4'h3383;
         4'he5eb 	:	val_out <= 4'h3383;
         4'he5f0 	:	val_out <= 4'h3397;
         4'he5f1 	:	val_out <= 4'h3397;
         4'he5f2 	:	val_out <= 4'h3397;
         4'he5f3 	:	val_out <= 4'h3397;
         4'he5f8 	:	val_out <= 4'h33ab;
         4'he5f9 	:	val_out <= 4'h33ab;
         4'he5fa 	:	val_out <= 4'h33ab;
         4'he5fb 	:	val_out <= 4'h33ab;
         4'he600 	:	val_out <= 4'h33c0;
         4'he601 	:	val_out <= 4'h33c0;
         4'he602 	:	val_out <= 4'h33c0;
         4'he603 	:	val_out <= 4'h33c0;
         4'he608 	:	val_out <= 4'h33d4;
         4'he609 	:	val_out <= 4'h33d4;
         4'he60a 	:	val_out <= 4'h33d4;
         4'he60b 	:	val_out <= 4'h33d4;
         4'he610 	:	val_out <= 4'h33e8;
         4'he611 	:	val_out <= 4'h33e8;
         4'he612 	:	val_out <= 4'h33e8;
         4'he613 	:	val_out <= 4'h33e8;
         4'he618 	:	val_out <= 4'h33fc;
         4'he619 	:	val_out <= 4'h33fc;
         4'he61a 	:	val_out <= 4'h33fc;
         4'he61b 	:	val_out <= 4'h33fc;
         4'he620 	:	val_out <= 4'h3410;
         4'he621 	:	val_out <= 4'h3410;
         4'he622 	:	val_out <= 4'h3410;
         4'he623 	:	val_out <= 4'h3410;
         4'he628 	:	val_out <= 4'h3425;
         4'he629 	:	val_out <= 4'h3425;
         4'he62a 	:	val_out <= 4'h3425;
         4'he62b 	:	val_out <= 4'h3425;
         4'he630 	:	val_out <= 4'h3439;
         4'he631 	:	val_out <= 4'h3439;
         4'he632 	:	val_out <= 4'h3439;
         4'he633 	:	val_out <= 4'h3439;
         4'he638 	:	val_out <= 4'h344d;
         4'he639 	:	val_out <= 4'h344d;
         4'he63a 	:	val_out <= 4'h344d;
         4'he63b 	:	val_out <= 4'h344d;
         4'he640 	:	val_out <= 4'h3461;
         4'he641 	:	val_out <= 4'h3461;
         4'he642 	:	val_out <= 4'h3461;
         4'he643 	:	val_out <= 4'h3461;
         4'he648 	:	val_out <= 4'h3476;
         4'he649 	:	val_out <= 4'h3476;
         4'he64a 	:	val_out <= 4'h3476;
         4'he64b 	:	val_out <= 4'h3476;
         4'he650 	:	val_out <= 4'h348a;
         4'he651 	:	val_out <= 4'h348a;
         4'he652 	:	val_out <= 4'h348a;
         4'he653 	:	val_out <= 4'h348a;
         4'he658 	:	val_out <= 4'h349e;
         4'he659 	:	val_out <= 4'h349e;
         4'he65a 	:	val_out <= 4'h349e;
         4'he65b 	:	val_out <= 4'h349e;
         4'he660 	:	val_out <= 4'h34b3;
         4'he661 	:	val_out <= 4'h34b3;
         4'he662 	:	val_out <= 4'h34b3;
         4'he663 	:	val_out <= 4'h34b3;
         4'he668 	:	val_out <= 4'h34c7;
         4'he669 	:	val_out <= 4'h34c7;
         4'he66a 	:	val_out <= 4'h34c7;
         4'he66b 	:	val_out <= 4'h34c7;
         4'he670 	:	val_out <= 4'h34db;
         4'he671 	:	val_out <= 4'h34db;
         4'he672 	:	val_out <= 4'h34db;
         4'he673 	:	val_out <= 4'h34db;
         4'he678 	:	val_out <= 4'h34f0;
         4'he679 	:	val_out <= 4'h34f0;
         4'he67a 	:	val_out <= 4'h34f0;
         4'he67b 	:	val_out <= 4'h34f0;
         4'he680 	:	val_out <= 4'h3504;
         4'he681 	:	val_out <= 4'h3504;
         4'he682 	:	val_out <= 4'h3504;
         4'he683 	:	val_out <= 4'h3504;
         4'he688 	:	val_out <= 4'h3518;
         4'he689 	:	val_out <= 4'h3518;
         4'he68a 	:	val_out <= 4'h3518;
         4'he68b 	:	val_out <= 4'h3518;
         4'he690 	:	val_out <= 4'h352d;
         4'he691 	:	val_out <= 4'h352d;
         4'he692 	:	val_out <= 4'h352d;
         4'he693 	:	val_out <= 4'h352d;
         4'he698 	:	val_out <= 4'h3541;
         4'he699 	:	val_out <= 4'h3541;
         4'he69a 	:	val_out <= 4'h3541;
         4'he69b 	:	val_out <= 4'h3541;
         4'he6a0 	:	val_out <= 4'h3556;
         4'he6a1 	:	val_out <= 4'h3556;
         4'he6a2 	:	val_out <= 4'h3556;
         4'he6a3 	:	val_out <= 4'h3556;
         4'he6a8 	:	val_out <= 4'h356a;
         4'he6a9 	:	val_out <= 4'h356a;
         4'he6aa 	:	val_out <= 4'h356a;
         4'he6ab 	:	val_out <= 4'h356a;
         4'he6b0 	:	val_out <= 4'h357e;
         4'he6b1 	:	val_out <= 4'h357e;
         4'he6b2 	:	val_out <= 4'h357e;
         4'he6b3 	:	val_out <= 4'h357e;
         4'he6b8 	:	val_out <= 4'h3593;
         4'he6b9 	:	val_out <= 4'h3593;
         4'he6ba 	:	val_out <= 4'h3593;
         4'he6bb 	:	val_out <= 4'h3593;
         4'he6c0 	:	val_out <= 4'h35a7;
         4'he6c1 	:	val_out <= 4'h35a7;
         4'he6c2 	:	val_out <= 4'h35a7;
         4'he6c3 	:	val_out <= 4'h35a7;
         4'he6c8 	:	val_out <= 4'h35bc;
         4'he6c9 	:	val_out <= 4'h35bc;
         4'he6ca 	:	val_out <= 4'h35bc;
         4'he6cb 	:	val_out <= 4'h35bc;
         4'he6d0 	:	val_out <= 4'h35d0;
         4'he6d1 	:	val_out <= 4'h35d0;
         4'he6d2 	:	val_out <= 4'h35d0;
         4'he6d3 	:	val_out <= 4'h35d0;
         4'he6d8 	:	val_out <= 4'h35e5;
         4'he6d9 	:	val_out <= 4'h35e5;
         4'he6da 	:	val_out <= 4'h35e5;
         4'he6db 	:	val_out <= 4'h35e5;
         4'he6e0 	:	val_out <= 4'h35f9;
         4'he6e1 	:	val_out <= 4'h35f9;
         4'he6e2 	:	val_out <= 4'h35f9;
         4'he6e3 	:	val_out <= 4'h35f9;
         4'he6e8 	:	val_out <= 4'h360e;
         4'he6e9 	:	val_out <= 4'h360e;
         4'he6ea 	:	val_out <= 4'h360e;
         4'he6eb 	:	val_out <= 4'h360e;
         4'he6f0 	:	val_out <= 4'h3622;
         4'he6f1 	:	val_out <= 4'h3622;
         4'he6f2 	:	val_out <= 4'h3622;
         4'he6f3 	:	val_out <= 4'h3622;
         4'he6f8 	:	val_out <= 4'h3637;
         4'he6f9 	:	val_out <= 4'h3637;
         4'he6fa 	:	val_out <= 4'h3637;
         4'he6fb 	:	val_out <= 4'h3637;
         4'he700 	:	val_out <= 4'h364b;
         4'he701 	:	val_out <= 4'h364b;
         4'he702 	:	val_out <= 4'h364b;
         4'he703 	:	val_out <= 4'h364b;
         4'he708 	:	val_out <= 4'h3660;
         4'he709 	:	val_out <= 4'h3660;
         4'he70a 	:	val_out <= 4'h3660;
         4'he70b 	:	val_out <= 4'h3660;
         4'he710 	:	val_out <= 4'h3675;
         4'he711 	:	val_out <= 4'h3675;
         4'he712 	:	val_out <= 4'h3675;
         4'he713 	:	val_out <= 4'h3675;
         4'he718 	:	val_out <= 4'h3689;
         4'he719 	:	val_out <= 4'h3689;
         4'he71a 	:	val_out <= 4'h3689;
         4'he71b 	:	val_out <= 4'h3689;
         4'he720 	:	val_out <= 4'h369e;
         4'he721 	:	val_out <= 4'h369e;
         4'he722 	:	val_out <= 4'h369e;
         4'he723 	:	val_out <= 4'h369e;
         4'he728 	:	val_out <= 4'h36b2;
         4'he729 	:	val_out <= 4'h36b2;
         4'he72a 	:	val_out <= 4'h36b2;
         4'he72b 	:	val_out <= 4'h36b2;
         4'he730 	:	val_out <= 4'h36c7;
         4'he731 	:	val_out <= 4'h36c7;
         4'he732 	:	val_out <= 4'h36c7;
         4'he733 	:	val_out <= 4'h36c7;
         4'he738 	:	val_out <= 4'h36dc;
         4'he739 	:	val_out <= 4'h36dc;
         4'he73a 	:	val_out <= 4'h36dc;
         4'he73b 	:	val_out <= 4'h36dc;
         4'he740 	:	val_out <= 4'h36f0;
         4'he741 	:	val_out <= 4'h36f0;
         4'he742 	:	val_out <= 4'h36f0;
         4'he743 	:	val_out <= 4'h36f0;
         4'he748 	:	val_out <= 4'h3705;
         4'he749 	:	val_out <= 4'h3705;
         4'he74a 	:	val_out <= 4'h3705;
         4'he74b 	:	val_out <= 4'h3705;
         4'he750 	:	val_out <= 4'h3719;
         4'he751 	:	val_out <= 4'h3719;
         4'he752 	:	val_out <= 4'h3719;
         4'he753 	:	val_out <= 4'h3719;
         4'he758 	:	val_out <= 4'h372e;
         4'he759 	:	val_out <= 4'h372e;
         4'he75a 	:	val_out <= 4'h372e;
         4'he75b 	:	val_out <= 4'h372e;
         4'he760 	:	val_out <= 4'h3743;
         4'he761 	:	val_out <= 4'h3743;
         4'he762 	:	val_out <= 4'h3743;
         4'he763 	:	val_out <= 4'h3743;
         4'he768 	:	val_out <= 4'h3757;
         4'he769 	:	val_out <= 4'h3757;
         4'he76a 	:	val_out <= 4'h3757;
         4'he76b 	:	val_out <= 4'h3757;
         4'he770 	:	val_out <= 4'h376c;
         4'he771 	:	val_out <= 4'h376c;
         4'he772 	:	val_out <= 4'h376c;
         4'he773 	:	val_out <= 4'h376c;
         4'he778 	:	val_out <= 4'h3781;
         4'he779 	:	val_out <= 4'h3781;
         4'he77a 	:	val_out <= 4'h3781;
         4'he77b 	:	val_out <= 4'h3781;
         4'he780 	:	val_out <= 4'h3796;
         4'he781 	:	val_out <= 4'h3796;
         4'he782 	:	val_out <= 4'h3796;
         4'he783 	:	val_out <= 4'h3796;
         4'he788 	:	val_out <= 4'h37aa;
         4'he789 	:	val_out <= 4'h37aa;
         4'he78a 	:	val_out <= 4'h37aa;
         4'he78b 	:	val_out <= 4'h37aa;
         4'he790 	:	val_out <= 4'h37bf;
         4'he791 	:	val_out <= 4'h37bf;
         4'he792 	:	val_out <= 4'h37bf;
         4'he793 	:	val_out <= 4'h37bf;
         4'he798 	:	val_out <= 4'h37d4;
         4'he799 	:	val_out <= 4'h37d4;
         4'he79a 	:	val_out <= 4'h37d4;
         4'he79b 	:	val_out <= 4'h37d4;
         4'he7a0 	:	val_out <= 4'h37e9;
         4'he7a1 	:	val_out <= 4'h37e9;
         4'he7a2 	:	val_out <= 4'h37e9;
         4'he7a3 	:	val_out <= 4'h37e9;
         4'he7a8 	:	val_out <= 4'h37fd;
         4'he7a9 	:	val_out <= 4'h37fd;
         4'he7aa 	:	val_out <= 4'h37fd;
         4'he7ab 	:	val_out <= 4'h37fd;
         4'he7b0 	:	val_out <= 4'h3812;
         4'he7b1 	:	val_out <= 4'h3812;
         4'he7b2 	:	val_out <= 4'h3812;
         4'he7b3 	:	val_out <= 4'h3812;
         4'he7b8 	:	val_out <= 4'h3827;
         4'he7b9 	:	val_out <= 4'h3827;
         4'he7ba 	:	val_out <= 4'h3827;
         4'he7bb 	:	val_out <= 4'h3827;
         4'he7c0 	:	val_out <= 4'h383c;
         4'he7c1 	:	val_out <= 4'h383c;
         4'he7c2 	:	val_out <= 4'h383c;
         4'he7c3 	:	val_out <= 4'h383c;
         4'he7c8 	:	val_out <= 4'h3851;
         4'he7c9 	:	val_out <= 4'h3851;
         4'he7ca 	:	val_out <= 4'h3851;
         4'he7cb 	:	val_out <= 4'h3851;
         4'he7d0 	:	val_out <= 4'h3865;
         4'he7d1 	:	val_out <= 4'h3865;
         4'he7d2 	:	val_out <= 4'h3865;
         4'he7d3 	:	val_out <= 4'h3865;
         4'he7d8 	:	val_out <= 4'h387a;
         4'he7d9 	:	val_out <= 4'h387a;
         4'he7da 	:	val_out <= 4'h387a;
         4'he7db 	:	val_out <= 4'h387a;
         4'he7e0 	:	val_out <= 4'h388f;
         4'he7e1 	:	val_out <= 4'h388f;
         4'he7e2 	:	val_out <= 4'h388f;
         4'he7e3 	:	val_out <= 4'h388f;
         4'he7e8 	:	val_out <= 4'h38a4;
         4'he7e9 	:	val_out <= 4'h38a4;
         4'he7ea 	:	val_out <= 4'h38a4;
         4'he7eb 	:	val_out <= 4'h38a4;
         4'he7f0 	:	val_out <= 4'h38b9;
         4'he7f1 	:	val_out <= 4'h38b9;
         4'he7f2 	:	val_out <= 4'h38b9;
         4'he7f3 	:	val_out <= 4'h38b9;
         4'he7f8 	:	val_out <= 4'h38ce;
         4'he7f9 	:	val_out <= 4'h38ce;
         4'he7fa 	:	val_out <= 4'h38ce;
         4'he7fb 	:	val_out <= 4'h38ce;
         4'he800 	:	val_out <= 4'h38e3;
         4'he801 	:	val_out <= 4'h38e3;
         4'he802 	:	val_out <= 4'h38e3;
         4'he803 	:	val_out <= 4'h38e3;
         4'he808 	:	val_out <= 4'h38f7;
         4'he809 	:	val_out <= 4'h38f7;
         4'he80a 	:	val_out <= 4'h38f7;
         4'he80b 	:	val_out <= 4'h38f7;
         4'he810 	:	val_out <= 4'h390c;
         4'he811 	:	val_out <= 4'h390c;
         4'he812 	:	val_out <= 4'h390c;
         4'he813 	:	val_out <= 4'h390c;
         4'he818 	:	val_out <= 4'h3921;
         4'he819 	:	val_out <= 4'h3921;
         4'he81a 	:	val_out <= 4'h3921;
         4'he81b 	:	val_out <= 4'h3921;
         4'he820 	:	val_out <= 4'h3936;
         4'he821 	:	val_out <= 4'h3936;
         4'he822 	:	val_out <= 4'h3936;
         4'he823 	:	val_out <= 4'h3936;
         4'he828 	:	val_out <= 4'h394b;
         4'he829 	:	val_out <= 4'h394b;
         4'he82a 	:	val_out <= 4'h394b;
         4'he82b 	:	val_out <= 4'h394b;
         4'he830 	:	val_out <= 4'h3960;
         4'he831 	:	val_out <= 4'h3960;
         4'he832 	:	val_out <= 4'h3960;
         4'he833 	:	val_out <= 4'h3960;
         4'he838 	:	val_out <= 4'h3975;
         4'he839 	:	val_out <= 4'h3975;
         4'he83a 	:	val_out <= 4'h3975;
         4'he83b 	:	val_out <= 4'h3975;
         4'he840 	:	val_out <= 4'h398a;
         4'he841 	:	val_out <= 4'h398a;
         4'he842 	:	val_out <= 4'h398a;
         4'he843 	:	val_out <= 4'h398a;
         4'he848 	:	val_out <= 4'h399f;
         4'he849 	:	val_out <= 4'h399f;
         4'he84a 	:	val_out <= 4'h399f;
         4'he84b 	:	val_out <= 4'h399f;
         4'he850 	:	val_out <= 4'h39b4;
         4'he851 	:	val_out <= 4'h39b4;
         4'he852 	:	val_out <= 4'h39b4;
         4'he853 	:	val_out <= 4'h39b4;
         4'he858 	:	val_out <= 4'h39c9;
         4'he859 	:	val_out <= 4'h39c9;
         4'he85a 	:	val_out <= 4'h39c9;
         4'he85b 	:	val_out <= 4'h39c9;
         4'he860 	:	val_out <= 4'h39de;
         4'he861 	:	val_out <= 4'h39de;
         4'he862 	:	val_out <= 4'h39de;
         4'he863 	:	val_out <= 4'h39de;
         4'he868 	:	val_out <= 4'h39f3;
         4'he869 	:	val_out <= 4'h39f3;
         4'he86a 	:	val_out <= 4'h39f3;
         4'he86b 	:	val_out <= 4'h39f3;
         4'he870 	:	val_out <= 4'h3a08;
         4'he871 	:	val_out <= 4'h3a08;
         4'he872 	:	val_out <= 4'h3a08;
         4'he873 	:	val_out <= 4'h3a08;
         4'he878 	:	val_out <= 4'h3a1d;
         4'he879 	:	val_out <= 4'h3a1d;
         4'he87a 	:	val_out <= 4'h3a1d;
         4'he87b 	:	val_out <= 4'h3a1d;
         4'he880 	:	val_out <= 4'h3a32;
         4'he881 	:	val_out <= 4'h3a32;
         4'he882 	:	val_out <= 4'h3a32;
         4'he883 	:	val_out <= 4'h3a32;
         4'he888 	:	val_out <= 4'h3a47;
         4'he889 	:	val_out <= 4'h3a47;
         4'he88a 	:	val_out <= 4'h3a47;
         4'he88b 	:	val_out <= 4'h3a47;
         4'he890 	:	val_out <= 4'h3a5c;
         4'he891 	:	val_out <= 4'h3a5c;
         4'he892 	:	val_out <= 4'h3a5c;
         4'he893 	:	val_out <= 4'h3a5c;
         4'he898 	:	val_out <= 4'h3a72;
         4'he899 	:	val_out <= 4'h3a72;
         4'he89a 	:	val_out <= 4'h3a72;
         4'he89b 	:	val_out <= 4'h3a72;
         4'he8a0 	:	val_out <= 4'h3a87;
         4'he8a1 	:	val_out <= 4'h3a87;
         4'he8a2 	:	val_out <= 4'h3a87;
         4'he8a3 	:	val_out <= 4'h3a87;
         4'he8a8 	:	val_out <= 4'h3a9c;
         4'he8a9 	:	val_out <= 4'h3a9c;
         4'he8aa 	:	val_out <= 4'h3a9c;
         4'he8ab 	:	val_out <= 4'h3a9c;
         4'he8b0 	:	val_out <= 4'h3ab1;
         4'he8b1 	:	val_out <= 4'h3ab1;
         4'he8b2 	:	val_out <= 4'h3ab1;
         4'he8b3 	:	val_out <= 4'h3ab1;
         4'he8b8 	:	val_out <= 4'h3ac6;
         4'he8b9 	:	val_out <= 4'h3ac6;
         4'he8ba 	:	val_out <= 4'h3ac6;
         4'he8bb 	:	val_out <= 4'h3ac6;
         4'he8c0 	:	val_out <= 4'h3adb;
         4'he8c1 	:	val_out <= 4'h3adb;
         4'he8c2 	:	val_out <= 4'h3adb;
         4'he8c3 	:	val_out <= 4'h3adb;
         4'he8c8 	:	val_out <= 4'h3af0;
         4'he8c9 	:	val_out <= 4'h3af0;
         4'he8ca 	:	val_out <= 4'h3af0;
         4'he8cb 	:	val_out <= 4'h3af0;
         4'he8d0 	:	val_out <= 4'h3b05;
         4'he8d1 	:	val_out <= 4'h3b05;
         4'he8d2 	:	val_out <= 4'h3b05;
         4'he8d3 	:	val_out <= 4'h3b05;
         4'he8d8 	:	val_out <= 4'h3b1b;
         4'he8d9 	:	val_out <= 4'h3b1b;
         4'he8da 	:	val_out <= 4'h3b1b;
         4'he8db 	:	val_out <= 4'h3b1b;
         4'he8e0 	:	val_out <= 4'h3b30;
         4'he8e1 	:	val_out <= 4'h3b30;
         4'he8e2 	:	val_out <= 4'h3b30;
         4'he8e3 	:	val_out <= 4'h3b30;
         4'he8e8 	:	val_out <= 4'h3b45;
         4'he8e9 	:	val_out <= 4'h3b45;
         4'he8ea 	:	val_out <= 4'h3b45;
         4'he8eb 	:	val_out <= 4'h3b45;
         4'he8f0 	:	val_out <= 4'h3b5a;
         4'he8f1 	:	val_out <= 4'h3b5a;
         4'he8f2 	:	val_out <= 4'h3b5a;
         4'he8f3 	:	val_out <= 4'h3b5a;
         4'he8f8 	:	val_out <= 4'h3b6f;
         4'he8f9 	:	val_out <= 4'h3b6f;
         4'he8fa 	:	val_out <= 4'h3b6f;
         4'he8fb 	:	val_out <= 4'h3b6f;
         4'he900 	:	val_out <= 4'h3b85;
         4'he901 	:	val_out <= 4'h3b85;
         4'he902 	:	val_out <= 4'h3b85;
         4'he903 	:	val_out <= 4'h3b85;
         4'he908 	:	val_out <= 4'h3b9a;
         4'he909 	:	val_out <= 4'h3b9a;
         4'he90a 	:	val_out <= 4'h3b9a;
         4'he90b 	:	val_out <= 4'h3b9a;
         4'he910 	:	val_out <= 4'h3baf;
         4'he911 	:	val_out <= 4'h3baf;
         4'he912 	:	val_out <= 4'h3baf;
         4'he913 	:	val_out <= 4'h3baf;
         4'he918 	:	val_out <= 4'h3bc4;
         4'he919 	:	val_out <= 4'h3bc4;
         4'he91a 	:	val_out <= 4'h3bc4;
         4'he91b 	:	val_out <= 4'h3bc4;
         4'he920 	:	val_out <= 4'h3bda;
         4'he921 	:	val_out <= 4'h3bda;
         4'he922 	:	val_out <= 4'h3bda;
         4'he923 	:	val_out <= 4'h3bda;
         4'he928 	:	val_out <= 4'h3bef;
         4'he929 	:	val_out <= 4'h3bef;
         4'he92a 	:	val_out <= 4'h3bef;
         4'he92b 	:	val_out <= 4'h3bef;
         4'he930 	:	val_out <= 4'h3c04;
         4'he931 	:	val_out <= 4'h3c04;
         4'he932 	:	val_out <= 4'h3c04;
         4'he933 	:	val_out <= 4'h3c04;
         4'he938 	:	val_out <= 4'h3c1a;
         4'he939 	:	val_out <= 4'h3c1a;
         4'he93a 	:	val_out <= 4'h3c1a;
         4'he93b 	:	val_out <= 4'h3c1a;
         4'he940 	:	val_out <= 4'h3c2f;
         4'he941 	:	val_out <= 4'h3c2f;
         4'he942 	:	val_out <= 4'h3c2f;
         4'he943 	:	val_out <= 4'h3c2f;
         4'he948 	:	val_out <= 4'h3c44;
         4'he949 	:	val_out <= 4'h3c44;
         4'he94a 	:	val_out <= 4'h3c44;
         4'he94b 	:	val_out <= 4'h3c44;
         4'he950 	:	val_out <= 4'h3c5a;
         4'he951 	:	val_out <= 4'h3c5a;
         4'he952 	:	val_out <= 4'h3c5a;
         4'he953 	:	val_out <= 4'h3c5a;
         4'he958 	:	val_out <= 4'h3c6f;
         4'he959 	:	val_out <= 4'h3c6f;
         4'he95a 	:	val_out <= 4'h3c6f;
         4'he95b 	:	val_out <= 4'h3c6f;
         4'he960 	:	val_out <= 4'h3c84;
         4'he961 	:	val_out <= 4'h3c84;
         4'he962 	:	val_out <= 4'h3c84;
         4'he963 	:	val_out <= 4'h3c84;
         4'he968 	:	val_out <= 4'h3c9a;
         4'he969 	:	val_out <= 4'h3c9a;
         4'he96a 	:	val_out <= 4'h3c9a;
         4'he96b 	:	val_out <= 4'h3c9a;
         4'he970 	:	val_out <= 4'h3caf;
         4'he971 	:	val_out <= 4'h3caf;
         4'he972 	:	val_out <= 4'h3caf;
         4'he973 	:	val_out <= 4'h3caf;
         4'he978 	:	val_out <= 4'h3cc4;
         4'he979 	:	val_out <= 4'h3cc4;
         4'he97a 	:	val_out <= 4'h3cc4;
         4'he97b 	:	val_out <= 4'h3cc4;
         4'he980 	:	val_out <= 4'h3cda;
         4'he981 	:	val_out <= 4'h3cda;
         4'he982 	:	val_out <= 4'h3cda;
         4'he983 	:	val_out <= 4'h3cda;
         4'he988 	:	val_out <= 4'h3cef;
         4'he989 	:	val_out <= 4'h3cef;
         4'he98a 	:	val_out <= 4'h3cef;
         4'he98b 	:	val_out <= 4'h3cef;
         4'he990 	:	val_out <= 4'h3d05;
         4'he991 	:	val_out <= 4'h3d05;
         4'he992 	:	val_out <= 4'h3d05;
         4'he993 	:	val_out <= 4'h3d05;
         4'he998 	:	val_out <= 4'h3d1a;
         4'he999 	:	val_out <= 4'h3d1a;
         4'he99a 	:	val_out <= 4'h3d1a;
         4'he99b 	:	val_out <= 4'h3d1a;
         4'he9a0 	:	val_out <= 4'h3d2f;
         4'he9a1 	:	val_out <= 4'h3d2f;
         4'he9a2 	:	val_out <= 4'h3d2f;
         4'he9a3 	:	val_out <= 4'h3d2f;
         4'he9a8 	:	val_out <= 4'h3d45;
         4'he9a9 	:	val_out <= 4'h3d45;
         4'he9aa 	:	val_out <= 4'h3d45;
         4'he9ab 	:	val_out <= 4'h3d45;
         4'he9b0 	:	val_out <= 4'h3d5a;
         4'he9b1 	:	val_out <= 4'h3d5a;
         4'he9b2 	:	val_out <= 4'h3d5a;
         4'he9b3 	:	val_out <= 4'h3d5a;
         4'he9b8 	:	val_out <= 4'h3d70;
         4'he9b9 	:	val_out <= 4'h3d70;
         4'he9ba 	:	val_out <= 4'h3d70;
         4'he9bb 	:	val_out <= 4'h3d70;
         4'he9c0 	:	val_out <= 4'h3d85;
         4'he9c1 	:	val_out <= 4'h3d85;
         4'he9c2 	:	val_out <= 4'h3d85;
         4'he9c3 	:	val_out <= 4'h3d85;
         4'he9c8 	:	val_out <= 4'h3d9b;
         4'he9c9 	:	val_out <= 4'h3d9b;
         4'he9ca 	:	val_out <= 4'h3d9b;
         4'he9cb 	:	val_out <= 4'h3d9b;
         4'he9d0 	:	val_out <= 4'h3db0;
         4'he9d1 	:	val_out <= 4'h3db0;
         4'he9d2 	:	val_out <= 4'h3db0;
         4'he9d3 	:	val_out <= 4'h3db0;
         4'he9d8 	:	val_out <= 4'h3dc6;
         4'he9d9 	:	val_out <= 4'h3dc6;
         4'he9da 	:	val_out <= 4'h3dc6;
         4'he9db 	:	val_out <= 4'h3dc6;
         4'he9e0 	:	val_out <= 4'h3ddb;
         4'he9e1 	:	val_out <= 4'h3ddb;
         4'he9e2 	:	val_out <= 4'h3ddb;
         4'he9e3 	:	val_out <= 4'h3ddb;
         4'he9e8 	:	val_out <= 4'h3df1;
         4'he9e9 	:	val_out <= 4'h3df1;
         4'he9ea 	:	val_out <= 4'h3df1;
         4'he9eb 	:	val_out <= 4'h3df1;
         4'he9f0 	:	val_out <= 4'h3e06;
         4'he9f1 	:	val_out <= 4'h3e06;
         4'he9f2 	:	val_out <= 4'h3e06;
         4'he9f3 	:	val_out <= 4'h3e06;
         4'he9f8 	:	val_out <= 4'h3e1c;
         4'he9f9 	:	val_out <= 4'h3e1c;
         4'he9fa 	:	val_out <= 4'h3e1c;
         4'he9fb 	:	val_out <= 4'h3e1c;
         4'hea00 	:	val_out <= 4'h3e31;
         4'hea01 	:	val_out <= 4'h3e31;
         4'hea02 	:	val_out <= 4'h3e31;
         4'hea03 	:	val_out <= 4'h3e31;
         4'hea08 	:	val_out <= 4'h3e47;
         4'hea09 	:	val_out <= 4'h3e47;
         4'hea0a 	:	val_out <= 4'h3e47;
         4'hea0b 	:	val_out <= 4'h3e47;
         4'hea10 	:	val_out <= 4'h3e5d;
         4'hea11 	:	val_out <= 4'h3e5d;
         4'hea12 	:	val_out <= 4'h3e5d;
         4'hea13 	:	val_out <= 4'h3e5d;
         4'hea18 	:	val_out <= 4'h3e72;
         4'hea19 	:	val_out <= 4'h3e72;
         4'hea1a 	:	val_out <= 4'h3e72;
         4'hea1b 	:	val_out <= 4'h3e72;
         4'hea20 	:	val_out <= 4'h3e88;
         4'hea21 	:	val_out <= 4'h3e88;
         4'hea22 	:	val_out <= 4'h3e88;
         4'hea23 	:	val_out <= 4'h3e88;
         4'hea28 	:	val_out <= 4'h3e9d;
         4'hea29 	:	val_out <= 4'h3e9d;
         4'hea2a 	:	val_out <= 4'h3e9d;
         4'hea2b 	:	val_out <= 4'h3e9d;
         4'hea30 	:	val_out <= 4'h3eb3;
         4'hea31 	:	val_out <= 4'h3eb3;
         4'hea32 	:	val_out <= 4'h3eb3;
         4'hea33 	:	val_out <= 4'h3eb3;
         4'hea38 	:	val_out <= 4'h3ec9;
         4'hea39 	:	val_out <= 4'h3ec9;
         4'hea3a 	:	val_out <= 4'h3ec9;
         4'hea3b 	:	val_out <= 4'h3ec9;
         4'hea40 	:	val_out <= 4'h3ede;
         4'hea41 	:	val_out <= 4'h3ede;
         4'hea42 	:	val_out <= 4'h3ede;
         4'hea43 	:	val_out <= 4'h3ede;
         4'hea48 	:	val_out <= 4'h3ef4;
         4'hea49 	:	val_out <= 4'h3ef4;
         4'hea4a 	:	val_out <= 4'h3ef4;
         4'hea4b 	:	val_out <= 4'h3ef4;
         4'hea50 	:	val_out <= 4'h3f09;
         4'hea51 	:	val_out <= 4'h3f09;
         4'hea52 	:	val_out <= 4'h3f09;
         4'hea53 	:	val_out <= 4'h3f09;
         4'hea58 	:	val_out <= 4'h3f1f;
         4'hea59 	:	val_out <= 4'h3f1f;
         4'hea5a 	:	val_out <= 4'h3f1f;
         4'hea5b 	:	val_out <= 4'h3f1f;
         4'hea60 	:	val_out <= 4'h3f35;
         4'hea61 	:	val_out <= 4'h3f35;
         4'hea62 	:	val_out <= 4'h3f35;
         4'hea63 	:	val_out <= 4'h3f35;
         4'hea68 	:	val_out <= 4'h3f4a;
         4'hea69 	:	val_out <= 4'h3f4a;
         4'hea6a 	:	val_out <= 4'h3f4a;
         4'hea6b 	:	val_out <= 4'h3f4a;
         4'hea70 	:	val_out <= 4'h3f60;
         4'hea71 	:	val_out <= 4'h3f60;
         4'hea72 	:	val_out <= 4'h3f60;
         4'hea73 	:	val_out <= 4'h3f60;
         4'hea78 	:	val_out <= 4'h3f76;
         4'hea79 	:	val_out <= 4'h3f76;
         4'hea7a 	:	val_out <= 4'h3f76;
         4'hea7b 	:	val_out <= 4'h3f76;
         4'hea80 	:	val_out <= 4'h3f8c;
         4'hea81 	:	val_out <= 4'h3f8c;
         4'hea82 	:	val_out <= 4'h3f8c;
         4'hea83 	:	val_out <= 4'h3f8c;
         4'hea88 	:	val_out <= 4'h3fa1;
         4'hea89 	:	val_out <= 4'h3fa1;
         4'hea8a 	:	val_out <= 4'h3fa1;
         4'hea8b 	:	val_out <= 4'h3fa1;
         4'hea90 	:	val_out <= 4'h3fb7;
         4'hea91 	:	val_out <= 4'h3fb7;
         4'hea92 	:	val_out <= 4'h3fb7;
         4'hea93 	:	val_out <= 4'h3fb7;
         4'hea98 	:	val_out <= 4'h3fcd;
         4'hea99 	:	val_out <= 4'h3fcd;
         4'hea9a 	:	val_out <= 4'h3fcd;
         4'hea9b 	:	val_out <= 4'h3fcd;
         4'heaa0 	:	val_out <= 4'h3fe2;
         4'heaa1 	:	val_out <= 4'h3fe2;
         4'heaa2 	:	val_out <= 4'h3fe2;
         4'heaa3 	:	val_out <= 4'h3fe2;
         4'heaa8 	:	val_out <= 4'h3ff8;
         4'heaa9 	:	val_out <= 4'h3ff8;
         4'heaaa 	:	val_out <= 4'h3ff8;
         4'heaab 	:	val_out <= 4'h3ff8;
         4'heab0 	:	val_out <= 4'h400e;
         4'heab1 	:	val_out <= 4'h400e;
         4'heab2 	:	val_out <= 4'h400e;
         4'heab3 	:	val_out <= 4'h400e;
         4'heab8 	:	val_out <= 4'h4024;
         4'heab9 	:	val_out <= 4'h4024;
         4'heaba 	:	val_out <= 4'h4024;
         4'heabb 	:	val_out <= 4'h4024;
         4'heac0 	:	val_out <= 4'h403a;
         4'heac1 	:	val_out <= 4'h403a;
         4'heac2 	:	val_out <= 4'h403a;
         4'heac3 	:	val_out <= 4'h403a;
         4'heac8 	:	val_out <= 4'h404f;
         4'heac9 	:	val_out <= 4'h404f;
         4'heaca 	:	val_out <= 4'h404f;
         4'heacb 	:	val_out <= 4'h404f;
         4'head0 	:	val_out <= 4'h4065;
         4'head1 	:	val_out <= 4'h4065;
         4'head2 	:	val_out <= 4'h4065;
         4'head3 	:	val_out <= 4'h4065;
         4'head8 	:	val_out <= 4'h407b;
         4'head9 	:	val_out <= 4'h407b;
         4'heada 	:	val_out <= 4'h407b;
         4'headb 	:	val_out <= 4'h407b;
         4'heae0 	:	val_out <= 4'h4091;
         4'heae1 	:	val_out <= 4'h4091;
         4'heae2 	:	val_out <= 4'h4091;
         4'heae3 	:	val_out <= 4'h4091;
         4'heae8 	:	val_out <= 4'h40a7;
         4'heae9 	:	val_out <= 4'h40a7;
         4'heaea 	:	val_out <= 4'h40a7;
         4'heaeb 	:	val_out <= 4'h40a7;
         4'heaf0 	:	val_out <= 4'h40bc;
         4'heaf1 	:	val_out <= 4'h40bc;
         4'heaf2 	:	val_out <= 4'h40bc;
         4'heaf3 	:	val_out <= 4'h40bc;
         4'heaf8 	:	val_out <= 4'h40d2;
         4'heaf9 	:	val_out <= 4'h40d2;
         4'heafa 	:	val_out <= 4'h40d2;
         4'heafb 	:	val_out <= 4'h40d2;
         4'heb00 	:	val_out <= 4'h40e8;
         4'heb01 	:	val_out <= 4'h40e8;
         4'heb02 	:	val_out <= 4'h40e8;
         4'heb03 	:	val_out <= 4'h40e8;
         4'heb08 	:	val_out <= 4'h40fe;
         4'heb09 	:	val_out <= 4'h40fe;
         4'heb0a 	:	val_out <= 4'h40fe;
         4'heb0b 	:	val_out <= 4'h40fe;
         4'heb10 	:	val_out <= 4'h4114;
         4'heb11 	:	val_out <= 4'h4114;
         4'heb12 	:	val_out <= 4'h4114;
         4'heb13 	:	val_out <= 4'h4114;
         4'heb18 	:	val_out <= 4'h412a;
         4'heb19 	:	val_out <= 4'h412a;
         4'heb1a 	:	val_out <= 4'h412a;
         4'heb1b 	:	val_out <= 4'h412a;
         4'heb20 	:	val_out <= 4'h4140;
         4'heb21 	:	val_out <= 4'h4140;
         4'heb22 	:	val_out <= 4'h4140;
         4'heb23 	:	val_out <= 4'h4140;
         4'heb28 	:	val_out <= 4'h4156;
         4'heb29 	:	val_out <= 4'h4156;
         4'heb2a 	:	val_out <= 4'h4156;
         4'heb2b 	:	val_out <= 4'h4156;
         4'heb30 	:	val_out <= 4'h416c;
         4'heb31 	:	val_out <= 4'h416c;
         4'heb32 	:	val_out <= 4'h416c;
         4'heb33 	:	val_out <= 4'h416c;
         4'heb38 	:	val_out <= 4'h4182;
         4'heb39 	:	val_out <= 4'h4182;
         4'heb3a 	:	val_out <= 4'h4182;
         4'heb3b 	:	val_out <= 4'h4182;
         4'heb40 	:	val_out <= 4'h4197;
         4'heb41 	:	val_out <= 4'h4197;
         4'heb42 	:	val_out <= 4'h4197;
         4'heb43 	:	val_out <= 4'h4197;
         4'heb48 	:	val_out <= 4'h41ad;
         4'heb49 	:	val_out <= 4'h41ad;
         4'heb4a 	:	val_out <= 4'h41ad;
         4'heb4b 	:	val_out <= 4'h41ad;
         4'heb50 	:	val_out <= 4'h41c3;
         4'heb51 	:	val_out <= 4'h41c3;
         4'heb52 	:	val_out <= 4'h41c3;
         4'heb53 	:	val_out <= 4'h41c3;
         4'heb58 	:	val_out <= 4'h41d9;
         4'heb59 	:	val_out <= 4'h41d9;
         4'heb5a 	:	val_out <= 4'h41d9;
         4'heb5b 	:	val_out <= 4'h41d9;
         4'heb60 	:	val_out <= 4'h41ef;
         4'heb61 	:	val_out <= 4'h41ef;
         4'heb62 	:	val_out <= 4'h41ef;
         4'heb63 	:	val_out <= 4'h41ef;
         4'heb68 	:	val_out <= 4'h4205;
         4'heb69 	:	val_out <= 4'h4205;
         4'heb6a 	:	val_out <= 4'h4205;
         4'heb6b 	:	val_out <= 4'h4205;
         4'heb70 	:	val_out <= 4'h421b;
         4'heb71 	:	val_out <= 4'h421b;
         4'heb72 	:	val_out <= 4'h421b;
         4'heb73 	:	val_out <= 4'h421b;
         4'heb78 	:	val_out <= 4'h4231;
         4'heb79 	:	val_out <= 4'h4231;
         4'heb7a 	:	val_out <= 4'h4231;
         4'heb7b 	:	val_out <= 4'h4231;
         4'heb80 	:	val_out <= 4'h4247;
         4'heb81 	:	val_out <= 4'h4247;
         4'heb82 	:	val_out <= 4'h4247;
         4'heb83 	:	val_out <= 4'h4247;
         4'heb88 	:	val_out <= 4'h425d;
         4'heb89 	:	val_out <= 4'h425d;
         4'heb8a 	:	val_out <= 4'h425d;
         4'heb8b 	:	val_out <= 4'h425d;
         4'heb90 	:	val_out <= 4'h4273;
         4'heb91 	:	val_out <= 4'h4273;
         4'heb92 	:	val_out <= 4'h4273;
         4'heb93 	:	val_out <= 4'h4273;
         4'heb98 	:	val_out <= 4'h4289;
         4'heb99 	:	val_out <= 4'h4289;
         4'heb9a 	:	val_out <= 4'h4289;
         4'heb9b 	:	val_out <= 4'h4289;
         4'heba0 	:	val_out <= 4'h429f;
         4'heba1 	:	val_out <= 4'h429f;
         4'heba2 	:	val_out <= 4'h429f;
         4'heba3 	:	val_out <= 4'h429f;
         4'heba8 	:	val_out <= 4'h42b6;
         4'heba9 	:	val_out <= 4'h42b6;
         4'hebaa 	:	val_out <= 4'h42b6;
         4'hebab 	:	val_out <= 4'h42b6;
         4'hebb0 	:	val_out <= 4'h42cc;
         4'hebb1 	:	val_out <= 4'h42cc;
         4'hebb2 	:	val_out <= 4'h42cc;
         4'hebb3 	:	val_out <= 4'h42cc;
         4'hebb8 	:	val_out <= 4'h42e2;
         4'hebb9 	:	val_out <= 4'h42e2;
         4'hebba 	:	val_out <= 4'h42e2;
         4'hebbb 	:	val_out <= 4'h42e2;
         4'hebc0 	:	val_out <= 4'h42f8;
         4'hebc1 	:	val_out <= 4'h42f8;
         4'hebc2 	:	val_out <= 4'h42f8;
         4'hebc3 	:	val_out <= 4'h42f8;
         4'hebc8 	:	val_out <= 4'h430e;
         4'hebc9 	:	val_out <= 4'h430e;
         4'hebca 	:	val_out <= 4'h430e;
         4'hebcb 	:	val_out <= 4'h430e;
         4'hebd0 	:	val_out <= 4'h4324;
         4'hebd1 	:	val_out <= 4'h4324;
         4'hebd2 	:	val_out <= 4'h4324;
         4'hebd3 	:	val_out <= 4'h4324;
         4'hebd8 	:	val_out <= 4'h433a;
         4'hebd9 	:	val_out <= 4'h433a;
         4'hebda 	:	val_out <= 4'h433a;
         4'hebdb 	:	val_out <= 4'h433a;
         4'hebe0 	:	val_out <= 4'h4350;
         4'hebe1 	:	val_out <= 4'h4350;
         4'hebe2 	:	val_out <= 4'h4350;
         4'hebe3 	:	val_out <= 4'h4350;
         4'hebe8 	:	val_out <= 4'h4366;
         4'hebe9 	:	val_out <= 4'h4366;
         4'hebea 	:	val_out <= 4'h4366;
         4'hebeb 	:	val_out <= 4'h4366;
         4'hebf0 	:	val_out <= 4'h437c;
         4'hebf1 	:	val_out <= 4'h437c;
         4'hebf2 	:	val_out <= 4'h437c;
         4'hebf3 	:	val_out <= 4'h437c;
         4'hebf8 	:	val_out <= 4'h4393;
         4'hebf9 	:	val_out <= 4'h4393;
         4'hebfa 	:	val_out <= 4'h4393;
         4'hebfb 	:	val_out <= 4'h4393;
         4'hec00 	:	val_out <= 4'h43a9;
         4'hec01 	:	val_out <= 4'h43a9;
         4'hec02 	:	val_out <= 4'h43a9;
         4'hec03 	:	val_out <= 4'h43a9;
         4'hec08 	:	val_out <= 4'h43bf;
         4'hec09 	:	val_out <= 4'h43bf;
         4'hec0a 	:	val_out <= 4'h43bf;
         4'hec0b 	:	val_out <= 4'h43bf;
         4'hec10 	:	val_out <= 4'h43d5;
         4'hec11 	:	val_out <= 4'h43d5;
         4'hec12 	:	val_out <= 4'h43d5;
         4'hec13 	:	val_out <= 4'h43d5;
         4'hec18 	:	val_out <= 4'h43eb;
         4'hec19 	:	val_out <= 4'h43eb;
         4'hec1a 	:	val_out <= 4'h43eb;
         4'hec1b 	:	val_out <= 4'h43eb;
         4'hec20 	:	val_out <= 4'h4402;
         4'hec21 	:	val_out <= 4'h4402;
         4'hec22 	:	val_out <= 4'h4402;
         4'hec23 	:	val_out <= 4'h4402;
         4'hec28 	:	val_out <= 4'h4418;
         4'hec29 	:	val_out <= 4'h4418;
         4'hec2a 	:	val_out <= 4'h4418;
         4'hec2b 	:	val_out <= 4'h4418;
         4'hec30 	:	val_out <= 4'h442e;
         4'hec31 	:	val_out <= 4'h442e;
         4'hec32 	:	val_out <= 4'h442e;
         4'hec33 	:	val_out <= 4'h442e;
         4'hec38 	:	val_out <= 4'h4444;
         4'hec39 	:	val_out <= 4'h4444;
         4'hec3a 	:	val_out <= 4'h4444;
         4'hec3b 	:	val_out <= 4'h4444;
         4'hec40 	:	val_out <= 4'h445a;
         4'hec41 	:	val_out <= 4'h445a;
         4'hec42 	:	val_out <= 4'h445a;
         4'hec43 	:	val_out <= 4'h445a;
         4'hec48 	:	val_out <= 4'h4471;
         4'hec49 	:	val_out <= 4'h4471;
         4'hec4a 	:	val_out <= 4'h4471;
         4'hec4b 	:	val_out <= 4'h4471;
         4'hec50 	:	val_out <= 4'h4487;
         4'hec51 	:	val_out <= 4'h4487;
         4'hec52 	:	val_out <= 4'h4487;
         4'hec53 	:	val_out <= 4'h4487;
         4'hec58 	:	val_out <= 4'h449d;
         4'hec59 	:	val_out <= 4'h449d;
         4'hec5a 	:	val_out <= 4'h449d;
         4'hec5b 	:	val_out <= 4'h449d;
         4'hec60 	:	val_out <= 4'h44b3;
         4'hec61 	:	val_out <= 4'h44b3;
         4'hec62 	:	val_out <= 4'h44b3;
         4'hec63 	:	val_out <= 4'h44b3;
         4'hec68 	:	val_out <= 4'h44ca;
         4'hec69 	:	val_out <= 4'h44ca;
         4'hec6a 	:	val_out <= 4'h44ca;
         4'hec6b 	:	val_out <= 4'h44ca;
         4'hec70 	:	val_out <= 4'h44e0;
         4'hec71 	:	val_out <= 4'h44e0;
         4'hec72 	:	val_out <= 4'h44e0;
         4'hec73 	:	val_out <= 4'h44e0;
         4'hec78 	:	val_out <= 4'h44f6;
         4'hec79 	:	val_out <= 4'h44f6;
         4'hec7a 	:	val_out <= 4'h44f6;
         4'hec7b 	:	val_out <= 4'h44f6;
         4'hec80 	:	val_out <= 4'h450d;
         4'hec81 	:	val_out <= 4'h450d;
         4'hec82 	:	val_out <= 4'h450d;
         4'hec83 	:	val_out <= 4'h450d;
         4'hec88 	:	val_out <= 4'h4523;
         4'hec89 	:	val_out <= 4'h4523;
         4'hec8a 	:	val_out <= 4'h4523;
         4'hec8b 	:	val_out <= 4'h4523;
         4'hec90 	:	val_out <= 4'h4539;
         4'hec91 	:	val_out <= 4'h4539;
         4'hec92 	:	val_out <= 4'h4539;
         4'hec93 	:	val_out <= 4'h4539;
         4'hec98 	:	val_out <= 4'h4550;
         4'hec99 	:	val_out <= 4'h4550;
         4'hec9a 	:	val_out <= 4'h4550;
         4'hec9b 	:	val_out <= 4'h4550;
         4'heca0 	:	val_out <= 4'h4566;
         4'heca1 	:	val_out <= 4'h4566;
         4'heca2 	:	val_out <= 4'h4566;
         4'heca3 	:	val_out <= 4'h4566;
         4'heca8 	:	val_out <= 4'h457c;
         4'heca9 	:	val_out <= 4'h457c;
         4'hecaa 	:	val_out <= 4'h457c;
         4'hecab 	:	val_out <= 4'h457c;
         4'hecb0 	:	val_out <= 4'h4593;
         4'hecb1 	:	val_out <= 4'h4593;
         4'hecb2 	:	val_out <= 4'h4593;
         4'hecb3 	:	val_out <= 4'h4593;
         4'hecb8 	:	val_out <= 4'h45a9;
         4'hecb9 	:	val_out <= 4'h45a9;
         4'hecba 	:	val_out <= 4'h45a9;
         4'hecbb 	:	val_out <= 4'h45a9;
         4'hecc0 	:	val_out <= 4'h45bf;
         4'hecc1 	:	val_out <= 4'h45bf;
         4'hecc2 	:	val_out <= 4'h45bf;
         4'hecc3 	:	val_out <= 4'h45bf;
         4'hecc8 	:	val_out <= 4'h45d6;
         4'hecc9 	:	val_out <= 4'h45d6;
         4'hecca 	:	val_out <= 4'h45d6;
         4'heccb 	:	val_out <= 4'h45d6;
         4'hecd0 	:	val_out <= 4'h45ec;
         4'hecd1 	:	val_out <= 4'h45ec;
         4'hecd2 	:	val_out <= 4'h45ec;
         4'hecd3 	:	val_out <= 4'h45ec;
         4'hecd8 	:	val_out <= 4'h4602;
         4'hecd9 	:	val_out <= 4'h4602;
         4'hecda 	:	val_out <= 4'h4602;
         4'hecdb 	:	val_out <= 4'h4602;
         4'hece0 	:	val_out <= 4'h4619;
         4'hece1 	:	val_out <= 4'h4619;
         4'hece2 	:	val_out <= 4'h4619;
         4'hece3 	:	val_out <= 4'h4619;
         4'hece8 	:	val_out <= 4'h462f;
         4'hece9 	:	val_out <= 4'h462f;
         4'hecea 	:	val_out <= 4'h462f;
         4'heceb 	:	val_out <= 4'h462f;
         4'hecf0 	:	val_out <= 4'h4646;
         4'hecf1 	:	val_out <= 4'h4646;
         4'hecf2 	:	val_out <= 4'h4646;
         4'hecf3 	:	val_out <= 4'h4646;
         4'hecf8 	:	val_out <= 4'h465c;
         4'hecf9 	:	val_out <= 4'h465c;
         4'hecfa 	:	val_out <= 4'h465c;
         4'hecfb 	:	val_out <= 4'h465c;
         4'hed00 	:	val_out <= 4'h4673;
         4'hed01 	:	val_out <= 4'h4673;
         4'hed02 	:	val_out <= 4'h4673;
         4'hed03 	:	val_out <= 4'h4673;
         4'hed08 	:	val_out <= 4'h4689;
         4'hed09 	:	val_out <= 4'h4689;
         4'hed0a 	:	val_out <= 4'h4689;
         4'hed0b 	:	val_out <= 4'h4689;
         4'hed10 	:	val_out <= 4'h46a0;
         4'hed11 	:	val_out <= 4'h46a0;
         4'hed12 	:	val_out <= 4'h46a0;
         4'hed13 	:	val_out <= 4'h46a0;
         4'hed18 	:	val_out <= 4'h46b6;
         4'hed19 	:	val_out <= 4'h46b6;
         4'hed1a 	:	val_out <= 4'h46b6;
         4'hed1b 	:	val_out <= 4'h46b6;
         4'hed20 	:	val_out <= 4'h46cd;
         4'hed21 	:	val_out <= 4'h46cd;
         4'hed22 	:	val_out <= 4'h46cd;
         4'hed23 	:	val_out <= 4'h46cd;
         4'hed28 	:	val_out <= 4'h46e3;
         4'hed29 	:	val_out <= 4'h46e3;
         4'hed2a 	:	val_out <= 4'h46e3;
         4'hed2b 	:	val_out <= 4'h46e3;
         4'hed30 	:	val_out <= 4'h46f9;
         4'hed31 	:	val_out <= 4'h46f9;
         4'hed32 	:	val_out <= 4'h46f9;
         4'hed33 	:	val_out <= 4'h46f9;
         4'hed38 	:	val_out <= 4'h4710;
         4'hed39 	:	val_out <= 4'h4710;
         4'hed3a 	:	val_out <= 4'h4710;
         4'hed3b 	:	val_out <= 4'h4710;
         4'hed40 	:	val_out <= 4'h4727;
         4'hed41 	:	val_out <= 4'h4727;
         4'hed42 	:	val_out <= 4'h4727;
         4'hed43 	:	val_out <= 4'h4727;
         4'hed48 	:	val_out <= 4'h473d;
         4'hed49 	:	val_out <= 4'h473d;
         4'hed4a 	:	val_out <= 4'h473d;
         4'hed4b 	:	val_out <= 4'h473d;
         4'hed50 	:	val_out <= 4'h4754;
         4'hed51 	:	val_out <= 4'h4754;
         4'hed52 	:	val_out <= 4'h4754;
         4'hed53 	:	val_out <= 4'h4754;
         4'hed58 	:	val_out <= 4'h476a;
         4'hed59 	:	val_out <= 4'h476a;
         4'hed5a 	:	val_out <= 4'h476a;
         4'hed5b 	:	val_out <= 4'h476a;
         4'hed60 	:	val_out <= 4'h4781;
         4'hed61 	:	val_out <= 4'h4781;
         4'hed62 	:	val_out <= 4'h4781;
         4'hed63 	:	val_out <= 4'h4781;
         4'hed68 	:	val_out <= 4'h4797;
         4'hed69 	:	val_out <= 4'h4797;
         4'hed6a 	:	val_out <= 4'h4797;
         4'hed6b 	:	val_out <= 4'h4797;
         4'hed70 	:	val_out <= 4'h47ae;
         4'hed71 	:	val_out <= 4'h47ae;
         4'hed72 	:	val_out <= 4'h47ae;
         4'hed73 	:	val_out <= 4'h47ae;
         4'hed78 	:	val_out <= 4'h47c4;
         4'hed79 	:	val_out <= 4'h47c4;
         4'hed7a 	:	val_out <= 4'h47c4;
         4'hed7b 	:	val_out <= 4'h47c4;
         4'hed80 	:	val_out <= 4'h47db;
         4'hed81 	:	val_out <= 4'h47db;
         4'hed82 	:	val_out <= 4'h47db;
         4'hed83 	:	val_out <= 4'h47db;
         4'hed88 	:	val_out <= 4'h47f2;
         4'hed89 	:	val_out <= 4'h47f2;
         4'hed8a 	:	val_out <= 4'h47f2;
         4'hed8b 	:	val_out <= 4'h47f2;
         4'hed90 	:	val_out <= 4'h4808;
         4'hed91 	:	val_out <= 4'h4808;
         4'hed92 	:	val_out <= 4'h4808;
         4'hed93 	:	val_out <= 4'h4808;
         4'hed98 	:	val_out <= 4'h481f;
         4'hed99 	:	val_out <= 4'h481f;
         4'hed9a 	:	val_out <= 4'h481f;
         4'hed9b 	:	val_out <= 4'h481f;
         4'heda0 	:	val_out <= 4'h4835;
         4'heda1 	:	val_out <= 4'h4835;
         4'heda2 	:	val_out <= 4'h4835;
         4'heda3 	:	val_out <= 4'h4835;
         4'heda8 	:	val_out <= 4'h484c;
         4'heda9 	:	val_out <= 4'h484c;
         4'hedaa 	:	val_out <= 4'h484c;
         4'hedab 	:	val_out <= 4'h484c;
         4'hedb0 	:	val_out <= 4'h4863;
         4'hedb1 	:	val_out <= 4'h4863;
         4'hedb2 	:	val_out <= 4'h4863;
         4'hedb3 	:	val_out <= 4'h4863;
         4'hedb8 	:	val_out <= 4'h4879;
         4'hedb9 	:	val_out <= 4'h4879;
         4'hedba 	:	val_out <= 4'h4879;
         4'hedbb 	:	val_out <= 4'h4879;
         4'hedc0 	:	val_out <= 4'h4890;
         4'hedc1 	:	val_out <= 4'h4890;
         4'hedc2 	:	val_out <= 4'h4890;
         4'hedc3 	:	val_out <= 4'h4890;
         4'hedc8 	:	val_out <= 4'h48a7;
         4'hedc9 	:	val_out <= 4'h48a7;
         4'hedca 	:	val_out <= 4'h48a7;
         4'hedcb 	:	val_out <= 4'h48a7;
         4'hedd0 	:	val_out <= 4'h48bd;
         4'hedd1 	:	val_out <= 4'h48bd;
         4'hedd2 	:	val_out <= 4'h48bd;
         4'hedd3 	:	val_out <= 4'h48bd;
         4'hedd8 	:	val_out <= 4'h48d4;
         4'hedd9 	:	val_out <= 4'h48d4;
         4'hedda 	:	val_out <= 4'h48d4;
         4'heddb 	:	val_out <= 4'h48d4;
         4'hede0 	:	val_out <= 4'h48eb;
         4'hede1 	:	val_out <= 4'h48eb;
         4'hede2 	:	val_out <= 4'h48eb;
         4'hede3 	:	val_out <= 4'h48eb;
         4'hede8 	:	val_out <= 4'h4901;
         4'hede9 	:	val_out <= 4'h4901;
         4'hedea 	:	val_out <= 4'h4901;
         4'hedeb 	:	val_out <= 4'h4901;
         4'hedf0 	:	val_out <= 4'h4918;
         4'hedf1 	:	val_out <= 4'h4918;
         4'hedf2 	:	val_out <= 4'h4918;
         4'hedf3 	:	val_out <= 4'h4918;
         4'hedf8 	:	val_out <= 4'h492f;
         4'hedf9 	:	val_out <= 4'h492f;
         4'hedfa 	:	val_out <= 4'h492f;
         4'hedfb 	:	val_out <= 4'h492f;
         4'hee00 	:	val_out <= 4'h4945;
         4'hee01 	:	val_out <= 4'h4945;
         4'hee02 	:	val_out <= 4'h4945;
         4'hee03 	:	val_out <= 4'h4945;
         4'hee08 	:	val_out <= 4'h495c;
         4'hee09 	:	val_out <= 4'h495c;
         4'hee0a 	:	val_out <= 4'h495c;
         4'hee0b 	:	val_out <= 4'h495c;
         4'hee10 	:	val_out <= 4'h4973;
         4'hee11 	:	val_out <= 4'h4973;
         4'hee12 	:	val_out <= 4'h4973;
         4'hee13 	:	val_out <= 4'h4973;
         4'hee18 	:	val_out <= 4'h498a;
         4'hee19 	:	val_out <= 4'h498a;
         4'hee1a 	:	val_out <= 4'h498a;
         4'hee1b 	:	val_out <= 4'h498a;
         4'hee20 	:	val_out <= 4'h49a0;
         4'hee21 	:	val_out <= 4'h49a0;
         4'hee22 	:	val_out <= 4'h49a0;
         4'hee23 	:	val_out <= 4'h49a0;
         4'hee28 	:	val_out <= 4'h49b7;
         4'hee29 	:	val_out <= 4'h49b7;
         4'hee2a 	:	val_out <= 4'h49b7;
         4'hee2b 	:	val_out <= 4'h49b7;
         4'hee30 	:	val_out <= 4'h49ce;
         4'hee31 	:	val_out <= 4'h49ce;
         4'hee32 	:	val_out <= 4'h49ce;
         4'hee33 	:	val_out <= 4'h49ce;
         4'hee38 	:	val_out <= 4'h49e5;
         4'hee39 	:	val_out <= 4'h49e5;
         4'hee3a 	:	val_out <= 4'h49e5;
         4'hee3b 	:	val_out <= 4'h49e5;
         4'hee40 	:	val_out <= 4'h49fb;
         4'hee41 	:	val_out <= 4'h49fb;
         4'hee42 	:	val_out <= 4'h49fb;
         4'hee43 	:	val_out <= 4'h49fb;
         4'hee48 	:	val_out <= 4'h4a12;
         4'hee49 	:	val_out <= 4'h4a12;
         4'hee4a 	:	val_out <= 4'h4a12;
         4'hee4b 	:	val_out <= 4'h4a12;
         4'hee50 	:	val_out <= 4'h4a29;
         4'hee51 	:	val_out <= 4'h4a29;
         4'hee52 	:	val_out <= 4'h4a29;
         4'hee53 	:	val_out <= 4'h4a29;
         4'hee58 	:	val_out <= 4'h4a40;
         4'hee59 	:	val_out <= 4'h4a40;
         4'hee5a 	:	val_out <= 4'h4a40;
         4'hee5b 	:	val_out <= 4'h4a40;
         4'hee60 	:	val_out <= 4'h4a57;
         4'hee61 	:	val_out <= 4'h4a57;
         4'hee62 	:	val_out <= 4'h4a57;
         4'hee63 	:	val_out <= 4'h4a57;
         4'hee68 	:	val_out <= 4'h4a6d;
         4'hee69 	:	val_out <= 4'h4a6d;
         4'hee6a 	:	val_out <= 4'h4a6d;
         4'hee6b 	:	val_out <= 4'h4a6d;
         4'hee70 	:	val_out <= 4'h4a84;
         4'hee71 	:	val_out <= 4'h4a84;
         4'hee72 	:	val_out <= 4'h4a84;
         4'hee73 	:	val_out <= 4'h4a84;
         4'hee78 	:	val_out <= 4'h4a9b;
         4'hee79 	:	val_out <= 4'h4a9b;
         4'hee7a 	:	val_out <= 4'h4a9b;
         4'hee7b 	:	val_out <= 4'h4a9b;
         4'hee80 	:	val_out <= 4'h4ab2;
         4'hee81 	:	val_out <= 4'h4ab2;
         4'hee82 	:	val_out <= 4'h4ab2;
         4'hee83 	:	val_out <= 4'h4ab2;
         4'hee88 	:	val_out <= 4'h4ac9;
         4'hee89 	:	val_out <= 4'h4ac9;
         4'hee8a 	:	val_out <= 4'h4ac9;
         4'hee8b 	:	val_out <= 4'h4ac9;
         4'hee90 	:	val_out <= 4'h4ae0;
         4'hee91 	:	val_out <= 4'h4ae0;
         4'hee92 	:	val_out <= 4'h4ae0;
         4'hee93 	:	val_out <= 4'h4ae0;
         4'hee98 	:	val_out <= 4'h4af7;
         4'hee99 	:	val_out <= 4'h4af7;
         4'hee9a 	:	val_out <= 4'h4af7;
         4'hee9b 	:	val_out <= 4'h4af7;
         4'heea0 	:	val_out <= 4'h4b0d;
         4'heea1 	:	val_out <= 4'h4b0d;
         4'heea2 	:	val_out <= 4'h4b0d;
         4'heea3 	:	val_out <= 4'h4b0d;
         4'heea8 	:	val_out <= 4'h4b24;
         4'heea9 	:	val_out <= 4'h4b24;
         4'heeaa 	:	val_out <= 4'h4b24;
         4'heeab 	:	val_out <= 4'h4b24;
         4'heeb0 	:	val_out <= 4'h4b3b;
         4'heeb1 	:	val_out <= 4'h4b3b;
         4'heeb2 	:	val_out <= 4'h4b3b;
         4'heeb3 	:	val_out <= 4'h4b3b;
         4'heeb8 	:	val_out <= 4'h4b52;
         4'heeb9 	:	val_out <= 4'h4b52;
         4'heeba 	:	val_out <= 4'h4b52;
         4'heebb 	:	val_out <= 4'h4b52;
         4'heec0 	:	val_out <= 4'h4b69;
         4'heec1 	:	val_out <= 4'h4b69;
         4'heec2 	:	val_out <= 4'h4b69;
         4'heec3 	:	val_out <= 4'h4b69;
         4'heec8 	:	val_out <= 4'h4b80;
         4'heec9 	:	val_out <= 4'h4b80;
         4'heeca 	:	val_out <= 4'h4b80;
         4'heecb 	:	val_out <= 4'h4b80;
         4'heed0 	:	val_out <= 4'h4b97;
         4'heed1 	:	val_out <= 4'h4b97;
         4'heed2 	:	val_out <= 4'h4b97;
         4'heed3 	:	val_out <= 4'h4b97;
         4'heed8 	:	val_out <= 4'h4bae;
         4'heed9 	:	val_out <= 4'h4bae;
         4'heeda 	:	val_out <= 4'h4bae;
         4'heedb 	:	val_out <= 4'h4bae;
         4'heee0 	:	val_out <= 4'h4bc5;
         4'heee1 	:	val_out <= 4'h4bc5;
         4'heee2 	:	val_out <= 4'h4bc5;
         4'heee3 	:	val_out <= 4'h4bc5;
         4'heee8 	:	val_out <= 4'h4bdc;
         4'heee9 	:	val_out <= 4'h4bdc;
         4'heeea 	:	val_out <= 4'h4bdc;
         4'heeeb 	:	val_out <= 4'h4bdc;
         4'heef0 	:	val_out <= 4'h4bf3;
         4'heef1 	:	val_out <= 4'h4bf3;
         4'heef2 	:	val_out <= 4'h4bf3;
         4'heef3 	:	val_out <= 4'h4bf3;
         4'heef8 	:	val_out <= 4'h4c0a;
         4'heef9 	:	val_out <= 4'h4c0a;
         4'heefa 	:	val_out <= 4'h4c0a;
         4'heefb 	:	val_out <= 4'h4c0a;
         4'hef00 	:	val_out <= 4'h4c21;
         4'hef01 	:	val_out <= 4'h4c21;
         4'hef02 	:	val_out <= 4'h4c21;
         4'hef03 	:	val_out <= 4'h4c21;
         4'hef08 	:	val_out <= 4'h4c38;
         4'hef09 	:	val_out <= 4'h4c38;
         4'hef0a 	:	val_out <= 4'h4c38;
         4'hef0b 	:	val_out <= 4'h4c38;
         4'hef10 	:	val_out <= 4'h4c4f;
         4'hef11 	:	val_out <= 4'h4c4f;
         4'hef12 	:	val_out <= 4'h4c4f;
         4'hef13 	:	val_out <= 4'h4c4f;
         4'hef18 	:	val_out <= 4'h4c66;
         4'hef19 	:	val_out <= 4'h4c66;
         4'hef1a 	:	val_out <= 4'h4c66;
         4'hef1b 	:	val_out <= 4'h4c66;
         4'hef20 	:	val_out <= 4'h4c7d;
         4'hef21 	:	val_out <= 4'h4c7d;
         4'hef22 	:	val_out <= 4'h4c7d;
         4'hef23 	:	val_out <= 4'h4c7d;
         4'hef28 	:	val_out <= 4'h4c94;
         4'hef29 	:	val_out <= 4'h4c94;
         4'hef2a 	:	val_out <= 4'h4c94;
         4'hef2b 	:	val_out <= 4'h4c94;
         4'hef30 	:	val_out <= 4'h4cab;
         4'hef31 	:	val_out <= 4'h4cab;
         4'hef32 	:	val_out <= 4'h4cab;
         4'hef33 	:	val_out <= 4'h4cab;
         4'hef38 	:	val_out <= 4'h4cc2;
         4'hef39 	:	val_out <= 4'h4cc2;
         4'hef3a 	:	val_out <= 4'h4cc2;
         4'hef3b 	:	val_out <= 4'h4cc2;
         4'hef40 	:	val_out <= 4'h4cd9;
         4'hef41 	:	val_out <= 4'h4cd9;
         4'hef42 	:	val_out <= 4'h4cd9;
         4'hef43 	:	val_out <= 4'h4cd9;
         4'hef48 	:	val_out <= 4'h4cf0;
         4'hef49 	:	val_out <= 4'h4cf0;
         4'hef4a 	:	val_out <= 4'h4cf0;
         4'hef4b 	:	val_out <= 4'h4cf0;
         4'hef50 	:	val_out <= 4'h4d07;
         4'hef51 	:	val_out <= 4'h4d07;
         4'hef52 	:	val_out <= 4'h4d07;
         4'hef53 	:	val_out <= 4'h4d07;
         4'hef58 	:	val_out <= 4'h4d1e;
         4'hef59 	:	val_out <= 4'h4d1e;
         4'hef5a 	:	val_out <= 4'h4d1e;
         4'hef5b 	:	val_out <= 4'h4d1e;
         4'hef60 	:	val_out <= 4'h4d35;
         4'hef61 	:	val_out <= 4'h4d35;
         4'hef62 	:	val_out <= 4'h4d35;
         4'hef63 	:	val_out <= 4'h4d35;
         4'hef68 	:	val_out <= 4'h4d4c;
         4'hef69 	:	val_out <= 4'h4d4c;
         4'hef6a 	:	val_out <= 4'h4d4c;
         4'hef6b 	:	val_out <= 4'h4d4c;
         4'hef70 	:	val_out <= 4'h4d63;
         4'hef71 	:	val_out <= 4'h4d63;
         4'hef72 	:	val_out <= 4'h4d63;
         4'hef73 	:	val_out <= 4'h4d63;
         4'hef78 	:	val_out <= 4'h4d7a;
         4'hef79 	:	val_out <= 4'h4d7a;
         4'hef7a 	:	val_out <= 4'h4d7a;
         4'hef7b 	:	val_out <= 4'h4d7a;
         4'hef80 	:	val_out <= 4'h4d91;
         4'hef81 	:	val_out <= 4'h4d91;
         4'hef82 	:	val_out <= 4'h4d91;
         4'hef83 	:	val_out <= 4'h4d91;
         4'hef88 	:	val_out <= 4'h4da8;
         4'hef89 	:	val_out <= 4'h4da8;
         4'hef8a 	:	val_out <= 4'h4da8;
         4'hef8b 	:	val_out <= 4'h4da8;
         4'hef90 	:	val_out <= 4'h4dbf;
         4'hef91 	:	val_out <= 4'h4dbf;
         4'hef92 	:	val_out <= 4'h4dbf;
         4'hef93 	:	val_out <= 4'h4dbf;
         4'hef98 	:	val_out <= 4'h4dd7;
         4'hef99 	:	val_out <= 4'h4dd7;
         4'hef9a 	:	val_out <= 4'h4dd7;
         4'hef9b 	:	val_out <= 4'h4dd7;
         4'hefa0 	:	val_out <= 4'h4dee;
         4'hefa1 	:	val_out <= 4'h4dee;
         4'hefa2 	:	val_out <= 4'h4dee;
         4'hefa3 	:	val_out <= 4'h4dee;
         4'hefa8 	:	val_out <= 4'h4e05;
         4'hefa9 	:	val_out <= 4'h4e05;
         4'hefaa 	:	val_out <= 4'h4e05;
         4'hefab 	:	val_out <= 4'h4e05;
         4'hefb0 	:	val_out <= 4'h4e1c;
         4'hefb1 	:	val_out <= 4'h4e1c;
         4'hefb2 	:	val_out <= 4'h4e1c;
         4'hefb3 	:	val_out <= 4'h4e1c;
         4'hefb8 	:	val_out <= 4'h4e33;
         4'hefb9 	:	val_out <= 4'h4e33;
         4'hefba 	:	val_out <= 4'h4e33;
         4'hefbb 	:	val_out <= 4'h4e33;
         4'hefc0 	:	val_out <= 4'h4e4a;
         4'hefc1 	:	val_out <= 4'h4e4a;
         4'hefc2 	:	val_out <= 4'h4e4a;
         4'hefc3 	:	val_out <= 4'h4e4a;
         4'hefc8 	:	val_out <= 4'h4e61;
         4'hefc9 	:	val_out <= 4'h4e61;
         4'hefca 	:	val_out <= 4'h4e61;
         4'hefcb 	:	val_out <= 4'h4e61;
         4'hefd0 	:	val_out <= 4'h4e79;
         4'hefd1 	:	val_out <= 4'h4e79;
         4'hefd2 	:	val_out <= 4'h4e79;
         4'hefd3 	:	val_out <= 4'h4e79;
         4'hefd8 	:	val_out <= 4'h4e90;
         4'hefd9 	:	val_out <= 4'h4e90;
         4'hefda 	:	val_out <= 4'h4e90;
         4'hefdb 	:	val_out <= 4'h4e90;
         4'hefe0 	:	val_out <= 4'h4ea7;
         4'hefe1 	:	val_out <= 4'h4ea7;
         4'hefe2 	:	val_out <= 4'h4ea7;
         4'hefe3 	:	val_out <= 4'h4ea7;
         4'hefe8 	:	val_out <= 4'h4ebe;
         4'hefe9 	:	val_out <= 4'h4ebe;
         4'hefea 	:	val_out <= 4'h4ebe;
         4'hefeb 	:	val_out <= 4'h4ebe;
         4'heff0 	:	val_out <= 4'h4ed5;
         4'heff1 	:	val_out <= 4'h4ed5;
         4'heff2 	:	val_out <= 4'h4ed5;
         4'heff3 	:	val_out <= 4'h4ed5;
         4'heff8 	:	val_out <= 4'h4eed;
         4'heff9 	:	val_out <= 4'h4eed;
         4'heffa 	:	val_out <= 4'h4eed;
         4'heffb 	:	val_out <= 4'h4eed;
         4'hf000 	:	val_out <= 4'h4f04;
         4'hf001 	:	val_out <= 4'h4f04;
         4'hf002 	:	val_out <= 4'h4f04;
         4'hf003 	:	val_out <= 4'h4f04;
         4'hf008 	:	val_out <= 4'h4f1b;
         4'hf009 	:	val_out <= 4'h4f1b;
         4'hf00a 	:	val_out <= 4'h4f1b;
         4'hf00b 	:	val_out <= 4'h4f1b;
         4'hf010 	:	val_out <= 4'h4f32;
         4'hf011 	:	val_out <= 4'h4f32;
         4'hf012 	:	val_out <= 4'h4f32;
         4'hf013 	:	val_out <= 4'h4f32;
         4'hf018 	:	val_out <= 4'h4f49;
         4'hf019 	:	val_out <= 4'h4f49;
         4'hf01a 	:	val_out <= 4'h4f49;
         4'hf01b 	:	val_out <= 4'h4f49;
         4'hf020 	:	val_out <= 4'h4f61;
         4'hf021 	:	val_out <= 4'h4f61;
         4'hf022 	:	val_out <= 4'h4f61;
         4'hf023 	:	val_out <= 4'h4f61;
         4'hf028 	:	val_out <= 4'h4f78;
         4'hf029 	:	val_out <= 4'h4f78;
         4'hf02a 	:	val_out <= 4'h4f78;
         4'hf02b 	:	val_out <= 4'h4f78;
         4'hf030 	:	val_out <= 4'h4f8f;
         4'hf031 	:	val_out <= 4'h4f8f;
         4'hf032 	:	val_out <= 4'h4f8f;
         4'hf033 	:	val_out <= 4'h4f8f;
         4'hf038 	:	val_out <= 4'h4fa6;
         4'hf039 	:	val_out <= 4'h4fa6;
         4'hf03a 	:	val_out <= 4'h4fa6;
         4'hf03b 	:	val_out <= 4'h4fa6;
         4'hf040 	:	val_out <= 4'h4fbe;
         4'hf041 	:	val_out <= 4'h4fbe;
         4'hf042 	:	val_out <= 4'h4fbe;
         4'hf043 	:	val_out <= 4'h4fbe;
         4'hf048 	:	val_out <= 4'h4fd5;
         4'hf049 	:	val_out <= 4'h4fd5;
         4'hf04a 	:	val_out <= 4'h4fd5;
         4'hf04b 	:	val_out <= 4'h4fd5;
         4'hf050 	:	val_out <= 4'h4fec;
         4'hf051 	:	val_out <= 4'h4fec;
         4'hf052 	:	val_out <= 4'h4fec;
         4'hf053 	:	val_out <= 4'h4fec;
         4'hf058 	:	val_out <= 4'h5004;
         4'hf059 	:	val_out <= 4'h5004;
         4'hf05a 	:	val_out <= 4'h5004;
         4'hf05b 	:	val_out <= 4'h5004;
         4'hf060 	:	val_out <= 4'h501b;
         4'hf061 	:	val_out <= 4'h501b;
         4'hf062 	:	val_out <= 4'h501b;
         4'hf063 	:	val_out <= 4'h501b;
         4'hf068 	:	val_out <= 4'h5032;
         4'hf069 	:	val_out <= 4'h5032;
         4'hf06a 	:	val_out <= 4'h5032;
         4'hf06b 	:	val_out <= 4'h5032;
         4'hf070 	:	val_out <= 4'h504a;
         4'hf071 	:	val_out <= 4'h504a;
         4'hf072 	:	val_out <= 4'h504a;
         4'hf073 	:	val_out <= 4'h504a;
         4'hf078 	:	val_out <= 4'h5061;
         4'hf079 	:	val_out <= 4'h5061;
         4'hf07a 	:	val_out <= 4'h5061;
         4'hf07b 	:	val_out <= 4'h5061;
         4'hf080 	:	val_out <= 4'h5078;
         4'hf081 	:	val_out <= 4'h5078;
         4'hf082 	:	val_out <= 4'h5078;
         4'hf083 	:	val_out <= 4'h5078;
         4'hf088 	:	val_out <= 4'h5090;
         4'hf089 	:	val_out <= 4'h5090;
         4'hf08a 	:	val_out <= 4'h5090;
         4'hf08b 	:	val_out <= 4'h5090;
         4'hf090 	:	val_out <= 4'h50a7;
         4'hf091 	:	val_out <= 4'h50a7;
         4'hf092 	:	val_out <= 4'h50a7;
         4'hf093 	:	val_out <= 4'h50a7;
         4'hf098 	:	val_out <= 4'h50be;
         4'hf099 	:	val_out <= 4'h50be;
         4'hf09a 	:	val_out <= 4'h50be;
         4'hf09b 	:	val_out <= 4'h50be;
         4'hf0a0 	:	val_out <= 4'h50d6;
         4'hf0a1 	:	val_out <= 4'h50d6;
         4'hf0a2 	:	val_out <= 4'h50d6;
         4'hf0a3 	:	val_out <= 4'h50d6;
         4'hf0a8 	:	val_out <= 4'h50ed;
         4'hf0a9 	:	val_out <= 4'h50ed;
         4'hf0aa 	:	val_out <= 4'h50ed;
         4'hf0ab 	:	val_out <= 4'h50ed;
         4'hf0b0 	:	val_out <= 4'h5104;
         4'hf0b1 	:	val_out <= 4'h5104;
         4'hf0b2 	:	val_out <= 4'h5104;
         4'hf0b3 	:	val_out <= 4'h5104;
         4'hf0b8 	:	val_out <= 4'h511c;
         4'hf0b9 	:	val_out <= 4'h511c;
         4'hf0ba 	:	val_out <= 4'h511c;
         4'hf0bb 	:	val_out <= 4'h511c;
         4'hf0c0 	:	val_out <= 4'h5133;
         4'hf0c1 	:	val_out <= 4'h5133;
         4'hf0c2 	:	val_out <= 4'h5133;
         4'hf0c3 	:	val_out <= 4'h5133;
         4'hf0c8 	:	val_out <= 4'h514a;
         4'hf0c9 	:	val_out <= 4'h514a;
         4'hf0ca 	:	val_out <= 4'h514a;
         4'hf0cb 	:	val_out <= 4'h514a;
         4'hf0d0 	:	val_out <= 4'h5162;
         4'hf0d1 	:	val_out <= 4'h5162;
         4'hf0d2 	:	val_out <= 4'h5162;
         4'hf0d3 	:	val_out <= 4'h5162;
         4'hf0d8 	:	val_out <= 4'h5179;
         4'hf0d9 	:	val_out <= 4'h5179;
         4'hf0da 	:	val_out <= 4'h5179;
         4'hf0db 	:	val_out <= 4'h5179;
         4'hf0e0 	:	val_out <= 4'h5191;
         4'hf0e1 	:	val_out <= 4'h5191;
         4'hf0e2 	:	val_out <= 4'h5191;
         4'hf0e3 	:	val_out <= 4'h5191;
         4'hf0e8 	:	val_out <= 4'h51a8;
         4'hf0e9 	:	val_out <= 4'h51a8;
         4'hf0ea 	:	val_out <= 4'h51a8;
         4'hf0eb 	:	val_out <= 4'h51a8;
         4'hf0f0 	:	val_out <= 4'h51c0;
         4'hf0f1 	:	val_out <= 4'h51c0;
         4'hf0f2 	:	val_out <= 4'h51c0;
         4'hf0f3 	:	val_out <= 4'h51c0;
         4'hf0f8 	:	val_out <= 4'h51d7;
         4'hf0f9 	:	val_out <= 4'h51d7;
         4'hf0fa 	:	val_out <= 4'h51d7;
         4'hf0fb 	:	val_out <= 4'h51d7;
         4'hf100 	:	val_out <= 4'h51ee;
         4'hf101 	:	val_out <= 4'h51ee;
         4'hf102 	:	val_out <= 4'h51ee;
         4'hf103 	:	val_out <= 4'h51ee;
         4'hf108 	:	val_out <= 4'h5206;
         4'hf109 	:	val_out <= 4'h5206;
         4'hf10a 	:	val_out <= 4'h5206;
         4'hf10b 	:	val_out <= 4'h5206;
         4'hf110 	:	val_out <= 4'h521d;
         4'hf111 	:	val_out <= 4'h521d;
         4'hf112 	:	val_out <= 4'h521d;
         4'hf113 	:	val_out <= 4'h521d;
         4'hf118 	:	val_out <= 4'h5235;
         4'hf119 	:	val_out <= 4'h5235;
         4'hf11a 	:	val_out <= 4'h5235;
         4'hf11b 	:	val_out <= 4'h5235;
         4'hf120 	:	val_out <= 4'h524c;
         4'hf121 	:	val_out <= 4'h524c;
         4'hf122 	:	val_out <= 4'h524c;
         4'hf123 	:	val_out <= 4'h524c;
         4'hf128 	:	val_out <= 4'h5264;
         4'hf129 	:	val_out <= 4'h5264;
         4'hf12a 	:	val_out <= 4'h5264;
         4'hf12b 	:	val_out <= 4'h5264;
         4'hf130 	:	val_out <= 4'h527b;
         4'hf131 	:	val_out <= 4'h527b;
         4'hf132 	:	val_out <= 4'h527b;
         4'hf133 	:	val_out <= 4'h527b;
         4'hf138 	:	val_out <= 4'h5293;
         4'hf139 	:	val_out <= 4'h5293;
         4'hf13a 	:	val_out <= 4'h5293;
         4'hf13b 	:	val_out <= 4'h5293;
         4'hf140 	:	val_out <= 4'h52aa;
         4'hf141 	:	val_out <= 4'h52aa;
         4'hf142 	:	val_out <= 4'h52aa;
         4'hf143 	:	val_out <= 4'h52aa;
         4'hf148 	:	val_out <= 4'h52c2;
         4'hf149 	:	val_out <= 4'h52c2;
         4'hf14a 	:	val_out <= 4'h52c2;
         4'hf14b 	:	val_out <= 4'h52c2;
         4'hf150 	:	val_out <= 4'h52d9;
         4'hf151 	:	val_out <= 4'h52d9;
         4'hf152 	:	val_out <= 4'h52d9;
         4'hf153 	:	val_out <= 4'h52d9;
         4'hf158 	:	val_out <= 4'h52f1;
         4'hf159 	:	val_out <= 4'h52f1;
         4'hf15a 	:	val_out <= 4'h52f1;
         4'hf15b 	:	val_out <= 4'h52f1;
         4'hf160 	:	val_out <= 4'h5308;
         4'hf161 	:	val_out <= 4'h5308;
         4'hf162 	:	val_out <= 4'h5308;
         4'hf163 	:	val_out <= 4'h5308;
         4'hf168 	:	val_out <= 4'h5320;
         4'hf169 	:	val_out <= 4'h5320;
         4'hf16a 	:	val_out <= 4'h5320;
         4'hf16b 	:	val_out <= 4'h5320;
         4'hf170 	:	val_out <= 4'h5337;
         4'hf171 	:	val_out <= 4'h5337;
         4'hf172 	:	val_out <= 4'h5337;
         4'hf173 	:	val_out <= 4'h5337;
         4'hf178 	:	val_out <= 4'h534f;
         4'hf179 	:	val_out <= 4'h534f;
         4'hf17a 	:	val_out <= 4'h534f;
         4'hf17b 	:	val_out <= 4'h534f;
         4'hf180 	:	val_out <= 4'h5367;
         4'hf181 	:	val_out <= 4'h5367;
         4'hf182 	:	val_out <= 4'h5367;
         4'hf183 	:	val_out <= 4'h5367;
         4'hf188 	:	val_out <= 4'h537e;
         4'hf189 	:	val_out <= 4'h537e;
         4'hf18a 	:	val_out <= 4'h537e;
         4'hf18b 	:	val_out <= 4'h537e;
         4'hf190 	:	val_out <= 4'h5396;
         4'hf191 	:	val_out <= 4'h5396;
         4'hf192 	:	val_out <= 4'h5396;
         4'hf193 	:	val_out <= 4'h5396;
         4'hf198 	:	val_out <= 4'h53ad;
         4'hf199 	:	val_out <= 4'h53ad;
         4'hf19a 	:	val_out <= 4'h53ad;
         4'hf19b 	:	val_out <= 4'h53ad;
         4'hf1a0 	:	val_out <= 4'h53c5;
         4'hf1a1 	:	val_out <= 4'h53c5;
         4'hf1a2 	:	val_out <= 4'h53c5;
         4'hf1a3 	:	val_out <= 4'h53c5;
         4'hf1a8 	:	val_out <= 4'h53dc;
         4'hf1a9 	:	val_out <= 4'h53dc;
         4'hf1aa 	:	val_out <= 4'h53dc;
         4'hf1ab 	:	val_out <= 4'h53dc;
         4'hf1b0 	:	val_out <= 4'h53f4;
         4'hf1b1 	:	val_out <= 4'h53f4;
         4'hf1b2 	:	val_out <= 4'h53f4;
         4'hf1b3 	:	val_out <= 4'h53f4;
         4'hf1b8 	:	val_out <= 4'h540c;
         4'hf1b9 	:	val_out <= 4'h540c;
         4'hf1ba 	:	val_out <= 4'h540c;
         4'hf1bb 	:	val_out <= 4'h540c;
         4'hf1c0 	:	val_out <= 4'h5423;
         4'hf1c1 	:	val_out <= 4'h5423;
         4'hf1c2 	:	val_out <= 4'h5423;
         4'hf1c3 	:	val_out <= 4'h5423;
         4'hf1c8 	:	val_out <= 4'h543b;
         4'hf1c9 	:	val_out <= 4'h543b;
         4'hf1ca 	:	val_out <= 4'h543b;
         4'hf1cb 	:	val_out <= 4'h543b;
         4'hf1d0 	:	val_out <= 4'h5452;
         4'hf1d1 	:	val_out <= 4'h5452;
         4'hf1d2 	:	val_out <= 4'h5452;
         4'hf1d3 	:	val_out <= 4'h5452;
         4'hf1d8 	:	val_out <= 4'h546a;
         4'hf1d9 	:	val_out <= 4'h546a;
         4'hf1da 	:	val_out <= 4'h546a;
         4'hf1db 	:	val_out <= 4'h546a;
         4'hf1e0 	:	val_out <= 4'h5482;
         4'hf1e1 	:	val_out <= 4'h5482;
         4'hf1e2 	:	val_out <= 4'h5482;
         4'hf1e3 	:	val_out <= 4'h5482;
         4'hf1e8 	:	val_out <= 4'h5499;
         4'hf1e9 	:	val_out <= 4'h5499;
         4'hf1ea 	:	val_out <= 4'h5499;
         4'hf1eb 	:	val_out <= 4'h5499;
         4'hf1f0 	:	val_out <= 4'h54b1;
         4'hf1f1 	:	val_out <= 4'h54b1;
         4'hf1f2 	:	val_out <= 4'h54b1;
         4'hf1f3 	:	val_out <= 4'h54b1;
         4'hf1f8 	:	val_out <= 4'h54c9;
         4'hf1f9 	:	val_out <= 4'h54c9;
         4'hf1fa 	:	val_out <= 4'h54c9;
         4'hf1fb 	:	val_out <= 4'h54c9;
         4'hf200 	:	val_out <= 4'h54e0;
         4'hf201 	:	val_out <= 4'h54e0;
         4'hf202 	:	val_out <= 4'h54e0;
         4'hf203 	:	val_out <= 4'h54e0;
         4'hf208 	:	val_out <= 4'h54f8;
         4'hf209 	:	val_out <= 4'h54f8;
         4'hf20a 	:	val_out <= 4'h54f8;
         4'hf20b 	:	val_out <= 4'h54f8;
         4'hf210 	:	val_out <= 4'h5510;
         4'hf211 	:	val_out <= 4'h5510;
         4'hf212 	:	val_out <= 4'h5510;
         4'hf213 	:	val_out <= 4'h5510;
         4'hf218 	:	val_out <= 4'h5527;
         4'hf219 	:	val_out <= 4'h5527;
         4'hf21a 	:	val_out <= 4'h5527;
         4'hf21b 	:	val_out <= 4'h5527;
         4'hf220 	:	val_out <= 4'h553f;
         4'hf221 	:	val_out <= 4'h553f;
         4'hf222 	:	val_out <= 4'h553f;
         4'hf223 	:	val_out <= 4'h553f;
         4'hf228 	:	val_out <= 4'h5557;
         4'hf229 	:	val_out <= 4'h5557;
         4'hf22a 	:	val_out <= 4'h5557;
         4'hf22b 	:	val_out <= 4'h5557;
         4'hf230 	:	val_out <= 4'h556e;
         4'hf231 	:	val_out <= 4'h556e;
         4'hf232 	:	val_out <= 4'h556e;
         4'hf233 	:	val_out <= 4'h556e;
         4'hf238 	:	val_out <= 4'h5586;
         4'hf239 	:	val_out <= 4'h5586;
         4'hf23a 	:	val_out <= 4'h5586;
         4'hf23b 	:	val_out <= 4'h5586;
         4'hf240 	:	val_out <= 4'h559e;
         4'hf241 	:	val_out <= 4'h559e;
         4'hf242 	:	val_out <= 4'h559e;
         4'hf243 	:	val_out <= 4'h559e;
         4'hf248 	:	val_out <= 4'h55b6;
         4'hf249 	:	val_out <= 4'h55b6;
         4'hf24a 	:	val_out <= 4'h55b6;
         4'hf24b 	:	val_out <= 4'h55b6;
         4'hf250 	:	val_out <= 4'h55cd;
         4'hf251 	:	val_out <= 4'h55cd;
         4'hf252 	:	val_out <= 4'h55cd;
         4'hf253 	:	val_out <= 4'h55cd;
         4'hf258 	:	val_out <= 4'h55e5;
         4'hf259 	:	val_out <= 4'h55e5;
         4'hf25a 	:	val_out <= 4'h55e5;
         4'hf25b 	:	val_out <= 4'h55e5;
         4'hf260 	:	val_out <= 4'h55fd;
         4'hf261 	:	val_out <= 4'h55fd;
         4'hf262 	:	val_out <= 4'h55fd;
         4'hf263 	:	val_out <= 4'h55fd;
         4'hf268 	:	val_out <= 4'h5614;
         4'hf269 	:	val_out <= 4'h5614;
         4'hf26a 	:	val_out <= 4'h5614;
         4'hf26b 	:	val_out <= 4'h5614;
         4'hf270 	:	val_out <= 4'h562c;
         4'hf271 	:	val_out <= 4'h562c;
         4'hf272 	:	val_out <= 4'h562c;
         4'hf273 	:	val_out <= 4'h562c;
         4'hf278 	:	val_out <= 4'h5644;
         4'hf279 	:	val_out <= 4'h5644;
         4'hf27a 	:	val_out <= 4'h5644;
         4'hf27b 	:	val_out <= 4'h5644;
         4'hf280 	:	val_out <= 4'h565c;
         4'hf281 	:	val_out <= 4'h565c;
         4'hf282 	:	val_out <= 4'h565c;
         4'hf283 	:	val_out <= 4'h565c;
         4'hf288 	:	val_out <= 4'h5674;
         4'hf289 	:	val_out <= 4'h5674;
         4'hf28a 	:	val_out <= 4'h5674;
         4'hf28b 	:	val_out <= 4'h5674;
         4'hf290 	:	val_out <= 4'h568b;
         4'hf291 	:	val_out <= 4'h568b;
         4'hf292 	:	val_out <= 4'h568b;
         4'hf293 	:	val_out <= 4'h568b;
         4'hf298 	:	val_out <= 4'h56a3;
         4'hf299 	:	val_out <= 4'h56a3;
         4'hf29a 	:	val_out <= 4'h56a3;
         4'hf29b 	:	val_out <= 4'h56a3;
         4'hf2a0 	:	val_out <= 4'h56bb;
         4'hf2a1 	:	val_out <= 4'h56bb;
         4'hf2a2 	:	val_out <= 4'h56bb;
         4'hf2a3 	:	val_out <= 4'h56bb;
         4'hf2a8 	:	val_out <= 4'h56d3;
         4'hf2a9 	:	val_out <= 4'h56d3;
         4'hf2aa 	:	val_out <= 4'h56d3;
         4'hf2ab 	:	val_out <= 4'h56d3;
         4'hf2b0 	:	val_out <= 4'h56ea;
         4'hf2b1 	:	val_out <= 4'h56ea;
         4'hf2b2 	:	val_out <= 4'h56ea;
         4'hf2b3 	:	val_out <= 4'h56ea;
         4'hf2b8 	:	val_out <= 4'h5702;
         4'hf2b9 	:	val_out <= 4'h5702;
         4'hf2ba 	:	val_out <= 4'h5702;
         4'hf2bb 	:	val_out <= 4'h5702;
         4'hf2c0 	:	val_out <= 4'h571a;
         4'hf2c1 	:	val_out <= 4'h571a;
         4'hf2c2 	:	val_out <= 4'h571a;
         4'hf2c3 	:	val_out <= 4'h571a;
         4'hf2c8 	:	val_out <= 4'h5732;
         4'hf2c9 	:	val_out <= 4'h5732;
         4'hf2ca 	:	val_out <= 4'h5732;
         4'hf2cb 	:	val_out <= 4'h5732;
         4'hf2d0 	:	val_out <= 4'h574a;
         4'hf2d1 	:	val_out <= 4'h574a;
         4'hf2d2 	:	val_out <= 4'h574a;
         4'hf2d3 	:	val_out <= 4'h574a;
         4'hf2d8 	:	val_out <= 4'h5762;
         4'hf2d9 	:	val_out <= 4'h5762;
         4'hf2da 	:	val_out <= 4'h5762;
         4'hf2db 	:	val_out <= 4'h5762;
         4'hf2e0 	:	val_out <= 4'h5779;
         4'hf2e1 	:	val_out <= 4'h5779;
         4'hf2e2 	:	val_out <= 4'h5779;
         4'hf2e3 	:	val_out <= 4'h5779;
         4'hf2e8 	:	val_out <= 4'h5791;
         4'hf2e9 	:	val_out <= 4'h5791;
         4'hf2ea 	:	val_out <= 4'h5791;
         4'hf2eb 	:	val_out <= 4'h5791;
         4'hf2f0 	:	val_out <= 4'h57a9;
         4'hf2f1 	:	val_out <= 4'h57a9;
         4'hf2f2 	:	val_out <= 4'h57a9;
         4'hf2f3 	:	val_out <= 4'h57a9;
         4'hf2f8 	:	val_out <= 4'h57c1;
         4'hf2f9 	:	val_out <= 4'h57c1;
         4'hf2fa 	:	val_out <= 4'h57c1;
         4'hf2fb 	:	val_out <= 4'h57c1;
         4'hf300 	:	val_out <= 4'h57d9;
         4'hf301 	:	val_out <= 4'h57d9;
         4'hf302 	:	val_out <= 4'h57d9;
         4'hf303 	:	val_out <= 4'h57d9;
         4'hf308 	:	val_out <= 4'h57f1;
         4'hf309 	:	val_out <= 4'h57f1;
         4'hf30a 	:	val_out <= 4'h57f1;
         4'hf30b 	:	val_out <= 4'h57f1;
         4'hf310 	:	val_out <= 4'h5809;
         4'hf311 	:	val_out <= 4'h5809;
         4'hf312 	:	val_out <= 4'h5809;
         4'hf313 	:	val_out <= 4'h5809;
         4'hf318 	:	val_out <= 4'h5820;
         4'hf319 	:	val_out <= 4'h5820;
         4'hf31a 	:	val_out <= 4'h5820;
         4'hf31b 	:	val_out <= 4'h5820;
         4'hf320 	:	val_out <= 4'h5838;
         4'hf321 	:	val_out <= 4'h5838;
         4'hf322 	:	val_out <= 4'h5838;
         4'hf323 	:	val_out <= 4'h5838;
         4'hf328 	:	val_out <= 4'h5850;
         4'hf329 	:	val_out <= 4'h5850;
         4'hf32a 	:	val_out <= 4'h5850;
         4'hf32b 	:	val_out <= 4'h5850;
         4'hf330 	:	val_out <= 4'h5868;
         4'hf331 	:	val_out <= 4'h5868;
         4'hf332 	:	val_out <= 4'h5868;
         4'hf333 	:	val_out <= 4'h5868;
         4'hf338 	:	val_out <= 4'h5880;
         4'hf339 	:	val_out <= 4'h5880;
         4'hf33a 	:	val_out <= 4'h5880;
         4'hf33b 	:	val_out <= 4'h5880;
         4'hf340 	:	val_out <= 4'h5898;
         4'hf341 	:	val_out <= 4'h5898;
         4'hf342 	:	val_out <= 4'h5898;
         4'hf343 	:	val_out <= 4'h5898;
         4'hf348 	:	val_out <= 4'h58b0;
         4'hf349 	:	val_out <= 4'h58b0;
         4'hf34a 	:	val_out <= 4'h58b0;
         4'hf34b 	:	val_out <= 4'h58b0;
         4'hf350 	:	val_out <= 4'h58c8;
         4'hf351 	:	val_out <= 4'h58c8;
         4'hf352 	:	val_out <= 4'h58c8;
         4'hf353 	:	val_out <= 4'h58c8;
         4'hf358 	:	val_out <= 4'h58e0;
         4'hf359 	:	val_out <= 4'h58e0;
         4'hf35a 	:	val_out <= 4'h58e0;
         4'hf35b 	:	val_out <= 4'h58e0;
         4'hf360 	:	val_out <= 4'h58f8;
         4'hf361 	:	val_out <= 4'h58f8;
         4'hf362 	:	val_out <= 4'h58f8;
         4'hf363 	:	val_out <= 4'h58f8;
         4'hf368 	:	val_out <= 4'h5910;
         4'hf369 	:	val_out <= 4'h5910;
         4'hf36a 	:	val_out <= 4'h5910;
         4'hf36b 	:	val_out <= 4'h5910;
         4'hf370 	:	val_out <= 4'h5927;
         4'hf371 	:	val_out <= 4'h5927;
         4'hf372 	:	val_out <= 4'h5927;
         4'hf373 	:	val_out <= 4'h5927;
         4'hf378 	:	val_out <= 4'h593f;
         4'hf379 	:	val_out <= 4'h593f;
         4'hf37a 	:	val_out <= 4'h593f;
         4'hf37b 	:	val_out <= 4'h593f;
         4'hf380 	:	val_out <= 4'h5957;
         4'hf381 	:	val_out <= 4'h5957;
         4'hf382 	:	val_out <= 4'h5957;
         4'hf383 	:	val_out <= 4'h5957;
         4'hf388 	:	val_out <= 4'h596f;
         4'hf389 	:	val_out <= 4'h596f;
         4'hf38a 	:	val_out <= 4'h596f;
         4'hf38b 	:	val_out <= 4'h596f;
         4'hf390 	:	val_out <= 4'h5987;
         4'hf391 	:	val_out <= 4'h5987;
         4'hf392 	:	val_out <= 4'h5987;
         4'hf393 	:	val_out <= 4'h5987;
         4'hf398 	:	val_out <= 4'h599f;
         4'hf399 	:	val_out <= 4'h599f;
         4'hf39a 	:	val_out <= 4'h599f;
         4'hf39b 	:	val_out <= 4'h599f;
         4'hf3a0 	:	val_out <= 4'h59b7;
         4'hf3a1 	:	val_out <= 4'h59b7;
         4'hf3a2 	:	val_out <= 4'h59b7;
         4'hf3a3 	:	val_out <= 4'h59b7;
         4'hf3a8 	:	val_out <= 4'h59cf;
         4'hf3a9 	:	val_out <= 4'h59cf;
         4'hf3aa 	:	val_out <= 4'h59cf;
         4'hf3ab 	:	val_out <= 4'h59cf;
         4'hf3b0 	:	val_out <= 4'h59e7;
         4'hf3b1 	:	val_out <= 4'h59e7;
         4'hf3b2 	:	val_out <= 4'h59e7;
         4'hf3b3 	:	val_out <= 4'h59e7;
         4'hf3b8 	:	val_out <= 4'h59ff;
         4'hf3b9 	:	val_out <= 4'h59ff;
         4'hf3ba 	:	val_out <= 4'h59ff;
         4'hf3bb 	:	val_out <= 4'h59ff;
         4'hf3c0 	:	val_out <= 4'h5a17;
         4'hf3c1 	:	val_out <= 4'h5a17;
         4'hf3c2 	:	val_out <= 4'h5a17;
         4'hf3c3 	:	val_out <= 4'h5a17;
         4'hf3c8 	:	val_out <= 4'h5a2f;
         4'hf3c9 	:	val_out <= 4'h5a2f;
         4'hf3ca 	:	val_out <= 4'h5a2f;
         4'hf3cb 	:	val_out <= 4'h5a2f;
         4'hf3d0 	:	val_out <= 4'h5a47;
         4'hf3d1 	:	val_out <= 4'h5a47;
         4'hf3d2 	:	val_out <= 4'h5a47;
         4'hf3d3 	:	val_out <= 4'h5a47;
         4'hf3d8 	:	val_out <= 4'h5a5f;
         4'hf3d9 	:	val_out <= 4'h5a5f;
         4'hf3da 	:	val_out <= 4'h5a5f;
         4'hf3db 	:	val_out <= 4'h5a5f;
         4'hf3e0 	:	val_out <= 4'h5a77;
         4'hf3e1 	:	val_out <= 4'h5a77;
         4'hf3e2 	:	val_out <= 4'h5a77;
         4'hf3e3 	:	val_out <= 4'h5a77;
         4'hf3e8 	:	val_out <= 4'h5a8f;
         4'hf3e9 	:	val_out <= 4'h5a8f;
         4'hf3ea 	:	val_out <= 4'h5a8f;
         4'hf3eb 	:	val_out <= 4'h5a8f;
         4'hf3f0 	:	val_out <= 4'h5aa7;
         4'hf3f1 	:	val_out <= 4'h5aa7;
         4'hf3f2 	:	val_out <= 4'h5aa7;
         4'hf3f3 	:	val_out <= 4'h5aa7;
         4'hf3f8 	:	val_out <= 4'h5abf;
         4'hf3f9 	:	val_out <= 4'h5abf;
         4'hf3fa 	:	val_out <= 4'h5abf;
         4'hf3fb 	:	val_out <= 4'h5abf;
         4'hf400 	:	val_out <= 4'h5ad7;
         4'hf401 	:	val_out <= 4'h5ad7;
         4'hf402 	:	val_out <= 4'h5ad7;
         4'hf403 	:	val_out <= 4'h5ad7;
         4'hf408 	:	val_out <= 4'h5af0;
         4'hf409 	:	val_out <= 4'h5af0;
         4'hf40a 	:	val_out <= 4'h5af0;
         4'hf40b 	:	val_out <= 4'h5af0;
         4'hf410 	:	val_out <= 4'h5b08;
         4'hf411 	:	val_out <= 4'h5b08;
         4'hf412 	:	val_out <= 4'h5b08;
         4'hf413 	:	val_out <= 4'h5b08;
         4'hf418 	:	val_out <= 4'h5b20;
         4'hf419 	:	val_out <= 4'h5b20;
         4'hf41a 	:	val_out <= 4'h5b20;
         4'hf41b 	:	val_out <= 4'h5b20;
         4'hf420 	:	val_out <= 4'h5b38;
         4'hf421 	:	val_out <= 4'h5b38;
         4'hf422 	:	val_out <= 4'h5b38;
         4'hf423 	:	val_out <= 4'h5b38;
         4'hf428 	:	val_out <= 4'h5b50;
         4'hf429 	:	val_out <= 4'h5b50;
         4'hf42a 	:	val_out <= 4'h5b50;
         4'hf42b 	:	val_out <= 4'h5b50;
         4'hf430 	:	val_out <= 4'h5b68;
         4'hf431 	:	val_out <= 4'h5b68;
         4'hf432 	:	val_out <= 4'h5b68;
         4'hf433 	:	val_out <= 4'h5b68;
         4'hf438 	:	val_out <= 4'h5b80;
         4'hf439 	:	val_out <= 4'h5b80;
         4'hf43a 	:	val_out <= 4'h5b80;
         4'hf43b 	:	val_out <= 4'h5b80;
         4'hf440 	:	val_out <= 4'h5b98;
         4'hf441 	:	val_out <= 4'h5b98;
         4'hf442 	:	val_out <= 4'h5b98;
         4'hf443 	:	val_out <= 4'h5b98;
         4'hf448 	:	val_out <= 4'h5bb0;
         4'hf449 	:	val_out <= 4'h5bb0;
         4'hf44a 	:	val_out <= 4'h5bb0;
         4'hf44b 	:	val_out <= 4'h5bb0;
         4'hf450 	:	val_out <= 4'h5bc8;
         4'hf451 	:	val_out <= 4'h5bc8;
         4'hf452 	:	val_out <= 4'h5bc8;
         4'hf453 	:	val_out <= 4'h5bc8;
         4'hf458 	:	val_out <= 4'h5be0;
         4'hf459 	:	val_out <= 4'h5be0;
         4'hf45a 	:	val_out <= 4'h5be0;
         4'hf45b 	:	val_out <= 4'h5be0;
         4'hf460 	:	val_out <= 4'h5bf8;
         4'hf461 	:	val_out <= 4'h5bf8;
         4'hf462 	:	val_out <= 4'h5bf8;
         4'hf463 	:	val_out <= 4'h5bf8;
         4'hf468 	:	val_out <= 4'h5c11;
         4'hf469 	:	val_out <= 4'h5c11;
         4'hf46a 	:	val_out <= 4'h5c11;
         4'hf46b 	:	val_out <= 4'h5c11;
         4'hf470 	:	val_out <= 4'h5c29;
         4'hf471 	:	val_out <= 4'h5c29;
         4'hf472 	:	val_out <= 4'h5c29;
         4'hf473 	:	val_out <= 4'h5c29;
         4'hf478 	:	val_out <= 4'h5c41;
         4'hf479 	:	val_out <= 4'h5c41;
         4'hf47a 	:	val_out <= 4'h5c41;
         4'hf47b 	:	val_out <= 4'h5c41;
         4'hf480 	:	val_out <= 4'h5c59;
         4'hf481 	:	val_out <= 4'h5c59;
         4'hf482 	:	val_out <= 4'h5c59;
         4'hf483 	:	val_out <= 4'h5c59;
         4'hf488 	:	val_out <= 4'h5c71;
         4'hf489 	:	val_out <= 4'h5c71;
         4'hf48a 	:	val_out <= 4'h5c71;
         4'hf48b 	:	val_out <= 4'h5c71;
         4'hf490 	:	val_out <= 4'h5c89;
         4'hf491 	:	val_out <= 4'h5c89;
         4'hf492 	:	val_out <= 4'h5c89;
         4'hf493 	:	val_out <= 4'h5c89;
         4'hf498 	:	val_out <= 4'h5ca1;
         4'hf499 	:	val_out <= 4'h5ca1;
         4'hf49a 	:	val_out <= 4'h5ca1;
         4'hf49b 	:	val_out <= 4'h5ca1;
         4'hf4a0 	:	val_out <= 4'h5cba;
         4'hf4a1 	:	val_out <= 4'h5cba;
         4'hf4a2 	:	val_out <= 4'h5cba;
         4'hf4a3 	:	val_out <= 4'h5cba;
         4'hf4a8 	:	val_out <= 4'h5cd2;
         4'hf4a9 	:	val_out <= 4'h5cd2;
         4'hf4aa 	:	val_out <= 4'h5cd2;
         4'hf4ab 	:	val_out <= 4'h5cd2;
         4'hf4b0 	:	val_out <= 4'h5cea;
         4'hf4b1 	:	val_out <= 4'h5cea;
         4'hf4b2 	:	val_out <= 4'h5cea;
         4'hf4b3 	:	val_out <= 4'h5cea;
         4'hf4b8 	:	val_out <= 4'h5d02;
         4'hf4b9 	:	val_out <= 4'h5d02;
         4'hf4ba 	:	val_out <= 4'h5d02;
         4'hf4bb 	:	val_out <= 4'h5d02;
         4'hf4c0 	:	val_out <= 4'h5d1a;
         4'hf4c1 	:	val_out <= 4'h5d1a;
         4'hf4c2 	:	val_out <= 4'h5d1a;
         4'hf4c3 	:	val_out <= 4'h5d1a;
         4'hf4c8 	:	val_out <= 4'h5d32;
         4'hf4c9 	:	val_out <= 4'h5d32;
         4'hf4ca 	:	val_out <= 4'h5d32;
         4'hf4cb 	:	val_out <= 4'h5d32;
         4'hf4d0 	:	val_out <= 4'h5d4b;
         4'hf4d1 	:	val_out <= 4'h5d4b;
         4'hf4d2 	:	val_out <= 4'h5d4b;
         4'hf4d3 	:	val_out <= 4'h5d4b;
         4'hf4d8 	:	val_out <= 4'h5d63;
         4'hf4d9 	:	val_out <= 4'h5d63;
         4'hf4da 	:	val_out <= 4'h5d63;
         4'hf4db 	:	val_out <= 4'h5d63;
         4'hf4e0 	:	val_out <= 4'h5d7b;
         4'hf4e1 	:	val_out <= 4'h5d7b;
         4'hf4e2 	:	val_out <= 4'h5d7b;
         4'hf4e3 	:	val_out <= 4'h5d7b;
         4'hf4e8 	:	val_out <= 4'h5d93;
         4'hf4e9 	:	val_out <= 4'h5d93;
         4'hf4ea 	:	val_out <= 4'h5d93;
         4'hf4eb 	:	val_out <= 4'h5d93;
         4'hf4f0 	:	val_out <= 4'h5dab;
         4'hf4f1 	:	val_out <= 4'h5dab;
         4'hf4f2 	:	val_out <= 4'h5dab;
         4'hf4f3 	:	val_out <= 4'h5dab;
         4'hf4f8 	:	val_out <= 4'h5dc4;
         4'hf4f9 	:	val_out <= 4'h5dc4;
         4'hf4fa 	:	val_out <= 4'h5dc4;
         4'hf4fb 	:	val_out <= 4'h5dc4;
         4'hf500 	:	val_out <= 4'h5ddc;
         4'hf501 	:	val_out <= 4'h5ddc;
         4'hf502 	:	val_out <= 4'h5ddc;
         4'hf503 	:	val_out <= 4'h5ddc;
         4'hf508 	:	val_out <= 4'h5df4;
         4'hf509 	:	val_out <= 4'h5df4;
         4'hf50a 	:	val_out <= 4'h5df4;
         4'hf50b 	:	val_out <= 4'h5df4;
         4'hf510 	:	val_out <= 4'h5e0c;
         4'hf511 	:	val_out <= 4'h5e0c;
         4'hf512 	:	val_out <= 4'h5e0c;
         4'hf513 	:	val_out <= 4'h5e0c;
         4'hf518 	:	val_out <= 4'h5e25;
         4'hf519 	:	val_out <= 4'h5e25;
         4'hf51a 	:	val_out <= 4'h5e25;
         4'hf51b 	:	val_out <= 4'h5e25;
         4'hf520 	:	val_out <= 4'h5e3d;
         4'hf521 	:	val_out <= 4'h5e3d;
         4'hf522 	:	val_out <= 4'h5e3d;
         4'hf523 	:	val_out <= 4'h5e3d;
         4'hf528 	:	val_out <= 4'h5e55;
         4'hf529 	:	val_out <= 4'h5e55;
         4'hf52a 	:	val_out <= 4'h5e55;
         4'hf52b 	:	val_out <= 4'h5e55;
         4'hf530 	:	val_out <= 4'h5e6d;
         4'hf531 	:	val_out <= 4'h5e6d;
         4'hf532 	:	val_out <= 4'h5e6d;
         4'hf533 	:	val_out <= 4'h5e6d;
         4'hf538 	:	val_out <= 4'h5e86;
         4'hf539 	:	val_out <= 4'h5e86;
         4'hf53a 	:	val_out <= 4'h5e86;
         4'hf53b 	:	val_out <= 4'h5e86;
         4'hf540 	:	val_out <= 4'h5e9e;
         4'hf541 	:	val_out <= 4'h5e9e;
         4'hf542 	:	val_out <= 4'h5e9e;
         4'hf543 	:	val_out <= 4'h5e9e;
         4'hf548 	:	val_out <= 4'h5eb6;
         4'hf549 	:	val_out <= 4'h5eb6;
         4'hf54a 	:	val_out <= 4'h5eb6;
         4'hf54b 	:	val_out <= 4'h5eb6;
         4'hf550 	:	val_out <= 4'h5ece;
         4'hf551 	:	val_out <= 4'h5ece;
         4'hf552 	:	val_out <= 4'h5ece;
         4'hf553 	:	val_out <= 4'h5ece;
         4'hf558 	:	val_out <= 4'h5ee7;
         4'hf559 	:	val_out <= 4'h5ee7;
         4'hf55a 	:	val_out <= 4'h5ee7;
         4'hf55b 	:	val_out <= 4'h5ee7;
         4'hf560 	:	val_out <= 4'h5eff;
         4'hf561 	:	val_out <= 4'h5eff;
         4'hf562 	:	val_out <= 4'h5eff;
         4'hf563 	:	val_out <= 4'h5eff;
         4'hf568 	:	val_out <= 4'h5f17;
         4'hf569 	:	val_out <= 4'h5f17;
         4'hf56a 	:	val_out <= 4'h5f17;
         4'hf56b 	:	val_out <= 4'h5f17;
         4'hf570 	:	val_out <= 4'h5f2f;
         4'hf571 	:	val_out <= 4'h5f2f;
         4'hf572 	:	val_out <= 4'h5f2f;
         4'hf573 	:	val_out <= 4'h5f2f;
         4'hf578 	:	val_out <= 4'h5f48;
         4'hf579 	:	val_out <= 4'h5f48;
         4'hf57a 	:	val_out <= 4'h5f48;
         4'hf57b 	:	val_out <= 4'h5f48;
         4'hf580 	:	val_out <= 4'h5f60;
         4'hf581 	:	val_out <= 4'h5f60;
         4'hf582 	:	val_out <= 4'h5f60;
         4'hf583 	:	val_out <= 4'h5f60;
         4'hf588 	:	val_out <= 4'h5f78;
         4'hf589 	:	val_out <= 4'h5f78;
         4'hf58a 	:	val_out <= 4'h5f78;
         4'hf58b 	:	val_out <= 4'h5f78;
         4'hf590 	:	val_out <= 4'h5f91;
         4'hf591 	:	val_out <= 4'h5f91;
         4'hf592 	:	val_out <= 4'h5f91;
         4'hf593 	:	val_out <= 4'h5f91;
         4'hf598 	:	val_out <= 4'h5fa9;
         4'hf599 	:	val_out <= 4'h5fa9;
         4'hf59a 	:	val_out <= 4'h5fa9;
         4'hf59b 	:	val_out <= 4'h5fa9;
         4'hf5a0 	:	val_out <= 4'h5fc1;
         4'hf5a1 	:	val_out <= 4'h5fc1;
         4'hf5a2 	:	val_out <= 4'h5fc1;
         4'hf5a3 	:	val_out <= 4'h5fc1;
         4'hf5a8 	:	val_out <= 4'h5fda;
         4'hf5a9 	:	val_out <= 4'h5fda;
         4'hf5aa 	:	val_out <= 4'h5fda;
         4'hf5ab 	:	val_out <= 4'h5fda;
         4'hf5b0 	:	val_out <= 4'h5ff2;
         4'hf5b1 	:	val_out <= 4'h5ff2;
         4'hf5b2 	:	val_out <= 4'h5ff2;
         4'hf5b3 	:	val_out <= 4'h5ff2;
         4'hf5b8 	:	val_out <= 4'h600a;
         4'hf5b9 	:	val_out <= 4'h600a;
         4'hf5ba 	:	val_out <= 4'h600a;
         4'hf5bb 	:	val_out <= 4'h600a;
         4'hf5c0 	:	val_out <= 4'h6023;
         4'hf5c1 	:	val_out <= 4'h6023;
         4'hf5c2 	:	val_out <= 4'h6023;
         4'hf5c3 	:	val_out <= 4'h6023;
         4'hf5c8 	:	val_out <= 4'h603b;
         4'hf5c9 	:	val_out <= 4'h603b;
         4'hf5ca 	:	val_out <= 4'h603b;
         4'hf5cb 	:	val_out <= 4'h603b;
         4'hf5d0 	:	val_out <= 4'h6053;
         4'hf5d1 	:	val_out <= 4'h6053;
         4'hf5d2 	:	val_out <= 4'h6053;
         4'hf5d3 	:	val_out <= 4'h6053;
         4'hf5d8 	:	val_out <= 4'h606c;
         4'hf5d9 	:	val_out <= 4'h606c;
         4'hf5da 	:	val_out <= 4'h606c;
         4'hf5db 	:	val_out <= 4'h606c;
         4'hf5e0 	:	val_out <= 4'h6084;
         4'hf5e1 	:	val_out <= 4'h6084;
         4'hf5e2 	:	val_out <= 4'h6084;
         4'hf5e3 	:	val_out <= 4'h6084;
         4'hf5e8 	:	val_out <= 4'h609c;
         4'hf5e9 	:	val_out <= 4'h609c;
         4'hf5ea 	:	val_out <= 4'h609c;
         4'hf5eb 	:	val_out <= 4'h609c;
         4'hf5f0 	:	val_out <= 4'h60b5;
         4'hf5f1 	:	val_out <= 4'h60b5;
         4'hf5f2 	:	val_out <= 4'h60b5;
         4'hf5f3 	:	val_out <= 4'h60b5;
         4'hf5f8 	:	val_out <= 4'h60cd;
         4'hf5f9 	:	val_out <= 4'h60cd;
         4'hf5fa 	:	val_out <= 4'h60cd;
         4'hf5fb 	:	val_out <= 4'h60cd;
         4'hf600 	:	val_out <= 4'h60e6;
         4'hf601 	:	val_out <= 4'h60e6;
         4'hf602 	:	val_out <= 4'h60e6;
         4'hf603 	:	val_out <= 4'h60e6;
         4'hf608 	:	val_out <= 4'h60fe;
         4'hf609 	:	val_out <= 4'h60fe;
         4'hf60a 	:	val_out <= 4'h60fe;
         4'hf60b 	:	val_out <= 4'h60fe;
         4'hf610 	:	val_out <= 4'h6116;
         4'hf611 	:	val_out <= 4'h6116;
         4'hf612 	:	val_out <= 4'h6116;
         4'hf613 	:	val_out <= 4'h6116;
         4'hf618 	:	val_out <= 4'h612f;
         4'hf619 	:	val_out <= 4'h612f;
         4'hf61a 	:	val_out <= 4'h612f;
         4'hf61b 	:	val_out <= 4'h612f;
         4'hf620 	:	val_out <= 4'h6147;
         4'hf621 	:	val_out <= 4'h6147;
         4'hf622 	:	val_out <= 4'h6147;
         4'hf623 	:	val_out <= 4'h6147;
         4'hf628 	:	val_out <= 4'h615f;
         4'hf629 	:	val_out <= 4'h615f;
         4'hf62a 	:	val_out <= 4'h615f;
         4'hf62b 	:	val_out <= 4'h615f;
         4'hf630 	:	val_out <= 4'h6178;
         4'hf631 	:	val_out <= 4'h6178;
         4'hf632 	:	val_out <= 4'h6178;
         4'hf633 	:	val_out <= 4'h6178;
         4'hf638 	:	val_out <= 4'h6190;
         4'hf639 	:	val_out <= 4'h6190;
         4'hf63a 	:	val_out <= 4'h6190;
         4'hf63b 	:	val_out <= 4'h6190;
         4'hf640 	:	val_out <= 4'h61a9;
         4'hf641 	:	val_out <= 4'h61a9;
         4'hf642 	:	val_out <= 4'h61a9;
         4'hf643 	:	val_out <= 4'h61a9;
         4'hf648 	:	val_out <= 4'h61c1;
         4'hf649 	:	val_out <= 4'h61c1;
         4'hf64a 	:	val_out <= 4'h61c1;
         4'hf64b 	:	val_out <= 4'h61c1;
         4'hf650 	:	val_out <= 4'h61da;
         4'hf651 	:	val_out <= 4'h61da;
         4'hf652 	:	val_out <= 4'h61da;
         4'hf653 	:	val_out <= 4'h61da;
         4'hf658 	:	val_out <= 4'h61f2;
         4'hf659 	:	val_out <= 4'h61f2;
         4'hf65a 	:	val_out <= 4'h61f2;
         4'hf65b 	:	val_out <= 4'h61f2;
         4'hf660 	:	val_out <= 4'h620a;
         4'hf661 	:	val_out <= 4'h620a;
         4'hf662 	:	val_out <= 4'h620a;
         4'hf663 	:	val_out <= 4'h620a;
         4'hf668 	:	val_out <= 4'h6223;
         4'hf669 	:	val_out <= 4'h6223;
         4'hf66a 	:	val_out <= 4'h6223;
         4'hf66b 	:	val_out <= 4'h6223;
         4'hf670 	:	val_out <= 4'h623b;
         4'hf671 	:	val_out <= 4'h623b;
         4'hf672 	:	val_out <= 4'h623b;
         4'hf673 	:	val_out <= 4'h623b;
         4'hf678 	:	val_out <= 4'h6254;
         4'hf679 	:	val_out <= 4'h6254;
         4'hf67a 	:	val_out <= 4'h6254;
         4'hf67b 	:	val_out <= 4'h6254;
         4'hf680 	:	val_out <= 4'h626c;
         4'hf681 	:	val_out <= 4'h626c;
         4'hf682 	:	val_out <= 4'h626c;
         4'hf683 	:	val_out <= 4'h626c;
         4'hf688 	:	val_out <= 4'h6285;
         4'hf689 	:	val_out <= 4'h6285;
         4'hf68a 	:	val_out <= 4'h6285;
         4'hf68b 	:	val_out <= 4'h6285;
         4'hf690 	:	val_out <= 4'h629d;
         4'hf691 	:	val_out <= 4'h629d;
         4'hf692 	:	val_out <= 4'h629d;
         4'hf693 	:	val_out <= 4'h629d;
         4'hf698 	:	val_out <= 4'h62b6;
         4'hf699 	:	val_out <= 4'h62b6;
         4'hf69a 	:	val_out <= 4'h62b6;
         4'hf69b 	:	val_out <= 4'h62b6;
         4'hf6a0 	:	val_out <= 4'h62ce;
         4'hf6a1 	:	val_out <= 4'h62ce;
         4'hf6a2 	:	val_out <= 4'h62ce;
         4'hf6a3 	:	val_out <= 4'h62ce;
         4'hf6a8 	:	val_out <= 4'h62e7;
         4'hf6a9 	:	val_out <= 4'h62e7;
         4'hf6aa 	:	val_out <= 4'h62e7;
         4'hf6ab 	:	val_out <= 4'h62e7;
         4'hf6b0 	:	val_out <= 4'h62ff;
         4'hf6b1 	:	val_out <= 4'h62ff;
         4'hf6b2 	:	val_out <= 4'h62ff;
         4'hf6b3 	:	val_out <= 4'h62ff;
         4'hf6b8 	:	val_out <= 4'h6317;
         4'hf6b9 	:	val_out <= 4'h6317;
         4'hf6ba 	:	val_out <= 4'h6317;
         4'hf6bb 	:	val_out <= 4'h6317;
         4'hf6c0 	:	val_out <= 4'h6330;
         4'hf6c1 	:	val_out <= 4'h6330;
         4'hf6c2 	:	val_out <= 4'h6330;
         4'hf6c3 	:	val_out <= 4'h6330;
         4'hf6c8 	:	val_out <= 4'h6348;
         4'hf6c9 	:	val_out <= 4'h6348;
         4'hf6ca 	:	val_out <= 4'h6348;
         4'hf6cb 	:	val_out <= 4'h6348;
         4'hf6d0 	:	val_out <= 4'h6361;
         4'hf6d1 	:	val_out <= 4'h6361;
         4'hf6d2 	:	val_out <= 4'h6361;
         4'hf6d3 	:	val_out <= 4'h6361;
         4'hf6d8 	:	val_out <= 4'h6379;
         4'hf6d9 	:	val_out <= 4'h6379;
         4'hf6da 	:	val_out <= 4'h6379;
         4'hf6db 	:	val_out <= 4'h6379;
         4'hf6e0 	:	val_out <= 4'h6392;
         4'hf6e1 	:	val_out <= 4'h6392;
         4'hf6e2 	:	val_out <= 4'h6392;
         4'hf6e3 	:	val_out <= 4'h6392;
         4'hf6e8 	:	val_out <= 4'h63aa;
         4'hf6e9 	:	val_out <= 4'h63aa;
         4'hf6ea 	:	val_out <= 4'h63aa;
         4'hf6eb 	:	val_out <= 4'h63aa;
         4'hf6f0 	:	val_out <= 4'h63c3;
         4'hf6f1 	:	val_out <= 4'h63c3;
         4'hf6f2 	:	val_out <= 4'h63c3;
         4'hf6f3 	:	val_out <= 4'h63c3;
         4'hf6f8 	:	val_out <= 4'h63db;
         4'hf6f9 	:	val_out <= 4'h63db;
         4'hf6fa 	:	val_out <= 4'h63db;
         4'hf6fb 	:	val_out <= 4'h63db;
         4'hf700 	:	val_out <= 4'h63f4;
         4'hf701 	:	val_out <= 4'h63f4;
         4'hf702 	:	val_out <= 4'h63f4;
         4'hf703 	:	val_out <= 4'h63f4;
         4'hf708 	:	val_out <= 4'h640d;
         4'hf709 	:	val_out <= 4'h640d;
         4'hf70a 	:	val_out <= 4'h640d;
         4'hf70b 	:	val_out <= 4'h640d;
         4'hf710 	:	val_out <= 4'h6425;
         4'hf711 	:	val_out <= 4'h6425;
         4'hf712 	:	val_out <= 4'h6425;
         4'hf713 	:	val_out <= 4'h6425;
         4'hf718 	:	val_out <= 4'h643e;
         4'hf719 	:	val_out <= 4'h643e;
         4'hf71a 	:	val_out <= 4'h643e;
         4'hf71b 	:	val_out <= 4'h643e;
         4'hf720 	:	val_out <= 4'h6456;
         4'hf721 	:	val_out <= 4'h6456;
         4'hf722 	:	val_out <= 4'h6456;
         4'hf723 	:	val_out <= 4'h6456;
         4'hf728 	:	val_out <= 4'h646f;
         4'hf729 	:	val_out <= 4'h646f;
         4'hf72a 	:	val_out <= 4'h646f;
         4'hf72b 	:	val_out <= 4'h646f;
         4'hf730 	:	val_out <= 4'h6487;
         4'hf731 	:	val_out <= 4'h6487;
         4'hf732 	:	val_out <= 4'h6487;
         4'hf733 	:	val_out <= 4'h6487;
         4'hf738 	:	val_out <= 4'h64a0;
         4'hf739 	:	val_out <= 4'h64a0;
         4'hf73a 	:	val_out <= 4'h64a0;
         4'hf73b 	:	val_out <= 4'h64a0;
         4'hf740 	:	val_out <= 4'h64b8;
         4'hf741 	:	val_out <= 4'h64b8;
         4'hf742 	:	val_out <= 4'h64b8;
         4'hf743 	:	val_out <= 4'h64b8;
         4'hf748 	:	val_out <= 4'h64d1;
         4'hf749 	:	val_out <= 4'h64d1;
         4'hf74a 	:	val_out <= 4'h64d1;
         4'hf74b 	:	val_out <= 4'h64d1;
         4'hf750 	:	val_out <= 4'h64e9;
         4'hf751 	:	val_out <= 4'h64e9;
         4'hf752 	:	val_out <= 4'h64e9;
         4'hf753 	:	val_out <= 4'h64e9;
         4'hf758 	:	val_out <= 4'h6502;
         4'hf759 	:	val_out <= 4'h6502;
         4'hf75a 	:	val_out <= 4'h6502;
         4'hf75b 	:	val_out <= 4'h6502;
         4'hf760 	:	val_out <= 4'h651b;
         4'hf761 	:	val_out <= 4'h651b;
         4'hf762 	:	val_out <= 4'h651b;
         4'hf763 	:	val_out <= 4'h651b;
         4'hf768 	:	val_out <= 4'h6533;
         4'hf769 	:	val_out <= 4'h6533;
         4'hf76a 	:	val_out <= 4'h6533;
         4'hf76b 	:	val_out <= 4'h6533;
         4'hf770 	:	val_out <= 4'h654c;
         4'hf771 	:	val_out <= 4'h654c;
         4'hf772 	:	val_out <= 4'h654c;
         4'hf773 	:	val_out <= 4'h654c;
         4'hf778 	:	val_out <= 4'h6564;
         4'hf779 	:	val_out <= 4'h6564;
         4'hf77a 	:	val_out <= 4'h6564;
         4'hf77b 	:	val_out <= 4'h6564;
         4'hf780 	:	val_out <= 4'h657d;
         4'hf781 	:	val_out <= 4'h657d;
         4'hf782 	:	val_out <= 4'h657d;
         4'hf783 	:	val_out <= 4'h657d;
         4'hf788 	:	val_out <= 4'h6595;
         4'hf789 	:	val_out <= 4'h6595;
         4'hf78a 	:	val_out <= 4'h6595;
         4'hf78b 	:	val_out <= 4'h6595;
         4'hf790 	:	val_out <= 4'h65ae;
         4'hf791 	:	val_out <= 4'h65ae;
         4'hf792 	:	val_out <= 4'h65ae;
         4'hf793 	:	val_out <= 4'h65ae;
         4'hf798 	:	val_out <= 4'h65c7;
         4'hf799 	:	val_out <= 4'h65c7;
         4'hf79a 	:	val_out <= 4'h65c7;
         4'hf79b 	:	val_out <= 4'h65c7;
         4'hf7a0 	:	val_out <= 4'h65df;
         4'hf7a1 	:	val_out <= 4'h65df;
         4'hf7a2 	:	val_out <= 4'h65df;
         4'hf7a3 	:	val_out <= 4'h65df;
         4'hf7a8 	:	val_out <= 4'h65f8;
         4'hf7a9 	:	val_out <= 4'h65f8;
         4'hf7aa 	:	val_out <= 4'h65f8;
         4'hf7ab 	:	val_out <= 4'h65f8;
         4'hf7b0 	:	val_out <= 4'h6610;
         4'hf7b1 	:	val_out <= 4'h6610;
         4'hf7b2 	:	val_out <= 4'h6610;
         4'hf7b3 	:	val_out <= 4'h6610;
         4'hf7b8 	:	val_out <= 4'h6629;
         4'hf7b9 	:	val_out <= 4'h6629;
         4'hf7ba 	:	val_out <= 4'h6629;
         4'hf7bb 	:	val_out <= 4'h6629;
         4'hf7c0 	:	val_out <= 4'h6642;
         4'hf7c1 	:	val_out <= 4'h6642;
         4'hf7c2 	:	val_out <= 4'h6642;
         4'hf7c3 	:	val_out <= 4'h6642;
         4'hf7c8 	:	val_out <= 4'h665a;
         4'hf7c9 	:	val_out <= 4'h665a;
         4'hf7ca 	:	val_out <= 4'h665a;
         4'hf7cb 	:	val_out <= 4'h665a;
         4'hf7d0 	:	val_out <= 4'h6673;
         4'hf7d1 	:	val_out <= 4'h6673;
         4'hf7d2 	:	val_out <= 4'h6673;
         4'hf7d3 	:	val_out <= 4'h6673;
         4'hf7d8 	:	val_out <= 4'h668c;
         4'hf7d9 	:	val_out <= 4'h668c;
         4'hf7da 	:	val_out <= 4'h668c;
         4'hf7db 	:	val_out <= 4'h668c;
         4'hf7e0 	:	val_out <= 4'h66a4;
         4'hf7e1 	:	val_out <= 4'h66a4;
         4'hf7e2 	:	val_out <= 4'h66a4;
         4'hf7e3 	:	val_out <= 4'h66a4;
         4'hf7e8 	:	val_out <= 4'h66bd;
         4'hf7e9 	:	val_out <= 4'h66bd;
         4'hf7ea 	:	val_out <= 4'h66bd;
         4'hf7eb 	:	val_out <= 4'h66bd;
         4'hf7f0 	:	val_out <= 4'h66d5;
         4'hf7f1 	:	val_out <= 4'h66d5;
         4'hf7f2 	:	val_out <= 4'h66d5;
         4'hf7f3 	:	val_out <= 4'h66d5;
         4'hf7f8 	:	val_out <= 4'h66ee;
         4'hf7f9 	:	val_out <= 4'h66ee;
         4'hf7fa 	:	val_out <= 4'h66ee;
         4'hf7fb 	:	val_out <= 4'h66ee;
         4'hf800 	:	val_out <= 4'h6707;
         4'hf801 	:	val_out <= 4'h6707;
         4'hf802 	:	val_out <= 4'h6707;
         4'hf803 	:	val_out <= 4'h6707;
         4'hf808 	:	val_out <= 4'h671f;
         4'hf809 	:	val_out <= 4'h671f;
         4'hf80a 	:	val_out <= 4'h671f;
         4'hf80b 	:	val_out <= 4'h671f;
         4'hf810 	:	val_out <= 4'h6738;
         4'hf811 	:	val_out <= 4'h6738;
         4'hf812 	:	val_out <= 4'h6738;
         4'hf813 	:	val_out <= 4'h6738;
         4'hf818 	:	val_out <= 4'h6751;
         4'hf819 	:	val_out <= 4'h6751;
         4'hf81a 	:	val_out <= 4'h6751;
         4'hf81b 	:	val_out <= 4'h6751;
         4'hf820 	:	val_out <= 4'h6769;
         4'hf821 	:	val_out <= 4'h6769;
         4'hf822 	:	val_out <= 4'h6769;
         4'hf823 	:	val_out <= 4'h6769;
         4'hf828 	:	val_out <= 4'h6782;
         4'hf829 	:	val_out <= 4'h6782;
         4'hf82a 	:	val_out <= 4'h6782;
         4'hf82b 	:	val_out <= 4'h6782;
         4'hf830 	:	val_out <= 4'h679b;
         4'hf831 	:	val_out <= 4'h679b;
         4'hf832 	:	val_out <= 4'h679b;
         4'hf833 	:	val_out <= 4'h679b;
         4'hf838 	:	val_out <= 4'h67b3;
         4'hf839 	:	val_out <= 4'h67b3;
         4'hf83a 	:	val_out <= 4'h67b3;
         4'hf83b 	:	val_out <= 4'h67b3;
         4'hf840 	:	val_out <= 4'h67cc;
         4'hf841 	:	val_out <= 4'h67cc;
         4'hf842 	:	val_out <= 4'h67cc;
         4'hf843 	:	val_out <= 4'h67cc;
         4'hf848 	:	val_out <= 4'h67e5;
         4'hf849 	:	val_out <= 4'h67e5;
         4'hf84a 	:	val_out <= 4'h67e5;
         4'hf84b 	:	val_out <= 4'h67e5;
         4'hf850 	:	val_out <= 4'h67fd;
         4'hf851 	:	val_out <= 4'h67fd;
         4'hf852 	:	val_out <= 4'h67fd;
         4'hf853 	:	val_out <= 4'h67fd;
         4'hf858 	:	val_out <= 4'h6816;
         4'hf859 	:	val_out <= 4'h6816;
         4'hf85a 	:	val_out <= 4'h6816;
         4'hf85b 	:	val_out <= 4'h6816;
         4'hf860 	:	val_out <= 4'h682f;
         4'hf861 	:	val_out <= 4'h682f;
         4'hf862 	:	val_out <= 4'h682f;
         4'hf863 	:	val_out <= 4'h682f;
         4'hf868 	:	val_out <= 4'h6848;
         4'hf869 	:	val_out <= 4'h6848;
         4'hf86a 	:	val_out <= 4'h6848;
         4'hf86b 	:	val_out <= 4'h6848;
         4'hf870 	:	val_out <= 4'h6860;
         4'hf871 	:	val_out <= 4'h6860;
         4'hf872 	:	val_out <= 4'h6860;
         4'hf873 	:	val_out <= 4'h6860;
         4'hf878 	:	val_out <= 4'h6879;
         4'hf879 	:	val_out <= 4'h6879;
         4'hf87a 	:	val_out <= 4'h6879;
         4'hf87b 	:	val_out <= 4'h6879;
         4'hf880 	:	val_out <= 4'h6892;
         4'hf881 	:	val_out <= 4'h6892;
         4'hf882 	:	val_out <= 4'h6892;
         4'hf883 	:	val_out <= 4'h6892;
         4'hf888 	:	val_out <= 4'h68aa;
         4'hf889 	:	val_out <= 4'h68aa;
         4'hf88a 	:	val_out <= 4'h68aa;
         4'hf88b 	:	val_out <= 4'h68aa;
         4'hf890 	:	val_out <= 4'h68c3;
         4'hf891 	:	val_out <= 4'h68c3;
         4'hf892 	:	val_out <= 4'h68c3;
         4'hf893 	:	val_out <= 4'h68c3;
         4'hf898 	:	val_out <= 4'h68dc;
         4'hf899 	:	val_out <= 4'h68dc;
         4'hf89a 	:	val_out <= 4'h68dc;
         4'hf89b 	:	val_out <= 4'h68dc;
         4'hf8a0 	:	val_out <= 4'h68f5;
         4'hf8a1 	:	val_out <= 4'h68f5;
         4'hf8a2 	:	val_out <= 4'h68f5;
         4'hf8a3 	:	val_out <= 4'h68f5;
         4'hf8a8 	:	val_out <= 4'h690d;
         4'hf8a9 	:	val_out <= 4'h690d;
         4'hf8aa 	:	val_out <= 4'h690d;
         4'hf8ab 	:	val_out <= 4'h690d;
         4'hf8b0 	:	val_out <= 4'h6926;
         4'hf8b1 	:	val_out <= 4'h6926;
         4'hf8b2 	:	val_out <= 4'h6926;
         4'hf8b3 	:	val_out <= 4'h6926;
         4'hf8b8 	:	val_out <= 4'h693f;
         4'hf8b9 	:	val_out <= 4'h693f;
         4'hf8ba 	:	val_out <= 4'h693f;
         4'hf8bb 	:	val_out <= 4'h693f;
         4'hf8c0 	:	val_out <= 4'h6957;
         4'hf8c1 	:	val_out <= 4'h6957;
         4'hf8c2 	:	val_out <= 4'h6957;
         4'hf8c3 	:	val_out <= 4'h6957;
         4'hf8c8 	:	val_out <= 4'h6970;
         4'hf8c9 	:	val_out <= 4'h6970;
         4'hf8ca 	:	val_out <= 4'h6970;
         4'hf8cb 	:	val_out <= 4'h6970;
         4'hf8d0 	:	val_out <= 4'h6989;
         4'hf8d1 	:	val_out <= 4'h6989;
         4'hf8d2 	:	val_out <= 4'h6989;
         4'hf8d3 	:	val_out <= 4'h6989;
         4'hf8d8 	:	val_out <= 4'h69a2;
         4'hf8d9 	:	val_out <= 4'h69a2;
         4'hf8da 	:	val_out <= 4'h69a2;
         4'hf8db 	:	val_out <= 4'h69a2;
         4'hf8e0 	:	val_out <= 4'h69ba;
         4'hf8e1 	:	val_out <= 4'h69ba;
         4'hf8e2 	:	val_out <= 4'h69ba;
         4'hf8e3 	:	val_out <= 4'h69ba;
         4'hf8e8 	:	val_out <= 4'h69d3;
         4'hf8e9 	:	val_out <= 4'h69d3;
         4'hf8ea 	:	val_out <= 4'h69d3;
         4'hf8eb 	:	val_out <= 4'h69d3;
         4'hf8f0 	:	val_out <= 4'h69ec;
         4'hf8f1 	:	val_out <= 4'h69ec;
         4'hf8f2 	:	val_out <= 4'h69ec;
         4'hf8f3 	:	val_out <= 4'h69ec;
         4'hf8f8 	:	val_out <= 4'h6a05;
         4'hf8f9 	:	val_out <= 4'h6a05;
         4'hf8fa 	:	val_out <= 4'h6a05;
         4'hf8fb 	:	val_out <= 4'h6a05;
         4'hf900 	:	val_out <= 4'h6a1d;
         4'hf901 	:	val_out <= 4'h6a1d;
         4'hf902 	:	val_out <= 4'h6a1d;
         4'hf903 	:	val_out <= 4'h6a1d;
         4'hf908 	:	val_out <= 4'h6a36;
         4'hf909 	:	val_out <= 4'h6a36;
         4'hf90a 	:	val_out <= 4'h6a36;
         4'hf90b 	:	val_out <= 4'h6a36;
         4'hf910 	:	val_out <= 4'h6a4f;
         4'hf911 	:	val_out <= 4'h6a4f;
         4'hf912 	:	val_out <= 4'h6a4f;
         4'hf913 	:	val_out <= 4'h6a4f;
         4'hf918 	:	val_out <= 4'h6a68;
         4'hf919 	:	val_out <= 4'h6a68;
         4'hf91a 	:	val_out <= 4'h6a68;
         4'hf91b 	:	val_out <= 4'h6a68;
         4'hf920 	:	val_out <= 4'h6a80;
         4'hf921 	:	val_out <= 4'h6a80;
         4'hf922 	:	val_out <= 4'h6a80;
         4'hf923 	:	val_out <= 4'h6a80;
         4'hf928 	:	val_out <= 4'h6a99;
         4'hf929 	:	val_out <= 4'h6a99;
         4'hf92a 	:	val_out <= 4'h6a99;
         4'hf92b 	:	val_out <= 4'h6a99;
         4'hf930 	:	val_out <= 4'h6ab2;
         4'hf931 	:	val_out <= 4'h6ab2;
         4'hf932 	:	val_out <= 4'h6ab2;
         4'hf933 	:	val_out <= 4'h6ab2;
         4'hf938 	:	val_out <= 4'h6acb;
         4'hf939 	:	val_out <= 4'h6acb;
         4'hf93a 	:	val_out <= 4'h6acb;
         4'hf93b 	:	val_out <= 4'h6acb;
         4'hf940 	:	val_out <= 4'h6ae4;
         4'hf941 	:	val_out <= 4'h6ae4;
         4'hf942 	:	val_out <= 4'h6ae4;
         4'hf943 	:	val_out <= 4'h6ae4;
         4'hf948 	:	val_out <= 4'h6afc;
         4'hf949 	:	val_out <= 4'h6afc;
         4'hf94a 	:	val_out <= 4'h6afc;
         4'hf94b 	:	val_out <= 4'h6afc;
         4'hf950 	:	val_out <= 4'h6b15;
         4'hf951 	:	val_out <= 4'h6b15;
         4'hf952 	:	val_out <= 4'h6b15;
         4'hf953 	:	val_out <= 4'h6b15;
         4'hf958 	:	val_out <= 4'h6b2e;
         4'hf959 	:	val_out <= 4'h6b2e;
         4'hf95a 	:	val_out <= 4'h6b2e;
         4'hf95b 	:	val_out <= 4'h6b2e;
         4'hf960 	:	val_out <= 4'h6b47;
         4'hf961 	:	val_out <= 4'h6b47;
         4'hf962 	:	val_out <= 4'h6b47;
         4'hf963 	:	val_out <= 4'h6b47;
         4'hf968 	:	val_out <= 4'h6b60;
         4'hf969 	:	val_out <= 4'h6b60;
         4'hf96a 	:	val_out <= 4'h6b60;
         4'hf96b 	:	val_out <= 4'h6b60;
         4'hf970 	:	val_out <= 4'h6b78;
         4'hf971 	:	val_out <= 4'h6b78;
         4'hf972 	:	val_out <= 4'h6b78;
         4'hf973 	:	val_out <= 4'h6b78;
         4'hf978 	:	val_out <= 4'h6b91;
         4'hf979 	:	val_out <= 4'h6b91;
         4'hf97a 	:	val_out <= 4'h6b91;
         4'hf97b 	:	val_out <= 4'h6b91;
         4'hf980 	:	val_out <= 4'h6baa;
         4'hf981 	:	val_out <= 4'h6baa;
         4'hf982 	:	val_out <= 4'h6baa;
         4'hf983 	:	val_out <= 4'h6baa;
         4'hf988 	:	val_out <= 4'h6bc3;
         4'hf989 	:	val_out <= 4'h6bc3;
         4'hf98a 	:	val_out <= 4'h6bc3;
         4'hf98b 	:	val_out <= 4'h6bc3;
         4'hf990 	:	val_out <= 4'h6bdc;
         4'hf991 	:	val_out <= 4'h6bdc;
         4'hf992 	:	val_out <= 4'h6bdc;
         4'hf993 	:	val_out <= 4'h6bdc;
         4'hf998 	:	val_out <= 4'h6bf4;
         4'hf999 	:	val_out <= 4'h6bf4;
         4'hf99a 	:	val_out <= 4'h6bf4;
         4'hf99b 	:	val_out <= 4'h6bf4;
         4'hf9a0 	:	val_out <= 4'h6c0d;
         4'hf9a1 	:	val_out <= 4'h6c0d;
         4'hf9a2 	:	val_out <= 4'h6c0d;
         4'hf9a3 	:	val_out <= 4'h6c0d;
         4'hf9a8 	:	val_out <= 4'h6c26;
         4'hf9a9 	:	val_out <= 4'h6c26;
         4'hf9aa 	:	val_out <= 4'h6c26;
         4'hf9ab 	:	val_out <= 4'h6c26;
         4'hf9b0 	:	val_out <= 4'h6c3f;
         4'hf9b1 	:	val_out <= 4'h6c3f;
         4'hf9b2 	:	val_out <= 4'h6c3f;
         4'hf9b3 	:	val_out <= 4'h6c3f;
         4'hf9b8 	:	val_out <= 4'h6c58;
         4'hf9b9 	:	val_out <= 4'h6c58;
         4'hf9ba 	:	val_out <= 4'h6c58;
         4'hf9bb 	:	val_out <= 4'h6c58;
         4'hf9c0 	:	val_out <= 4'h6c71;
         4'hf9c1 	:	val_out <= 4'h6c71;
         4'hf9c2 	:	val_out <= 4'h6c71;
         4'hf9c3 	:	val_out <= 4'h6c71;
         4'hf9c8 	:	val_out <= 4'h6c89;
         4'hf9c9 	:	val_out <= 4'h6c89;
         4'hf9ca 	:	val_out <= 4'h6c89;
         4'hf9cb 	:	val_out <= 4'h6c89;
         4'hf9d0 	:	val_out <= 4'h6ca2;
         4'hf9d1 	:	val_out <= 4'h6ca2;
         4'hf9d2 	:	val_out <= 4'h6ca2;
         4'hf9d3 	:	val_out <= 4'h6ca2;
         4'hf9d8 	:	val_out <= 4'h6cbb;
         4'hf9d9 	:	val_out <= 4'h6cbb;
         4'hf9da 	:	val_out <= 4'h6cbb;
         4'hf9db 	:	val_out <= 4'h6cbb;
         4'hf9e0 	:	val_out <= 4'h6cd4;
         4'hf9e1 	:	val_out <= 4'h6cd4;
         4'hf9e2 	:	val_out <= 4'h6cd4;
         4'hf9e3 	:	val_out <= 4'h6cd4;
         4'hf9e8 	:	val_out <= 4'h6ced;
         4'hf9e9 	:	val_out <= 4'h6ced;
         4'hf9ea 	:	val_out <= 4'h6ced;
         4'hf9eb 	:	val_out <= 4'h6ced;
         4'hf9f0 	:	val_out <= 4'h6d06;
         4'hf9f1 	:	val_out <= 4'h6d06;
         4'hf9f2 	:	val_out <= 4'h6d06;
         4'hf9f3 	:	val_out <= 4'h6d06;
         4'hf9f8 	:	val_out <= 4'h6d1f;
         4'hf9f9 	:	val_out <= 4'h6d1f;
         4'hf9fa 	:	val_out <= 4'h6d1f;
         4'hf9fb 	:	val_out <= 4'h6d1f;
         4'hfa00 	:	val_out <= 4'h6d37;
         4'hfa01 	:	val_out <= 4'h6d37;
         4'hfa02 	:	val_out <= 4'h6d37;
         4'hfa03 	:	val_out <= 4'h6d37;
         4'hfa08 	:	val_out <= 4'h6d50;
         4'hfa09 	:	val_out <= 4'h6d50;
         4'hfa0a 	:	val_out <= 4'h6d50;
         4'hfa0b 	:	val_out <= 4'h6d50;
         4'hfa10 	:	val_out <= 4'h6d69;
         4'hfa11 	:	val_out <= 4'h6d69;
         4'hfa12 	:	val_out <= 4'h6d69;
         4'hfa13 	:	val_out <= 4'h6d69;
         4'hfa18 	:	val_out <= 4'h6d82;
         4'hfa19 	:	val_out <= 4'h6d82;
         4'hfa1a 	:	val_out <= 4'h6d82;
         4'hfa1b 	:	val_out <= 4'h6d82;
         4'hfa20 	:	val_out <= 4'h6d9b;
         4'hfa21 	:	val_out <= 4'h6d9b;
         4'hfa22 	:	val_out <= 4'h6d9b;
         4'hfa23 	:	val_out <= 4'h6d9b;
         4'hfa28 	:	val_out <= 4'h6db4;
         4'hfa29 	:	val_out <= 4'h6db4;
         4'hfa2a 	:	val_out <= 4'h6db4;
         4'hfa2b 	:	val_out <= 4'h6db4;
         4'hfa30 	:	val_out <= 4'h6dcd;
         4'hfa31 	:	val_out <= 4'h6dcd;
         4'hfa32 	:	val_out <= 4'h6dcd;
         4'hfa33 	:	val_out <= 4'h6dcd;
         4'hfa38 	:	val_out <= 4'h6de6;
         4'hfa39 	:	val_out <= 4'h6de6;
         4'hfa3a 	:	val_out <= 4'h6de6;
         4'hfa3b 	:	val_out <= 4'h6de6;
         4'hfa40 	:	val_out <= 4'h6dfe;
         4'hfa41 	:	val_out <= 4'h6dfe;
         4'hfa42 	:	val_out <= 4'h6dfe;
         4'hfa43 	:	val_out <= 4'h6dfe;
         4'hfa48 	:	val_out <= 4'h6e17;
         4'hfa49 	:	val_out <= 4'h6e17;
         4'hfa4a 	:	val_out <= 4'h6e17;
         4'hfa4b 	:	val_out <= 4'h6e17;
         4'hfa50 	:	val_out <= 4'h6e30;
         4'hfa51 	:	val_out <= 4'h6e30;
         4'hfa52 	:	val_out <= 4'h6e30;
         4'hfa53 	:	val_out <= 4'h6e30;
         4'hfa58 	:	val_out <= 4'h6e49;
         4'hfa59 	:	val_out <= 4'h6e49;
         4'hfa5a 	:	val_out <= 4'h6e49;
         4'hfa5b 	:	val_out <= 4'h6e49;
         4'hfa60 	:	val_out <= 4'h6e62;
         4'hfa61 	:	val_out <= 4'h6e62;
         4'hfa62 	:	val_out <= 4'h6e62;
         4'hfa63 	:	val_out <= 4'h6e62;
         4'hfa68 	:	val_out <= 4'h6e7b;
         4'hfa69 	:	val_out <= 4'h6e7b;
         4'hfa6a 	:	val_out <= 4'h6e7b;
         4'hfa6b 	:	val_out <= 4'h6e7b;
         4'hfa70 	:	val_out <= 4'h6e94;
         4'hfa71 	:	val_out <= 4'h6e94;
         4'hfa72 	:	val_out <= 4'h6e94;
         4'hfa73 	:	val_out <= 4'h6e94;
         4'hfa78 	:	val_out <= 4'h6ead;
         4'hfa79 	:	val_out <= 4'h6ead;
         4'hfa7a 	:	val_out <= 4'h6ead;
         4'hfa7b 	:	val_out <= 4'h6ead;
         4'hfa80 	:	val_out <= 4'h6ec6;
         4'hfa81 	:	val_out <= 4'h6ec6;
         4'hfa82 	:	val_out <= 4'h6ec6;
         4'hfa83 	:	val_out <= 4'h6ec6;
         4'hfa88 	:	val_out <= 4'h6ede;
         4'hfa89 	:	val_out <= 4'h6ede;
         4'hfa8a 	:	val_out <= 4'h6ede;
         4'hfa8b 	:	val_out <= 4'h6ede;
         4'hfa90 	:	val_out <= 4'h6ef7;
         4'hfa91 	:	val_out <= 4'h6ef7;
         4'hfa92 	:	val_out <= 4'h6ef7;
         4'hfa93 	:	val_out <= 4'h6ef7;
         4'hfa98 	:	val_out <= 4'h6f10;
         4'hfa99 	:	val_out <= 4'h6f10;
         4'hfa9a 	:	val_out <= 4'h6f10;
         4'hfa9b 	:	val_out <= 4'h6f10;
         4'hfaa0 	:	val_out <= 4'h6f29;
         4'hfaa1 	:	val_out <= 4'h6f29;
         4'hfaa2 	:	val_out <= 4'h6f29;
         4'hfaa3 	:	val_out <= 4'h6f29;
         4'hfaa8 	:	val_out <= 4'h6f42;
         4'hfaa9 	:	val_out <= 4'h6f42;
         4'hfaaa 	:	val_out <= 4'h6f42;
         4'hfaab 	:	val_out <= 4'h6f42;
         4'hfab0 	:	val_out <= 4'h6f5b;
         4'hfab1 	:	val_out <= 4'h6f5b;
         4'hfab2 	:	val_out <= 4'h6f5b;
         4'hfab3 	:	val_out <= 4'h6f5b;
         4'hfab8 	:	val_out <= 4'h6f74;
         4'hfab9 	:	val_out <= 4'h6f74;
         4'hfaba 	:	val_out <= 4'h6f74;
         4'hfabb 	:	val_out <= 4'h6f74;
         4'hfac0 	:	val_out <= 4'h6f8d;
         4'hfac1 	:	val_out <= 4'h6f8d;
         4'hfac2 	:	val_out <= 4'h6f8d;
         4'hfac3 	:	val_out <= 4'h6f8d;
         4'hfac8 	:	val_out <= 4'h6fa6;
         4'hfac9 	:	val_out <= 4'h6fa6;
         4'hfaca 	:	val_out <= 4'h6fa6;
         4'hfacb 	:	val_out <= 4'h6fa6;
         4'hfad0 	:	val_out <= 4'h6fbf;
         4'hfad1 	:	val_out <= 4'h6fbf;
         4'hfad2 	:	val_out <= 4'h6fbf;
         4'hfad3 	:	val_out <= 4'h6fbf;
         4'hfad8 	:	val_out <= 4'h6fd8;
         4'hfad9 	:	val_out <= 4'h6fd8;
         4'hfada 	:	val_out <= 4'h6fd8;
         4'hfadb 	:	val_out <= 4'h6fd8;
         4'hfae0 	:	val_out <= 4'h6ff1;
         4'hfae1 	:	val_out <= 4'h6ff1;
         4'hfae2 	:	val_out <= 4'h6ff1;
         4'hfae3 	:	val_out <= 4'h6ff1;
         4'hfae8 	:	val_out <= 4'h700a;
         4'hfae9 	:	val_out <= 4'h700a;
         4'hfaea 	:	val_out <= 4'h700a;
         4'hfaeb 	:	val_out <= 4'h700a;
         4'hfaf0 	:	val_out <= 4'h7022;
         4'hfaf1 	:	val_out <= 4'h7022;
         4'hfaf2 	:	val_out <= 4'h7022;
         4'hfaf3 	:	val_out <= 4'h7022;
         4'hfaf8 	:	val_out <= 4'h703b;
         4'hfaf9 	:	val_out <= 4'h703b;
         4'hfafa 	:	val_out <= 4'h703b;
         4'hfafb 	:	val_out <= 4'h703b;
         4'hfb00 	:	val_out <= 4'h7054;
         4'hfb01 	:	val_out <= 4'h7054;
         4'hfb02 	:	val_out <= 4'h7054;
         4'hfb03 	:	val_out <= 4'h7054;
         4'hfb08 	:	val_out <= 4'h706d;
         4'hfb09 	:	val_out <= 4'h706d;
         4'hfb0a 	:	val_out <= 4'h706d;
         4'hfb0b 	:	val_out <= 4'h706d;
         4'hfb10 	:	val_out <= 4'h7086;
         4'hfb11 	:	val_out <= 4'h7086;
         4'hfb12 	:	val_out <= 4'h7086;
         4'hfb13 	:	val_out <= 4'h7086;
         4'hfb18 	:	val_out <= 4'h709f;
         4'hfb19 	:	val_out <= 4'h709f;
         4'hfb1a 	:	val_out <= 4'h709f;
         4'hfb1b 	:	val_out <= 4'h709f;
         4'hfb20 	:	val_out <= 4'h70b8;
         4'hfb21 	:	val_out <= 4'h70b8;
         4'hfb22 	:	val_out <= 4'h70b8;
         4'hfb23 	:	val_out <= 4'h70b8;
         4'hfb28 	:	val_out <= 4'h70d1;
         4'hfb29 	:	val_out <= 4'h70d1;
         4'hfb2a 	:	val_out <= 4'h70d1;
         4'hfb2b 	:	val_out <= 4'h70d1;
         4'hfb30 	:	val_out <= 4'h70ea;
         4'hfb31 	:	val_out <= 4'h70ea;
         4'hfb32 	:	val_out <= 4'h70ea;
         4'hfb33 	:	val_out <= 4'h70ea;
         4'hfb38 	:	val_out <= 4'h7103;
         4'hfb39 	:	val_out <= 4'h7103;
         4'hfb3a 	:	val_out <= 4'h7103;
         4'hfb3b 	:	val_out <= 4'h7103;
         4'hfb40 	:	val_out <= 4'h711c;
         4'hfb41 	:	val_out <= 4'h711c;
         4'hfb42 	:	val_out <= 4'h711c;
         4'hfb43 	:	val_out <= 4'h711c;
         4'hfb48 	:	val_out <= 4'h7135;
         4'hfb49 	:	val_out <= 4'h7135;
         4'hfb4a 	:	val_out <= 4'h7135;
         4'hfb4b 	:	val_out <= 4'h7135;
         4'hfb50 	:	val_out <= 4'h714e;
         4'hfb51 	:	val_out <= 4'h714e;
         4'hfb52 	:	val_out <= 4'h714e;
         4'hfb53 	:	val_out <= 4'h714e;
         4'hfb58 	:	val_out <= 4'h7167;
         4'hfb59 	:	val_out <= 4'h7167;
         4'hfb5a 	:	val_out <= 4'h7167;
         4'hfb5b 	:	val_out <= 4'h7167;
         4'hfb60 	:	val_out <= 4'h7180;
         4'hfb61 	:	val_out <= 4'h7180;
         4'hfb62 	:	val_out <= 4'h7180;
         4'hfb63 	:	val_out <= 4'h7180;
         4'hfb68 	:	val_out <= 4'h7199;
         4'hfb69 	:	val_out <= 4'h7199;
         4'hfb6a 	:	val_out <= 4'h7199;
         4'hfb6b 	:	val_out <= 4'h7199;
         4'hfb70 	:	val_out <= 4'h71b2;
         4'hfb71 	:	val_out <= 4'h71b2;
         4'hfb72 	:	val_out <= 4'h71b2;
         4'hfb73 	:	val_out <= 4'h71b2;
         4'hfb78 	:	val_out <= 4'h71cb;
         4'hfb79 	:	val_out <= 4'h71cb;
         4'hfb7a 	:	val_out <= 4'h71cb;
         4'hfb7b 	:	val_out <= 4'h71cb;
         4'hfb80 	:	val_out <= 4'h71e4;
         4'hfb81 	:	val_out <= 4'h71e4;
         4'hfb82 	:	val_out <= 4'h71e4;
         4'hfb83 	:	val_out <= 4'h71e4;
         4'hfb88 	:	val_out <= 4'h71fd;
         4'hfb89 	:	val_out <= 4'h71fd;
         4'hfb8a 	:	val_out <= 4'h71fd;
         4'hfb8b 	:	val_out <= 4'h71fd;
         4'hfb90 	:	val_out <= 4'h7216;
         4'hfb91 	:	val_out <= 4'h7216;
         4'hfb92 	:	val_out <= 4'h7216;
         4'hfb93 	:	val_out <= 4'h7216;
         4'hfb98 	:	val_out <= 4'h722f;
         4'hfb99 	:	val_out <= 4'h722f;
         4'hfb9a 	:	val_out <= 4'h722f;
         4'hfb9b 	:	val_out <= 4'h722f;
         4'hfba0 	:	val_out <= 4'h7248;
         4'hfba1 	:	val_out <= 4'h7248;
         4'hfba2 	:	val_out <= 4'h7248;
         4'hfba3 	:	val_out <= 4'h7248;
         4'hfba8 	:	val_out <= 4'h7261;
         4'hfba9 	:	val_out <= 4'h7261;
         4'hfbaa 	:	val_out <= 4'h7261;
         4'hfbab 	:	val_out <= 4'h7261;
         4'hfbb0 	:	val_out <= 4'h727a;
         4'hfbb1 	:	val_out <= 4'h727a;
         4'hfbb2 	:	val_out <= 4'h727a;
         4'hfbb3 	:	val_out <= 4'h727a;
         4'hfbb8 	:	val_out <= 4'h7293;
         4'hfbb9 	:	val_out <= 4'h7293;
         4'hfbba 	:	val_out <= 4'h7293;
         4'hfbbb 	:	val_out <= 4'h7293;
         4'hfbc0 	:	val_out <= 4'h72ac;
         4'hfbc1 	:	val_out <= 4'h72ac;
         4'hfbc2 	:	val_out <= 4'h72ac;
         4'hfbc3 	:	val_out <= 4'h72ac;
         4'hfbc8 	:	val_out <= 4'h72c5;
         4'hfbc9 	:	val_out <= 4'h72c5;
         4'hfbca 	:	val_out <= 4'h72c5;
         4'hfbcb 	:	val_out <= 4'h72c5;
         4'hfbd0 	:	val_out <= 4'h72de;
         4'hfbd1 	:	val_out <= 4'h72de;
         4'hfbd2 	:	val_out <= 4'h72de;
         4'hfbd3 	:	val_out <= 4'h72de;
         4'hfbd8 	:	val_out <= 4'h72f7;
         4'hfbd9 	:	val_out <= 4'h72f7;
         4'hfbda 	:	val_out <= 4'h72f7;
         4'hfbdb 	:	val_out <= 4'h72f7;
         4'hfbe0 	:	val_out <= 4'h7310;
         4'hfbe1 	:	val_out <= 4'h7310;
         4'hfbe2 	:	val_out <= 4'h7310;
         4'hfbe3 	:	val_out <= 4'h7310;
         4'hfbe8 	:	val_out <= 4'h7329;
         4'hfbe9 	:	val_out <= 4'h7329;
         4'hfbea 	:	val_out <= 4'h7329;
         4'hfbeb 	:	val_out <= 4'h7329;
         4'hfbf0 	:	val_out <= 4'h7342;
         4'hfbf1 	:	val_out <= 4'h7342;
         4'hfbf2 	:	val_out <= 4'h7342;
         4'hfbf3 	:	val_out <= 4'h7342;
         4'hfbf8 	:	val_out <= 4'h735b;
         4'hfbf9 	:	val_out <= 4'h735b;
         4'hfbfa 	:	val_out <= 4'h735b;
         4'hfbfb 	:	val_out <= 4'h735b;
         4'hfc00 	:	val_out <= 4'h7374;
         4'hfc01 	:	val_out <= 4'h7374;
         4'hfc02 	:	val_out <= 4'h7374;
         4'hfc03 	:	val_out <= 4'h7374;
         4'hfc08 	:	val_out <= 4'h738d;
         4'hfc09 	:	val_out <= 4'h738d;
         4'hfc0a 	:	val_out <= 4'h738d;
         4'hfc0b 	:	val_out <= 4'h738d;
         4'hfc10 	:	val_out <= 4'h73a6;
         4'hfc11 	:	val_out <= 4'h73a6;
         4'hfc12 	:	val_out <= 4'h73a6;
         4'hfc13 	:	val_out <= 4'h73a6;
         4'hfc18 	:	val_out <= 4'h73bf;
         4'hfc19 	:	val_out <= 4'h73bf;
         4'hfc1a 	:	val_out <= 4'h73bf;
         4'hfc1b 	:	val_out <= 4'h73bf;
         4'hfc20 	:	val_out <= 4'h73d8;
         4'hfc21 	:	val_out <= 4'h73d8;
         4'hfc22 	:	val_out <= 4'h73d8;
         4'hfc23 	:	val_out <= 4'h73d8;
         4'hfc28 	:	val_out <= 4'h73f1;
         4'hfc29 	:	val_out <= 4'h73f1;
         4'hfc2a 	:	val_out <= 4'h73f1;
         4'hfc2b 	:	val_out <= 4'h73f1;
         4'hfc30 	:	val_out <= 4'h740a;
         4'hfc31 	:	val_out <= 4'h740a;
         4'hfc32 	:	val_out <= 4'h740a;
         4'hfc33 	:	val_out <= 4'h740a;
         4'hfc38 	:	val_out <= 4'h7423;
         4'hfc39 	:	val_out <= 4'h7423;
         4'hfc3a 	:	val_out <= 4'h7423;
         4'hfc3b 	:	val_out <= 4'h7423;
         4'hfc40 	:	val_out <= 4'h743c;
         4'hfc41 	:	val_out <= 4'h743c;
         4'hfc42 	:	val_out <= 4'h743c;
         4'hfc43 	:	val_out <= 4'h743c;
         4'hfc48 	:	val_out <= 4'h7455;
         4'hfc49 	:	val_out <= 4'h7455;
         4'hfc4a 	:	val_out <= 4'h7455;
         4'hfc4b 	:	val_out <= 4'h7455;
         4'hfc50 	:	val_out <= 4'h746e;
         4'hfc51 	:	val_out <= 4'h746e;
         4'hfc52 	:	val_out <= 4'h746e;
         4'hfc53 	:	val_out <= 4'h746e;
         4'hfc58 	:	val_out <= 4'h7487;
         4'hfc59 	:	val_out <= 4'h7487;
         4'hfc5a 	:	val_out <= 4'h7487;
         4'hfc5b 	:	val_out <= 4'h7487;
         4'hfc60 	:	val_out <= 4'h74a0;
         4'hfc61 	:	val_out <= 4'h74a0;
         4'hfc62 	:	val_out <= 4'h74a0;
         4'hfc63 	:	val_out <= 4'h74a0;
         4'hfc68 	:	val_out <= 4'h74b9;
         4'hfc69 	:	val_out <= 4'h74b9;
         4'hfc6a 	:	val_out <= 4'h74b9;
         4'hfc6b 	:	val_out <= 4'h74b9;
         4'hfc70 	:	val_out <= 4'h74d2;
         4'hfc71 	:	val_out <= 4'h74d2;
         4'hfc72 	:	val_out <= 4'h74d2;
         4'hfc73 	:	val_out <= 4'h74d2;
         4'hfc78 	:	val_out <= 4'h74eb;
         4'hfc79 	:	val_out <= 4'h74eb;
         4'hfc7a 	:	val_out <= 4'h74eb;
         4'hfc7b 	:	val_out <= 4'h74eb;
         4'hfc80 	:	val_out <= 4'h7504;
         4'hfc81 	:	val_out <= 4'h7504;
         4'hfc82 	:	val_out <= 4'h7504;
         4'hfc83 	:	val_out <= 4'h7504;
         4'hfc88 	:	val_out <= 4'h751d;
         4'hfc89 	:	val_out <= 4'h751d;
         4'hfc8a 	:	val_out <= 4'h751d;
         4'hfc8b 	:	val_out <= 4'h751d;
         4'hfc90 	:	val_out <= 4'h7536;
         4'hfc91 	:	val_out <= 4'h7536;
         4'hfc92 	:	val_out <= 4'h7536;
         4'hfc93 	:	val_out <= 4'h7536;
         4'hfc98 	:	val_out <= 4'h754f;
         4'hfc99 	:	val_out <= 4'h754f;
         4'hfc9a 	:	val_out <= 4'h754f;
         4'hfc9b 	:	val_out <= 4'h754f;
         4'hfca0 	:	val_out <= 4'h7568;
         4'hfca1 	:	val_out <= 4'h7568;
         4'hfca2 	:	val_out <= 4'h7568;
         4'hfca3 	:	val_out <= 4'h7568;
         4'hfca8 	:	val_out <= 4'h7581;
         4'hfca9 	:	val_out <= 4'h7581;
         4'hfcaa 	:	val_out <= 4'h7581;
         4'hfcab 	:	val_out <= 4'h7581;
         4'hfcb0 	:	val_out <= 4'h759a;
         4'hfcb1 	:	val_out <= 4'h759a;
         4'hfcb2 	:	val_out <= 4'h759a;
         4'hfcb3 	:	val_out <= 4'h759a;
         4'hfcb8 	:	val_out <= 4'h75b3;
         4'hfcb9 	:	val_out <= 4'h75b3;
         4'hfcba 	:	val_out <= 4'h75b3;
         4'hfcbb 	:	val_out <= 4'h75b3;
         4'hfcc0 	:	val_out <= 4'h75cc;
         4'hfcc1 	:	val_out <= 4'h75cc;
         4'hfcc2 	:	val_out <= 4'h75cc;
         4'hfcc3 	:	val_out <= 4'h75cc;
         4'hfcc8 	:	val_out <= 4'h75e6;
         4'hfcc9 	:	val_out <= 4'h75e6;
         4'hfcca 	:	val_out <= 4'h75e6;
         4'hfccb 	:	val_out <= 4'h75e6;
         4'hfcd0 	:	val_out <= 4'h75ff;
         4'hfcd1 	:	val_out <= 4'h75ff;
         4'hfcd2 	:	val_out <= 4'h75ff;
         4'hfcd3 	:	val_out <= 4'h75ff;
         4'hfcd8 	:	val_out <= 4'h7618;
         4'hfcd9 	:	val_out <= 4'h7618;
         4'hfcda 	:	val_out <= 4'h7618;
         4'hfcdb 	:	val_out <= 4'h7618;
         4'hfce0 	:	val_out <= 4'h7631;
         4'hfce1 	:	val_out <= 4'h7631;
         4'hfce2 	:	val_out <= 4'h7631;
         4'hfce3 	:	val_out <= 4'h7631;
         4'hfce8 	:	val_out <= 4'h764a;
         4'hfce9 	:	val_out <= 4'h764a;
         4'hfcea 	:	val_out <= 4'h764a;
         4'hfceb 	:	val_out <= 4'h764a;
         4'hfcf0 	:	val_out <= 4'h7663;
         4'hfcf1 	:	val_out <= 4'h7663;
         4'hfcf2 	:	val_out <= 4'h7663;
         4'hfcf3 	:	val_out <= 4'h7663;
         4'hfcf8 	:	val_out <= 4'h767c;
         4'hfcf9 	:	val_out <= 4'h767c;
         4'hfcfa 	:	val_out <= 4'h767c;
         4'hfcfb 	:	val_out <= 4'h767c;
         4'hfd00 	:	val_out <= 4'h7695;
         4'hfd01 	:	val_out <= 4'h7695;
         4'hfd02 	:	val_out <= 4'h7695;
         4'hfd03 	:	val_out <= 4'h7695;
         4'hfd08 	:	val_out <= 4'h76ae;
         4'hfd09 	:	val_out <= 4'h76ae;
         4'hfd0a 	:	val_out <= 4'h76ae;
         4'hfd0b 	:	val_out <= 4'h76ae;
         4'hfd10 	:	val_out <= 4'h76c7;
         4'hfd11 	:	val_out <= 4'h76c7;
         4'hfd12 	:	val_out <= 4'h76c7;
         4'hfd13 	:	val_out <= 4'h76c7;
         4'hfd18 	:	val_out <= 4'h76e0;
         4'hfd19 	:	val_out <= 4'h76e0;
         4'hfd1a 	:	val_out <= 4'h76e0;
         4'hfd1b 	:	val_out <= 4'h76e0;
         4'hfd20 	:	val_out <= 4'h76f9;
         4'hfd21 	:	val_out <= 4'h76f9;
         4'hfd22 	:	val_out <= 4'h76f9;
         4'hfd23 	:	val_out <= 4'h76f9;
         4'hfd28 	:	val_out <= 4'h7712;
         4'hfd29 	:	val_out <= 4'h7712;
         4'hfd2a 	:	val_out <= 4'h7712;
         4'hfd2b 	:	val_out <= 4'h7712;
         4'hfd30 	:	val_out <= 4'h772b;
         4'hfd31 	:	val_out <= 4'h772b;
         4'hfd32 	:	val_out <= 4'h772b;
         4'hfd33 	:	val_out <= 4'h772b;
         4'hfd38 	:	val_out <= 4'h7744;
         4'hfd39 	:	val_out <= 4'h7744;
         4'hfd3a 	:	val_out <= 4'h7744;
         4'hfd3b 	:	val_out <= 4'h7744;
         4'hfd40 	:	val_out <= 4'h775d;
         4'hfd41 	:	val_out <= 4'h775d;
         4'hfd42 	:	val_out <= 4'h775d;
         4'hfd43 	:	val_out <= 4'h775d;
         4'hfd48 	:	val_out <= 4'h7777;
         4'hfd49 	:	val_out <= 4'h7777;
         4'hfd4a 	:	val_out <= 4'h7777;
         4'hfd4b 	:	val_out <= 4'h7777;
         4'hfd50 	:	val_out <= 4'h7790;
         4'hfd51 	:	val_out <= 4'h7790;
         4'hfd52 	:	val_out <= 4'h7790;
         4'hfd53 	:	val_out <= 4'h7790;
         4'hfd58 	:	val_out <= 4'h77a9;
         4'hfd59 	:	val_out <= 4'h77a9;
         4'hfd5a 	:	val_out <= 4'h77a9;
         4'hfd5b 	:	val_out <= 4'h77a9;
         4'hfd60 	:	val_out <= 4'h77c2;
         4'hfd61 	:	val_out <= 4'h77c2;
         4'hfd62 	:	val_out <= 4'h77c2;
         4'hfd63 	:	val_out <= 4'h77c2;
         4'hfd68 	:	val_out <= 4'h77db;
         4'hfd69 	:	val_out <= 4'h77db;
         4'hfd6a 	:	val_out <= 4'h77db;
         4'hfd6b 	:	val_out <= 4'h77db;
         4'hfd70 	:	val_out <= 4'h77f4;
         4'hfd71 	:	val_out <= 4'h77f4;
         4'hfd72 	:	val_out <= 4'h77f4;
         4'hfd73 	:	val_out <= 4'h77f4;
         4'hfd78 	:	val_out <= 4'h780d;
         4'hfd79 	:	val_out <= 4'h780d;
         4'hfd7a 	:	val_out <= 4'h780d;
         4'hfd7b 	:	val_out <= 4'h780d;
         4'hfd80 	:	val_out <= 4'h7826;
         4'hfd81 	:	val_out <= 4'h7826;
         4'hfd82 	:	val_out <= 4'h7826;
         4'hfd83 	:	val_out <= 4'h7826;
         4'hfd88 	:	val_out <= 4'h783f;
         4'hfd89 	:	val_out <= 4'h783f;
         4'hfd8a 	:	val_out <= 4'h783f;
         4'hfd8b 	:	val_out <= 4'h783f;
         4'hfd90 	:	val_out <= 4'h7858;
         4'hfd91 	:	val_out <= 4'h7858;
         4'hfd92 	:	val_out <= 4'h7858;
         4'hfd93 	:	val_out <= 4'h7858;
         4'hfd98 	:	val_out <= 4'h7871;
         4'hfd99 	:	val_out <= 4'h7871;
         4'hfd9a 	:	val_out <= 4'h7871;
         4'hfd9b 	:	val_out <= 4'h7871;
         4'hfda0 	:	val_out <= 4'h788a;
         4'hfda1 	:	val_out <= 4'h788a;
         4'hfda2 	:	val_out <= 4'h788a;
         4'hfda3 	:	val_out <= 4'h788a;
         4'hfda8 	:	val_out <= 4'h78a4;
         4'hfda9 	:	val_out <= 4'h78a4;
         4'hfdaa 	:	val_out <= 4'h78a4;
         4'hfdab 	:	val_out <= 4'h78a4;
         4'hfdb0 	:	val_out <= 4'h78bd;
         4'hfdb1 	:	val_out <= 4'h78bd;
         4'hfdb2 	:	val_out <= 4'h78bd;
         4'hfdb3 	:	val_out <= 4'h78bd;
         4'hfdb8 	:	val_out <= 4'h78d6;
         4'hfdb9 	:	val_out <= 4'h78d6;
         4'hfdba 	:	val_out <= 4'h78d6;
         4'hfdbb 	:	val_out <= 4'h78d6;
         4'hfdc0 	:	val_out <= 4'h78ef;
         4'hfdc1 	:	val_out <= 4'h78ef;
         4'hfdc2 	:	val_out <= 4'h78ef;
         4'hfdc3 	:	val_out <= 4'h78ef;
         4'hfdc8 	:	val_out <= 4'h7908;
         4'hfdc9 	:	val_out <= 4'h7908;
         4'hfdca 	:	val_out <= 4'h7908;
         4'hfdcb 	:	val_out <= 4'h7908;
         4'hfdd0 	:	val_out <= 4'h7921;
         4'hfdd1 	:	val_out <= 4'h7921;
         4'hfdd2 	:	val_out <= 4'h7921;
         4'hfdd3 	:	val_out <= 4'h7921;
         4'hfdd8 	:	val_out <= 4'h793a;
         4'hfdd9 	:	val_out <= 4'h793a;
         4'hfdda 	:	val_out <= 4'h793a;
         4'hfddb 	:	val_out <= 4'h793a;
         4'hfde0 	:	val_out <= 4'h7953;
         4'hfde1 	:	val_out <= 4'h7953;
         4'hfde2 	:	val_out <= 4'h7953;
         4'hfde3 	:	val_out <= 4'h7953;
         4'hfde8 	:	val_out <= 4'h796c;
         4'hfde9 	:	val_out <= 4'h796c;
         4'hfdea 	:	val_out <= 4'h796c;
         4'hfdeb 	:	val_out <= 4'h796c;
         4'hfdf0 	:	val_out <= 4'h7985;
         4'hfdf1 	:	val_out <= 4'h7985;
         4'hfdf2 	:	val_out <= 4'h7985;
         4'hfdf3 	:	val_out <= 4'h7985;
         4'hfdf8 	:	val_out <= 4'h799f;
         4'hfdf9 	:	val_out <= 4'h799f;
         4'hfdfa 	:	val_out <= 4'h799f;
         4'hfdfb 	:	val_out <= 4'h799f;
         4'hfe00 	:	val_out <= 4'h79b8;
         4'hfe01 	:	val_out <= 4'h79b8;
         4'hfe02 	:	val_out <= 4'h79b8;
         4'hfe03 	:	val_out <= 4'h79b8;
         4'hfe08 	:	val_out <= 4'h79d1;
         4'hfe09 	:	val_out <= 4'h79d1;
         4'hfe0a 	:	val_out <= 4'h79d1;
         4'hfe0b 	:	val_out <= 4'h79d1;
         4'hfe10 	:	val_out <= 4'h79ea;
         4'hfe11 	:	val_out <= 4'h79ea;
         4'hfe12 	:	val_out <= 4'h79ea;
         4'hfe13 	:	val_out <= 4'h79ea;
         4'hfe18 	:	val_out <= 4'h7a03;
         4'hfe19 	:	val_out <= 4'h7a03;
         4'hfe1a 	:	val_out <= 4'h7a03;
         4'hfe1b 	:	val_out <= 4'h7a03;
         4'hfe20 	:	val_out <= 4'h7a1c;
         4'hfe21 	:	val_out <= 4'h7a1c;
         4'hfe22 	:	val_out <= 4'h7a1c;
         4'hfe23 	:	val_out <= 4'h7a1c;
         4'hfe28 	:	val_out <= 4'h7a35;
         4'hfe29 	:	val_out <= 4'h7a35;
         4'hfe2a 	:	val_out <= 4'h7a35;
         4'hfe2b 	:	val_out <= 4'h7a35;
         4'hfe30 	:	val_out <= 4'h7a4e;
         4'hfe31 	:	val_out <= 4'h7a4e;
         4'hfe32 	:	val_out <= 4'h7a4e;
         4'hfe33 	:	val_out <= 4'h7a4e;
         4'hfe38 	:	val_out <= 4'h7a67;
         4'hfe39 	:	val_out <= 4'h7a67;
         4'hfe3a 	:	val_out <= 4'h7a67;
         4'hfe3b 	:	val_out <= 4'h7a67;
         4'hfe40 	:	val_out <= 4'h7a80;
         4'hfe41 	:	val_out <= 4'h7a80;
         4'hfe42 	:	val_out <= 4'h7a80;
         4'hfe43 	:	val_out <= 4'h7a80;
         4'hfe48 	:	val_out <= 4'h7a9a;
         4'hfe49 	:	val_out <= 4'h7a9a;
         4'hfe4a 	:	val_out <= 4'h7a9a;
         4'hfe4b 	:	val_out <= 4'h7a9a;
         4'hfe50 	:	val_out <= 4'h7ab3;
         4'hfe51 	:	val_out <= 4'h7ab3;
         4'hfe52 	:	val_out <= 4'h7ab3;
         4'hfe53 	:	val_out <= 4'h7ab3;
         4'hfe58 	:	val_out <= 4'h7acc;
         4'hfe59 	:	val_out <= 4'h7acc;
         4'hfe5a 	:	val_out <= 4'h7acc;
         4'hfe5b 	:	val_out <= 4'h7acc;
         4'hfe60 	:	val_out <= 4'h7ae5;
         4'hfe61 	:	val_out <= 4'h7ae5;
         4'hfe62 	:	val_out <= 4'h7ae5;
         4'hfe63 	:	val_out <= 4'h7ae5;
         4'hfe68 	:	val_out <= 4'h7afe;
         4'hfe69 	:	val_out <= 4'h7afe;
         4'hfe6a 	:	val_out <= 4'h7afe;
         4'hfe6b 	:	val_out <= 4'h7afe;
         4'hfe70 	:	val_out <= 4'h7b17;
         4'hfe71 	:	val_out <= 4'h7b17;
         4'hfe72 	:	val_out <= 4'h7b17;
         4'hfe73 	:	val_out <= 4'h7b17;
         4'hfe78 	:	val_out <= 4'h7b30;
         4'hfe79 	:	val_out <= 4'h7b30;
         4'hfe7a 	:	val_out <= 4'h7b30;
         4'hfe7b 	:	val_out <= 4'h7b30;
         4'hfe80 	:	val_out <= 4'h7b49;
         4'hfe81 	:	val_out <= 4'h7b49;
         4'hfe82 	:	val_out <= 4'h7b49;
         4'hfe83 	:	val_out <= 4'h7b49;
         4'hfe88 	:	val_out <= 4'h7b63;
         4'hfe89 	:	val_out <= 4'h7b63;
         4'hfe8a 	:	val_out <= 4'h7b63;
         4'hfe8b 	:	val_out <= 4'h7b63;
         4'hfe90 	:	val_out <= 4'h7b7c;
         4'hfe91 	:	val_out <= 4'h7b7c;
         4'hfe92 	:	val_out <= 4'h7b7c;
         4'hfe93 	:	val_out <= 4'h7b7c;
         4'hfe98 	:	val_out <= 4'h7b95;
         4'hfe99 	:	val_out <= 4'h7b95;
         4'hfe9a 	:	val_out <= 4'h7b95;
         4'hfe9b 	:	val_out <= 4'h7b95;
         4'hfea0 	:	val_out <= 4'h7bae;
         4'hfea1 	:	val_out <= 4'h7bae;
         4'hfea2 	:	val_out <= 4'h7bae;
         4'hfea3 	:	val_out <= 4'h7bae;
         4'hfea8 	:	val_out <= 4'h7bc7;
         4'hfea9 	:	val_out <= 4'h7bc7;
         4'hfeaa 	:	val_out <= 4'h7bc7;
         4'hfeab 	:	val_out <= 4'h7bc7;
         4'hfeb0 	:	val_out <= 4'h7be0;
         4'hfeb1 	:	val_out <= 4'h7be0;
         4'hfeb2 	:	val_out <= 4'h7be0;
         4'hfeb3 	:	val_out <= 4'h7be0;
         4'hfeb8 	:	val_out <= 4'h7bf9;
         4'hfeb9 	:	val_out <= 4'h7bf9;
         4'hfeba 	:	val_out <= 4'h7bf9;
         4'hfebb 	:	val_out <= 4'h7bf9;
         4'hfec0 	:	val_out <= 4'h7c12;
         4'hfec1 	:	val_out <= 4'h7c12;
         4'hfec2 	:	val_out <= 4'h7c12;
         4'hfec3 	:	val_out <= 4'h7c12;
         4'hfec8 	:	val_out <= 4'h7c2b;
         4'hfec9 	:	val_out <= 4'h7c2b;
         4'hfeca 	:	val_out <= 4'h7c2b;
         4'hfecb 	:	val_out <= 4'h7c2b;
         4'hfed0 	:	val_out <= 4'h7c45;
         4'hfed1 	:	val_out <= 4'h7c45;
         4'hfed2 	:	val_out <= 4'h7c45;
         4'hfed3 	:	val_out <= 4'h7c45;
         4'hfed8 	:	val_out <= 4'h7c5e;
         4'hfed9 	:	val_out <= 4'h7c5e;
         4'hfeda 	:	val_out <= 4'h7c5e;
         4'hfedb 	:	val_out <= 4'h7c5e;
         4'hfee0 	:	val_out <= 4'h7c77;
         4'hfee1 	:	val_out <= 4'h7c77;
         4'hfee2 	:	val_out <= 4'h7c77;
         4'hfee3 	:	val_out <= 4'h7c77;
         4'hfee8 	:	val_out <= 4'h7c90;
         4'hfee9 	:	val_out <= 4'h7c90;
         4'hfeea 	:	val_out <= 4'h7c90;
         4'hfeeb 	:	val_out <= 4'h7c90;
         4'hfef0 	:	val_out <= 4'h7ca9;
         4'hfef1 	:	val_out <= 4'h7ca9;
         4'hfef2 	:	val_out <= 4'h7ca9;
         4'hfef3 	:	val_out <= 4'h7ca9;
         4'hfef8 	:	val_out <= 4'h7cc2;
         4'hfef9 	:	val_out <= 4'h7cc2;
         4'hfefa 	:	val_out <= 4'h7cc2;
         4'hfefb 	:	val_out <= 4'h7cc2;
         4'hff00 	:	val_out <= 4'h7cdb;
         4'hff01 	:	val_out <= 4'h7cdb;
         4'hff02 	:	val_out <= 4'h7cdb;
         4'hff03 	:	val_out <= 4'h7cdb;
         4'hff08 	:	val_out <= 4'h7cf4;
         4'hff09 	:	val_out <= 4'h7cf4;
         4'hff0a 	:	val_out <= 4'h7cf4;
         4'hff0b 	:	val_out <= 4'h7cf4;
         4'hff10 	:	val_out <= 4'h7d0e;
         4'hff11 	:	val_out <= 4'h7d0e;
         4'hff12 	:	val_out <= 4'h7d0e;
         4'hff13 	:	val_out <= 4'h7d0e;
         4'hff18 	:	val_out <= 4'h7d27;
         4'hff19 	:	val_out <= 4'h7d27;
         4'hff1a 	:	val_out <= 4'h7d27;
         4'hff1b 	:	val_out <= 4'h7d27;
         4'hff20 	:	val_out <= 4'h7d40;
         4'hff21 	:	val_out <= 4'h7d40;
         4'hff22 	:	val_out <= 4'h7d40;
         4'hff23 	:	val_out <= 4'h7d40;
         4'hff28 	:	val_out <= 4'h7d59;
         4'hff29 	:	val_out <= 4'h7d59;
         4'hff2a 	:	val_out <= 4'h7d59;
         4'hff2b 	:	val_out <= 4'h7d59;
         4'hff30 	:	val_out <= 4'h7d72;
         4'hff31 	:	val_out <= 4'h7d72;
         4'hff32 	:	val_out <= 4'h7d72;
         4'hff33 	:	val_out <= 4'h7d72;
         4'hff38 	:	val_out <= 4'h7d8b;
         4'hff39 	:	val_out <= 4'h7d8b;
         4'hff3a 	:	val_out <= 4'h7d8b;
         4'hff3b 	:	val_out <= 4'h7d8b;
         4'hff40 	:	val_out <= 4'h7da4;
         4'hff41 	:	val_out <= 4'h7da4;
         4'hff42 	:	val_out <= 4'h7da4;
         4'hff43 	:	val_out <= 4'h7da4;
         4'hff48 	:	val_out <= 4'h7dbd;
         4'hff49 	:	val_out <= 4'h7dbd;
         4'hff4a 	:	val_out <= 4'h7dbd;
         4'hff4b 	:	val_out <= 4'h7dbd;
         4'hff50 	:	val_out <= 4'h7dd7;
         4'hff51 	:	val_out <= 4'h7dd7;
         4'hff52 	:	val_out <= 4'h7dd7;
         4'hff53 	:	val_out <= 4'h7dd7;
         4'hff58 	:	val_out <= 4'h7df0;
         4'hff59 	:	val_out <= 4'h7df0;
         4'hff5a 	:	val_out <= 4'h7df0;
         4'hff5b 	:	val_out <= 4'h7df0;
         4'hff60 	:	val_out <= 4'h7e09;
         4'hff61 	:	val_out <= 4'h7e09;
         4'hff62 	:	val_out <= 4'h7e09;
         4'hff63 	:	val_out <= 4'h7e09;
         4'hff68 	:	val_out <= 4'h7e22;
         4'hff69 	:	val_out <= 4'h7e22;
         4'hff6a 	:	val_out <= 4'h7e22;
         4'hff6b 	:	val_out <= 4'h7e22;
         4'hff70 	:	val_out <= 4'h7e3b;
         4'hff71 	:	val_out <= 4'h7e3b;
         4'hff72 	:	val_out <= 4'h7e3b;
         4'hff73 	:	val_out <= 4'h7e3b;
         4'hff78 	:	val_out <= 4'h7e54;
         4'hff79 	:	val_out <= 4'h7e54;
         4'hff7a 	:	val_out <= 4'h7e54;
         4'hff7b 	:	val_out <= 4'h7e54;
         4'hff80 	:	val_out <= 4'h7e6d;
         4'hff81 	:	val_out <= 4'h7e6d;
         4'hff82 	:	val_out <= 4'h7e6d;
         4'hff83 	:	val_out <= 4'h7e6d;
         4'hff88 	:	val_out <= 4'h7e87;
         4'hff89 	:	val_out <= 4'h7e87;
         4'hff8a 	:	val_out <= 4'h7e87;
         4'hff8b 	:	val_out <= 4'h7e87;
         4'hff90 	:	val_out <= 4'h7ea0;
         4'hff91 	:	val_out <= 4'h7ea0;
         4'hff92 	:	val_out <= 4'h7ea0;
         4'hff93 	:	val_out <= 4'h7ea0;
         4'hff98 	:	val_out <= 4'h7eb9;
         4'hff99 	:	val_out <= 4'h7eb9;
         4'hff9a 	:	val_out <= 4'h7eb9;
         4'hff9b 	:	val_out <= 4'h7eb9;
         4'hffa0 	:	val_out <= 4'h7ed2;
         4'hffa1 	:	val_out <= 4'h7ed2;
         4'hffa2 	:	val_out <= 4'h7ed2;
         4'hffa3 	:	val_out <= 4'h7ed2;
         4'hffa8 	:	val_out <= 4'h7eeb;
         4'hffa9 	:	val_out <= 4'h7eeb;
         4'hffaa 	:	val_out <= 4'h7eeb;
         4'hffab 	:	val_out <= 4'h7eeb;
         4'hffb0 	:	val_out <= 4'h7f04;
         4'hffb1 	:	val_out <= 4'h7f04;
         4'hffb2 	:	val_out <= 4'h7f04;
         4'hffb3 	:	val_out <= 4'h7f04;
         4'hffb8 	:	val_out <= 4'h7f1d;
         4'hffb9 	:	val_out <= 4'h7f1d;
         4'hffba 	:	val_out <= 4'h7f1d;
         4'hffbb 	:	val_out <= 4'h7f1d;
         4'hffc0 	:	val_out <= 4'h7f36;
         4'hffc1 	:	val_out <= 4'h7f36;
         4'hffc2 	:	val_out <= 4'h7f36;
         4'hffc3 	:	val_out <= 4'h7f36;
         4'hffc8 	:	val_out <= 4'h7f50;
         4'hffc9 	:	val_out <= 4'h7f50;
         4'hffca 	:	val_out <= 4'h7f50;
         4'hffcb 	:	val_out <= 4'h7f50;
         4'hffd0 	:	val_out <= 4'h7f69;
         4'hffd1 	:	val_out <= 4'h7f69;
         4'hffd2 	:	val_out <= 4'h7f69;
         4'hffd3 	:	val_out <= 4'h7f69;
         4'hffd8 	:	val_out <= 4'h7f82;
         4'hffd9 	:	val_out <= 4'h7f82;
         4'hffda 	:	val_out <= 4'h7f82;
         4'hffdb 	:	val_out <= 4'h7f82;
         4'hffe0 	:	val_out <= 4'h7f9b;
         4'hffe1 	:	val_out <= 4'h7f9b;
         4'hffe2 	:	val_out <= 4'h7f9b;
         4'hffe3 	:	val_out <= 4'h7f9b;
         4'hffe8 	:	val_out <= 4'h7fb4;
         4'hffe9 	:	val_out <= 4'h7fb4;
         4'hffea 	:	val_out <= 4'h7fb4;
         4'hffeb 	:	val_out <= 4'h7fb4;
         4'hfff0 	:	val_out <= 4'h7fcd;
         4'hfff1 	:	val_out <= 4'h7fcd;
         4'hfff2 	:	val_out <= 4'h7fcd;
         4'hfff3 	:	val_out <= 4'h7fcd;
         4'hfff8 	:	val_out <= 4'h7fe6;
         4'hfff9 	:	val_out <= 4'h7fe6;
         4'hfffa 	:	val_out <= 4'h7fe6;
         4'hfffb 	:	val_out <= 4'h7fe6;
			default	:	val_out <= 4'h0000;
		endcase
	end
endmodule
