// Pipelined phase bank module

module phase_bank_p(input clk,
						input clk_en,
						input rst,
						input[6:0] i_midi,
						output reg[6:0] o_midi,
						output reg o_valid, 
						output reg[23:0] o_phase);
		parameter NBANKS = 10;
		
		// for now holding 24 bits, feeding LUT with only 16 upper bits of bank -> losing precision but frequency should be right
		// if want make phase interpolation then need to output both integer and fractional part then interpolate in sine
		reg[23:0] phase_banks[NBANKS-1:0];
		wire[23:0] w_tw;
		
		tuning_word_lut tw_lut(.i_midi(i_midi), .o_tw(w_tw));
		
		integer v_idx;
		integer i;
		
		initial begin
			o_phase = 16'b0;
			v_idx = 9;
			for (i = 0; i < NBANKS; i = i + 1) begin
				phase_banks[i] = 24'b0;
			end
			o_midi = 7'b0;
		end
		
		always @(posedge clk or posedge rst) begin
			if (rst) begin
				o_phase = 16'b0;
				v_idx = 9;
				for (i = 0; i < NBANKS; i = i + 1) begin
					phase_banks[i] <= 24'b0;
				end
				o_midi <= 7'b0;
			end else if (clk_en) begin
				if (i_midi !== 7'h0) begin
					phase_banks[v_idx] <= phase_banks[v_idx] + w_tw;
					o_phase <= phase_banks[v_idx]; // output a delayed value (one whole loop)
				end else begin
					o_phase <= 16'b0;
				end
					
				o_valid <= (i_midi == 7'h0) ? 1'b0 : 1'b1;
				o_midi <= i_midi;
				
				if (v_idx == NBANKS - 1)
					v_idx <= 0;
				else
					v_idx <= v_idx + 1;
			end
		end
						
endmodule

// right now increasing tw to 24 bits
module tuning_word_lut(input[6:0] i_midi,
								output reg[23:0] o_tw);
		initial o_tw = 24'b0;
		
		always @(i_midi) begin
			case(i_midi)
            7'h00 	:	o_tw <= 24'b000000000000010110010100;
            7'h01 	:	o_tw <= 24'b000000000000010111101001;
            7'h02 	:	o_tw <= 24'b000000000000011001000011;
            7'h03 	:	o_tw <= 24'b000000000000011010100011;
            7'h04 	:	o_tw <= 24'b000000000000011100001000;
            7'h05 	:	o_tw <= 24'b000000000000011101110011;
            7'h06 	:	o_tw <= 24'b000000000000011111100100;
            7'h07 	:	o_tw <= 24'b000000000000100001011100;
            7'h08 	:	o_tw <= 24'b000000000000100011011100;
            7'h09 	:	o_tw <= 24'b000000000000100101100010;
            7'h0a 	:	o_tw <= 24'b000000000000100111110001;
            7'h0b 	:	o_tw <= 24'b000000000000101010001001;
            7'h0c 	:	o_tw <= 24'b000000000000101100101001;
            7'h0d 	:	o_tw <= 24'b000000000000101111010011;
            7'h0e 	:	o_tw <= 24'b000000000000110010000111;
            7'h0f 	:	o_tw <= 24'b000000000000110101000110;
            7'h10 	:	o_tw <= 24'b000000000000111000010000;
            7'h11 	:	o_tw <= 24'b000000000000111011100110;
            7'h12 	:	o_tw <= 24'b000000000000111111001001;
            7'h13 	:	o_tw <= 24'b000000000001000010111001;
            7'h14 	:	o_tw <= 24'b000000000001000110111000;
            7'h15 	:	o_tw <= 24'b000000000001001011000101;
            7'h16 	:	o_tw <= 24'b000000000001001111100011;
            7'h17 	:	o_tw <= 24'b000000000001010100010010;
            7'h18 	:	o_tw <= 24'b000000000001011001010011;
            7'h19 	:	o_tw <= 24'b000000000001011110100111;
            7'h1a 	:	o_tw <= 24'b000000000001100100001111;
            7'h1b 	:	o_tw <= 24'b000000000001101010001100;
            7'h1c 	:	o_tw <= 24'b000000000001110000100000;
            7'h1d 	:	o_tw <= 24'b000000000001110111001101;
            7'h1e 	:	o_tw <= 24'b000000000001111110010010;
            7'h1f 	:	o_tw <= 24'b000000000010000101110011;
            7'h20 	:	o_tw <= 24'b000000000010001101110000;
            7'h21 	:	o_tw <= 24'b000000000010010110001011;
            7'h22 	:	o_tw <= 24'b000000000010011111000111;
            7'h23 	:	o_tw <= 24'b000000000010101000100101;
            7'h24 	:	o_tw <= 24'b000000000010110010100110;
            7'h25 	:	o_tw <= 24'b000000000010111101001110;
            7'h26 	:	o_tw <= 24'b000000000011001000011110;
            7'h27 	:	o_tw <= 24'b000000000011010100011001;
            7'h28 	:	o_tw <= 24'b000000000011100001000001;
            7'h29 	:	o_tw <= 24'b000000000011101110011010;
            7'h2a 	:	o_tw <= 24'b000000000011111100100101;
            7'h2b 	:	o_tw <= 24'b000000000100001011100110;
            7'h2c 	:	o_tw <= 24'b000000000100011011100000;
            7'h2d 	:	o_tw <= 24'b000000000100101100010111;
            7'h2e 	:	o_tw <= 24'b000000000100111110001111;
            7'h2f 	:	o_tw <= 24'b000000000101010001001010;
            7'h30 	:	o_tw <= 24'b000000000101100101001101;
            7'h31 	:	o_tw <= 24'b000000000101111010011100;
            7'h32 	:	o_tw <= 24'b000000000110010000111100;
            7'h33 	:	o_tw <= 24'b000000000110101000110010;
            7'h34 	:	o_tw <= 24'b000000000111000010000011;
            7'h35 	:	o_tw <= 24'b000000000111011100110100;
            7'h36 	:	o_tw <= 24'b000000000111111001001010;
            7'h37 	:	o_tw <= 24'b000000001000010111001101;
            7'h38 	:	o_tw <= 24'b000000001000110111000001;
            7'h39 	:	o_tw <= 24'b000000001001011000101111;
            7'h3a 	:	o_tw <= 24'b000000001001111100011110;
            7'h3b 	:	o_tw <= 24'b000000001010100010010100;
            7'h3c 	:	o_tw <= 24'b000000001011001010011010;
            7'h3d 	:	o_tw <= 24'b000000001011110100111001;
            7'h3e 	:	o_tw <= 24'b000000001100100001111001;
            7'h3f 	:	o_tw <= 24'b000000001101010001100101;
            7'h40 	:	o_tw <= 24'b000000001110000100000110;
            7'h41 	:	o_tw <= 24'b000000001110111001101000;
            7'h42 	:	o_tw <= 24'b000000001111110010010101;
            7'h43 	:	o_tw <= 24'b000000010000101110011010;
            7'h44 	:	o_tw <= 24'b000000010001101110000011;
            7'h45 	:	o_tw <= 24'b000000010010110001011111;
            7'h46 	:	o_tw <= 24'b000000010011111000111100;
            7'h47 	:	o_tw <= 24'b000000010101000100101000;
            7'h48 	:	o_tw <= 24'b000000010110010100110100;
            7'h49 	:	o_tw <= 24'b000000010111101001110010;
            7'h4a 	:	o_tw <= 24'b000000011001000011110011;
            7'h4b 	:	o_tw <= 24'b000000011010100011001010;
            7'h4c 	:	o_tw <= 24'b000000011100001000001101;
            7'h4d 	:	o_tw <= 24'b000000011101110011010000;
            7'h4e 	:	o_tw <= 24'b000000011111100100101010;
            7'h4f 	:	o_tw <= 24'b000000100001011100110100;
            7'h50 	:	o_tw <= 24'b000000100011011100000111;
            7'h51 	:	o_tw <= 24'b000000100101100010111111;
            7'h52 	:	o_tw <= 24'b000000100111110001111000;
            7'h53 	:	o_tw <= 24'b000000101010001001010000;
            7'h54 	:	o_tw <= 24'b000000101100101001101001;
            7'h55 	:	o_tw <= 24'b000000101111010011100100;
            7'h56 	:	o_tw <= 24'b000000110010000111100110;
            7'h57 	:	o_tw <= 24'b000000110101000110010101;
            7'h58 	:	o_tw <= 24'b000000111000010000011010;
            7'h59 	:	o_tw <= 24'b000000111011100110100000;
            7'h5a 	:	o_tw <= 24'b000000111111001001010100;
            7'h5b 	:	o_tw <= 24'b000001000010111001101000;
            7'h5c 	:	o_tw <= 24'b000001000110111000001111;
            7'h5d 	:	o_tw <= 24'b000001001011000101111110;
            7'h5e 	:	o_tw <= 24'b000001001111100011110000;
            7'h5f 	:	o_tw <= 24'b000001010100010010100001;
            7'h60 	:	o_tw <= 24'b000001011001010011010011;
            7'h61 	:	o_tw <= 24'b000001011110100111001001;
            7'h62 	:	o_tw <= 24'b000001100100001111001101;
            7'h63 	:	o_tw <= 24'b000001101010001100101011;
            7'h64 	:	o_tw <= 24'b000001110000100000110100;
            7'h65 	:	o_tw <= 24'b000001110111001101000000;
            7'h66 	:	o_tw <= 24'b000001111110010010101001;
            7'h67 	:	o_tw <= 24'b000010000101110011010001;
            7'h68 	:	o_tw <= 24'b000010001101110000011110;
            7'h69 	:	o_tw <= 24'b000010010110001011111100;
            7'h6a 	:	o_tw <= 24'b000010011111000111100000;
            7'h6b 	:	o_tw <= 24'b000010101000100101000010;
            7'h6c 	:	o_tw <= 24'b000010110010100110100110;
            7'h6d 	:	o_tw <= 24'b000010111101001110010010;
            7'h6e 	:	o_tw <= 24'b000011001000011110011010;
            7'h6f 	:	o_tw <= 24'b000011010100011001010110;
            7'h70 	:	o_tw <= 24'b000011100001000001101001;
            7'h71 	:	o_tw <= 24'b000011101110011010000000;
            7'h72 	:	o_tw <= 24'b000011111100100101010011;
            7'h73 	:	o_tw <= 24'b000100001011100110100010;
            7'h74 	:	o_tw <= 24'b000100011011100000111100;
            7'h75 	:	o_tw <= 24'b000100101100010111111001;
            7'h76 	:	o_tw <= 24'b000100111110001111000000;
            7'h77 	:	o_tw <= 24'b000101010001001010000101;
            7'h78 	:	o_tw <= 24'b000101100101001101001100;
            7'h79 	:	o_tw <= 24'b000101111010011100100101;
            7'h7a 	:	o_tw <= 24'b000110010000111100110100;
            7'h7b 	:	o_tw <= 24'b000110101000110010101100;
            7'h7c 	:	o_tw <= 24'b000111000010000011010010;
            7'h7d 	:	o_tw <= 24'b000111011100110100000001;
            7'h7e 	:	o_tw <= 24'b000111111001001010100110;
            7'h7f 	:	o_tw <= 24'b001000010111001101000101;
				default 	:	o_tw <= 24'h0000; // h00 is MIDI 0 value
			endcase
		end	
endmodule
