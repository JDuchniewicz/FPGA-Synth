

module quarter_sine_lut(input[13:0] i_phase,
								output reg signed[15:0] o_val); //is reg needed here? try removing
		always @(i_phase) begin
			case(i_phase)
                14'h000 	:	o_val <= 16'b0000000000000110;
                14'h001 	:	o_val <= 16'b0000000000010010;
                14'h002 	:	o_val <= 16'b0000000000011111;
                14'h003 	:	o_val <= 16'b0000000000101011;
                14'h004 	:	o_val <= 16'b0000000000111000;
                14'h005 	:	o_val <= 16'b0000000001000101;
                14'h006 	:	o_val <= 16'b0000000001010001;
                14'h007 	:	o_val <= 16'b0000000001011110;
                14'h008 	:	o_val <= 16'b0000000001101010;
                14'h009 	:	o_val <= 16'b0000000001110111;
                14'h00a 	:	o_val <= 16'b0000000010000011;
                14'h00b 	:	o_val <= 16'b0000000010010000;
                14'h00c 	:	o_val <= 16'b0000000010011101;
                14'h00d 	:	o_val <= 16'b0000000010101001;
                14'h00e 	:	o_val <= 16'b0000000010110110;
                14'h00f 	:	o_val <= 16'b0000000011000010;
                14'h010 	:	o_val <= 16'b0000000011001111;
                14'h011 	:	o_val <= 16'b0000000011011011;
                14'h012 	:	o_val <= 16'b0000000011101000;
                14'h013 	:	o_val <= 16'b0000000011110101;
                14'h014 	:	o_val <= 16'b0000000100000001;
                14'h015 	:	o_val <= 16'b0000000100001110;
                14'h016 	:	o_val <= 16'b0000000100011010;
                14'h017 	:	o_val <= 16'b0000000100100111;
                14'h018 	:	o_val <= 16'b0000000100110011;
                14'h019 	:	o_val <= 16'b0000000101000000;
                14'h01a 	:	o_val <= 16'b0000000101001101;
                14'h01b 	:	o_val <= 16'b0000000101011001;
                14'h01c 	:	o_val <= 16'b0000000101100110;
                14'h01d 	:	o_val <= 16'b0000000101110010;
                14'h01e 	:	o_val <= 16'b0000000101111111;
                14'h01f 	:	o_val <= 16'b0000000110001011;
                14'h020 	:	o_val <= 16'b0000000110011000;
                14'h021 	:	o_val <= 16'b0000000110100100;
                14'h022 	:	o_val <= 16'b0000000110110001;
                14'h023 	:	o_val <= 16'b0000000110111110;
                14'h024 	:	o_val <= 16'b0000000111001010;
                14'h025 	:	o_val <= 16'b0000000111010111;
                14'h026 	:	o_val <= 16'b0000000111100011;
                14'h027 	:	o_val <= 16'b0000000111110000;
                14'h028 	:	o_val <= 16'b0000000111111100;
                14'h029 	:	o_val <= 16'b0000001000001001;
                14'h02a 	:	o_val <= 16'b0000001000010110;
                14'h02b 	:	o_val <= 16'b0000001000100010;
                14'h02c 	:	o_val <= 16'b0000001000101111;
                14'h02d 	:	o_val <= 16'b0000001000111011;
                14'h02e 	:	o_val <= 16'b0000001001001000;
                14'h02f 	:	o_val <= 16'b0000001001010100;
                14'h030 	:	o_val <= 16'b0000001001100001;
                14'h031 	:	o_val <= 16'b0000001001101101;
                14'h032 	:	o_val <= 16'b0000001001111010;
                14'h033 	:	o_val <= 16'b0000001010000111;
                14'h034 	:	o_val <= 16'b0000001010010011;
                14'h035 	:	o_val <= 16'b0000001010100000;
                14'h036 	:	o_val <= 16'b0000001010101100;
                14'h037 	:	o_val <= 16'b0000001010111001;
                14'h038 	:	o_val <= 16'b0000001011000101;
                14'h039 	:	o_val <= 16'b0000001011010010;
                14'h03a 	:	o_val <= 16'b0000001011011111;
                14'h03b 	:	o_val <= 16'b0000001011101011;
                14'h03c 	:	o_val <= 16'b0000001011111000;
                14'h03d 	:	o_val <= 16'b0000001100000100;
                14'h03e 	:	o_val <= 16'b0000001100010001;
                14'h03f 	:	o_val <= 16'b0000001100011101;
                14'h040 	:	o_val <= 16'b0000001100101010;
                14'h041 	:	o_val <= 16'b0000001100110111;
                14'h042 	:	o_val <= 16'b0000001101000011;
                14'h043 	:	o_val <= 16'b0000001101010000;
                14'h044 	:	o_val <= 16'b0000001101011100;
                14'h045 	:	o_val <= 16'b0000001101101001;
                14'h046 	:	o_val <= 16'b0000001101110101;
                14'h047 	:	o_val <= 16'b0000001110000010;
                14'h048 	:	o_val <= 16'b0000001110001110;
                14'h049 	:	o_val <= 16'b0000001110011011;
                14'h04a 	:	o_val <= 16'b0000001110101000;
                14'h04b 	:	o_val <= 16'b0000001110110100;
                14'h04c 	:	o_val <= 16'b0000001111000001;
                14'h04d 	:	o_val <= 16'b0000001111001101;
                14'h04e 	:	o_val <= 16'b0000001111011010;
                14'h04f 	:	o_val <= 16'b0000001111100110;
                14'h050 	:	o_val <= 16'b0000001111110011;
                14'h051 	:	o_val <= 16'b0000001111111111;
                14'h052 	:	o_val <= 16'b0000010000001100;
                14'h053 	:	o_val <= 16'b0000010000011001;
                14'h054 	:	o_val <= 16'b0000010000100101;
                14'h055 	:	o_val <= 16'b0000010000110010;
                14'h056 	:	o_val <= 16'b0000010000111110;
                14'h057 	:	o_val <= 16'b0000010001001011;
                14'h058 	:	o_val <= 16'b0000010001010111;
                14'h059 	:	o_val <= 16'b0000010001100100;
                14'h05a 	:	o_val <= 16'b0000010001110001;
                14'h05b 	:	o_val <= 16'b0000010001111101;
                14'h05c 	:	o_val <= 16'b0000010010001010;
                14'h05d 	:	o_val <= 16'b0000010010010110;
                14'h05e 	:	o_val <= 16'b0000010010100011;
                14'h05f 	:	o_val <= 16'b0000010010101111;
                14'h060 	:	o_val <= 16'b0000010010111100;
                14'h061 	:	o_val <= 16'b0000010011001000;
                14'h062 	:	o_val <= 16'b0000010011010101;
                14'h063 	:	o_val <= 16'b0000010011100010;
                14'h064 	:	o_val <= 16'b0000010011101110;
                14'h065 	:	o_val <= 16'b0000010011111011;
                14'h066 	:	o_val <= 16'b0000010100000111;
                14'h067 	:	o_val <= 16'b0000010100010100;
                14'h068 	:	o_val <= 16'b0000010100100000;
                14'h069 	:	o_val <= 16'b0000010100101101;
                14'h06a 	:	o_val <= 16'b0000010100111001;
                14'h06b 	:	o_val <= 16'b0000010101000110;
                14'h06c 	:	o_val <= 16'b0000010101010011;
                14'h06d 	:	o_val <= 16'b0000010101011111;
                14'h06e 	:	o_val <= 16'b0000010101101100;
                14'h06f 	:	o_val <= 16'b0000010101111000;
                14'h070 	:	o_val <= 16'b0000010110000101;
                14'h071 	:	o_val <= 16'b0000010110010001;
                14'h072 	:	o_val <= 16'b0000010110011110;
                14'h073 	:	o_val <= 16'b0000010110101010;
                14'h074 	:	o_val <= 16'b0000010110110111;
                14'h075 	:	o_val <= 16'b0000010111000100;
                14'h076 	:	o_val <= 16'b0000010111010000;
                14'h077 	:	o_val <= 16'b0000010111011101;
                14'h078 	:	o_val <= 16'b0000010111101001;
                14'h079 	:	o_val <= 16'b0000010111110110;
                14'h07a 	:	o_val <= 16'b0000011000000010;
                14'h07b 	:	o_val <= 16'b0000011000001111;
                14'h07c 	:	o_val <= 16'b0000011000011011;
                14'h07d 	:	o_val <= 16'b0000011000101000;
                14'h07e 	:	o_val <= 16'b0000011000110101;
                14'h07f 	:	o_val <= 16'b0000011001000001;
                14'h080 	:	o_val <= 16'b0000011001001110;
                14'h081 	:	o_val <= 16'b0000011001011010;
                14'h082 	:	o_val <= 16'b0000011001100111;
                14'h083 	:	o_val <= 16'b0000011001110011;
                14'h084 	:	o_val <= 16'b0000011010000000;
                14'h085 	:	o_val <= 16'b0000011010001100;
                14'h086 	:	o_val <= 16'b0000011010011001;
                14'h087 	:	o_val <= 16'b0000011010100101;
                14'h088 	:	o_val <= 16'b0000011010110010;
                14'h089 	:	o_val <= 16'b0000011010111111;
                14'h08a 	:	o_val <= 16'b0000011011001011;
                14'h08b 	:	o_val <= 16'b0000011011011000;
                14'h08c 	:	o_val <= 16'b0000011011100100;
                14'h08d 	:	o_val <= 16'b0000011011110001;
                14'h08e 	:	o_val <= 16'b0000011011111101;
                14'h08f 	:	o_val <= 16'b0000011100001010;
                14'h090 	:	o_val <= 16'b0000011100010110;
                14'h091 	:	o_val <= 16'b0000011100100011;
                14'h092 	:	o_val <= 16'b0000011100110000;
                14'h093 	:	o_val <= 16'b0000011100111100;
                14'h094 	:	o_val <= 16'b0000011101001001;
                14'h095 	:	o_val <= 16'b0000011101010101;
                14'h096 	:	o_val <= 16'b0000011101100010;
                14'h097 	:	o_val <= 16'b0000011101101110;
                14'h098 	:	o_val <= 16'b0000011101111011;
                14'h099 	:	o_val <= 16'b0000011110000111;
                14'h09a 	:	o_val <= 16'b0000011110010100;
                14'h09b 	:	o_val <= 16'b0000011110100000;
                14'h09c 	:	o_val <= 16'b0000011110101101;
                14'h09d 	:	o_val <= 16'b0000011110111010;
                14'h09e 	:	o_val <= 16'b0000011111000110;
                14'h09f 	:	o_val <= 16'b0000011111010011;
                14'h0a0 	:	o_val <= 16'b0000011111011111;
                14'h0a1 	:	o_val <= 16'b0000011111101100;
                14'h0a2 	:	o_val <= 16'b0000011111111000;
                14'h0a3 	:	o_val <= 16'b0000100000000101;
                14'h0a4 	:	o_val <= 16'b0000100000010001;
                14'h0a5 	:	o_val <= 16'b0000100000011110;
                14'h0a6 	:	o_val <= 16'b0000100000101010;
                14'h0a7 	:	o_val <= 16'b0000100000110111;
                14'h0a8 	:	o_val <= 16'b0000100001000011;
                14'h0a9 	:	o_val <= 16'b0000100001010000;
                14'h0aa 	:	o_val <= 16'b0000100001011101;
                14'h0ab 	:	o_val <= 16'b0000100001101001;
                14'h0ac 	:	o_val <= 16'b0000100001110110;
                14'h0ad 	:	o_val <= 16'b0000100010000010;
                14'h0ae 	:	o_val <= 16'b0000100010001111;
                14'h0af 	:	o_val <= 16'b0000100010011011;
                14'h0b0 	:	o_val <= 16'b0000100010101000;
                14'h0b1 	:	o_val <= 16'b0000100010110100;
                14'h0b2 	:	o_val <= 16'b0000100011000001;
                14'h0b3 	:	o_val <= 16'b0000100011001101;
                14'h0b4 	:	o_val <= 16'b0000100011011010;
                14'h0b5 	:	o_val <= 16'b0000100011100110;
                14'h0b6 	:	o_val <= 16'b0000100011110011;
                14'h0b7 	:	o_val <= 16'b0000100100000000;
                14'h0b8 	:	o_val <= 16'b0000100100001100;
                14'h0b9 	:	o_val <= 16'b0000100100011001;
                14'h0ba 	:	o_val <= 16'b0000100100100101;
                14'h0bb 	:	o_val <= 16'b0000100100110010;
                14'h0bc 	:	o_val <= 16'b0000100100111110;
                14'h0bd 	:	o_val <= 16'b0000100101001011;
                14'h0be 	:	o_val <= 16'b0000100101010111;
                14'h0bf 	:	o_val <= 16'b0000100101100100;
                14'h0c0 	:	o_val <= 16'b0000100101110000;
                14'h0c1 	:	o_val <= 16'b0000100101111101;
                14'h0c2 	:	o_val <= 16'b0000100110001001;
                14'h0c3 	:	o_val <= 16'b0000100110010110;
                14'h0c4 	:	o_val <= 16'b0000100110100010;
                14'h0c5 	:	o_val <= 16'b0000100110101111;
                14'h0c6 	:	o_val <= 16'b0000100110111100;
                14'h0c7 	:	o_val <= 16'b0000100111001000;
                14'h0c8 	:	o_val <= 16'b0000100111010101;
                14'h0c9 	:	o_val <= 16'b0000100111100001;
                14'h0ca 	:	o_val <= 16'b0000100111101110;
                14'h0cb 	:	o_val <= 16'b0000100111111010;
                14'h0cc 	:	o_val <= 16'b0000101000000111;
                14'h0cd 	:	o_val <= 16'b0000101000010011;
                14'h0ce 	:	o_val <= 16'b0000101000100000;
                14'h0cf 	:	o_val <= 16'b0000101000101100;
                14'h0d0 	:	o_val <= 16'b0000101000111001;
                14'h0d1 	:	o_val <= 16'b0000101001000101;
                14'h0d2 	:	o_val <= 16'b0000101001010010;
                14'h0d3 	:	o_val <= 16'b0000101001011110;
                14'h0d4 	:	o_val <= 16'b0000101001101011;
                14'h0d5 	:	o_val <= 16'b0000101001110111;
                14'h0d6 	:	o_val <= 16'b0000101010000100;
                14'h0d7 	:	o_val <= 16'b0000101010010000;
                14'h0d8 	:	o_val <= 16'b0000101010011101;
                14'h0d9 	:	o_val <= 16'b0000101010101010;
                14'h0da 	:	o_val <= 16'b0000101010110110;
                14'h0db 	:	o_val <= 16'b0000101011000011;
                14'h0dc 	:	o_val <= 16'b0000101011001111;
                14'h0dd 	:	o_val <= 16'b0000101011011100;
                14'h0de 	:	o_val <= 16'b0000101011101000;
                14'h0df 	:	o_val <= 16'b0000101011110101;
                14'h0e0 	:	o_val <= 16'b0000101100000001;
                14'h0e1 	:	o_val <= 16'b0000101100001110;
                14'h0e2 	:	o_val <= 16'b0000101100011010;
                14'h0e3 	:	o_val <= 16'b0000101100100111;
                14'h0e4 	:	o_val <= 16'b0000101100110011;
                14'h0e5 	:	o_val <= 16'b0000101101000000;
                14'h0e6 	:	o_val <= 16'b0000101101001100;
                14'h0e7 	:	o_val <= 16'b0000101101011001;
                14'h0e8 	:	o_val <= 16'b0000101101100101;
                14'h0e9 	:	o_val <= 16'b0000101101110010;
                14'h0ea 	:	o_val <= 16'b0000101101111110;
                14'h0eb 	:	o_val <= 16'b0000101110001011;
                14'h0ec 	:	o_val <= 16'b0000101110010111;
                14'h0ed 	:	o_val <= 16'b0000101110100100;
                14'h0ee 	:	o_val <= 16'b0000101110110000;
                14'h0ef 	:	o_val <= 16'b0000101110111101;
                14'h0f0 	:	o_val <= 16'b0000101111001001;
                14'h0f1 	:	o_val <= 16'b0000101111010110;
                14'h0f2 	:	o_val <= 16'b0000101111100010;
                14'h0f3 	:	o_val <= 16'b0000101111101111;
                14'h0f4 	:	o_val <= 16'b0000101111111011;
                14'h0f5 	:	o_val <= 16'b0000110000001000;
                14'h0f6 	:	o_val <= 16'b0000110000010100;
                14'h0f7 	:	o_val <= 16'b0000110000100001;
                14'h0f8 	:	o_val <= 16'b0000110000101110;
                14'h0f9 	:	o_val <= 16'b0000110000111010;
                14'h0fa 	:	o_val <= 16'b0000110001000111;
                14'h0fb 	:	o_val <= 16'b0000110001010011;
                14'h0fc 	:	o_val <= 16'b0000110001100000;
                14'h0fd 	:	o_val <= 16'b0000110001101100;
                14'h0fe 	:	o_val <= 16'b0000110001111001;
                14'h0ff 	:	o_val <= 16'b0000110010000101;
                14'h100 	:	o_val <= 16'b0000110010010010;
                14'h101 	:	o_val <= 16'b0000110010011110;
                14'h102 	:	o_val <= 16'b0000110010101011;
                14'h103 	:	o_val <= 16'b0000110010110111;
                14'h104 	:	o_val <= 16'b0000110011000100;
                14'h105 	:	o_val <= 16'b0000110011010000;
                14'h106 	:	o_val <= 16'b0000110011011101;
                14'h107 	:	o_val <= 16'b0000110011101001;
                14'h108 	:	o_val <= 16'b0000110011110110;
                14'h109 	:	o_val <= 16'b0000110100000010;
                14'h10a 	:	o_val <= 16'b0000110100001111;
                14'h10b 	:	o_val <= 16'b0000110100011011;
                14'h10c 	:	o_val <= 16'b0000110100101000;
                14'h10d 	:	o_val <= 16'b0000110100110100;
                14'h10e 	:	o_val <= 16'b0000110101000001;
                14'h10f 	:	o_val <= 16'b0000110101001101;
                14'h110 	:	o_val <= 16'b0000110101011010;
                14'h111 	:	o_val <= 16'b0000110101100110;
                14'h112 	:	o_val <= 16'b0000110101110011;
                14'h113 	:	o_val <= 16'b0000110101111111;
                14'h114 	:	o_val <= 16'b0000110110001100;
                14'h115 	:	o_val <= 16'b0000110110011000;
                14'h116 	:	o_val <= 16'b0000110110100101;
                14'h117 	:	o_val <= 16'b0000110110110001;
                14'h118 	:	o_val <= 16'b0000110110111110;
                14'h119 	:	o_val <= 16'b0000110111001010;
                14'h11a 	:	o_val <= 16'b0000110111010111;
                14'h11b 	:	o_val <= 16'b0000110111100011;
                14'h11c 	:	o_val <= 16'b0000110111110000;
                14'h11d 	:	o_val <= 16'b0000110111111100;
                14'h11e 	:	o_val <= 16'b0000111000001001;
                14'h11f 	:	o_val <= 16'b0000111000010101;
                14'h120 	:	o_val <= 16'b0000111000100010;
                14'h121 	:	o_val <= 16'b0000111000101110;
                14'h122 	:	o_val <= 16'b0000111000111010;
                14'h123 	:	o_val <= 16'b0000111001000111;
                14'h124 	:	o_val <= 16'b0000111001010011;
                14'h125 	:	o_val <= 16'b0000111001100000;
                14'h126 	:	o_val <= 16'b0000111001101100;
                14'h127 	:	o_val <= 16'b0000111001111001;
                14'h128 	:	o_val <= 16'b0000111010000101;
                14'h129 	:	o_val <= 16'b0000111010010010;
                14'h12a 	:	o_val <= 16'b0000111010011110;
                14'h12b 	:	o_val <= 16'b0000111010101011;
                14'h12c 	:	o_val <= 16'b0000111010110111;
                14'h12d 	:	o_val <= 16'b0000111011000100;
                14'h12e 	:	o_val <= 16'b0000111011010000;
                14'h12f 	:	o_val <= 16'b0000111011011101;
                14'h130 	:	o_val <= 16'b0000111011101001;
                14'h131 	:	o_val <= 16'b0000111011110110;
                14'h132 	:	o_val <= 16'b0000111100000010;
                14'h133 	:	o_val <= 16'b0000111100001111;
                14'h134 	:	o_val <= 16'b0000111100011011;
                14'h135 	:	o_val <= 16'b0000111100101000;
                14'h136 	:	o_val <= 16'b0000111100110100;
                14'h137 	:	o_val <= 16'b0000111101000001;
                14'h138 	:	o_val <= 16'b0000111101001101;
                14'h139 	:	o_val <= 16'b0000111101011010;
                14'h13a 	:	o_val <= 16'b0000111101100110;
                14'h13b 	:	o_val <= 16'b0000111101110011;
                14'h13c 	:	o_val <= 16'b0000111101111111;
                14'h13d 	:	o_val <= 16'b0000111110001011;
                14'h13e 	:	o_val <= 16'b0000111110011000;
                14'h13f 	:	o_val <= 16'b0000111110100100;
                14'h140 	:	o_val <= 16'b0000111110110001;
                14'h141 	:	o_val <= 16'b0000111110111101;
                14'h142 	:	o_val <= 16'b0000111111001010;
                14'h143 	:	o_val <= 16'b0000111111010110;
                14'h144 	:	o_val <= 16'b0000111111100011;
                14'h145 	:	o_val <= 16'b0000111111101111;
                14'h146 	:	o_val <= 16'b0000111111111100;
                14'h147 	:	o_val <= 16'b0001000000001000;
                14'h148 	:	o_val <= 16'b0001000000010101;
                14'h149 	:	o_val <= 16'b0001000000100001;
                14'h14a 	:	o_val <= 16'b0001000000101110;
                14'h14b 	:	o_val <= 16'b0001000000111010;
                14'h14c 	:	o_val <= 16'b0001000001000111;
                14'h14d 	:	o_val <= 16'b0001000001010011;
                14'h14e 	:	o_val <= 16'b0001000001011111;
                14'h14f 	:	o_val <= 16'b0001000001101100;
                14'h150 	:	o_val <= 16'b0001000001111000;
                14'h151 	:	o_val <= 16'b0001000010000101;
                14'h152 	:	o_val <= 16'b0001000010010001;
                14'h153 	:	o_val <= 16'b0001000010011110;
                14'h154 	:	o_val <= 16'b0001000010101010;
                14'h155 	:	o_val <= 16'b0001000010110111;
                14'h156 	:	o_val <= 16'b0001000011000011;
                14'h157 	:	o_val <= 16'b0001000011010000;
                14'h158 	:	o_val <= 16'b0001000011011100;
                14'h159 	:	o_val <= 16'b0001000011101000;
                14'h15a 	:	o_val <= 16'b0001000011110101;
                14'h15b 	:	o_val <= 16'b0001000100000001;
                14'h15c 	:	o_val <= 16'b0001000100001110;
                14'h15d 	:	o_val <= 16'b0001000100011010;
                14'h15e 	:	o_val <= 16'b0001000100100111;
                14'h15f 	:	o_val <= 16'b0001000100110011;
                14'h160 	:	o_val <= 16'b0001000101000000;
                14'h161 	:	o_val <= 16'b0001000101001100;
                14'h162 	:	o_val <= 16'b0001000101011001;
                14'h163 	:	o_val <= 16'b0001000101100101;
                14'h164 	:	o_val <= 16'b0001000101110001;
                14'h165 	:	o_val <= 16'b0001000101111110;
                14'h166 	:	o_val <= 16'b0001000110001010;
                14'h167 	:	o_val <= 16'b0001000110010111;
                14'h168 	:	o_val <= 16'b0001000110100011;
                14'h169 	:	o_val <= 16'b0001000110110000;
                14'h16a 	:	o_val <= 16'b0001000110111100;
                14'h16b 	:	o_val <= 16'b0001000111001001;
                14'h16c 	:	o_val <= 16'b0001000111010101;
                14'h16d 	:	o_val <= 16'b0001000111100001;
                14'h16e 	:	o_val <= 16'b0001000111101110;
                14'h16f 	:	o_val <= 16'b0001000111111010;
                14'h170 	:	o_val <= 16'b0001001000000111;
                14'h171 	:	o_val <= 16'b0001001000010011;
                14'h172 	:	o_val <= 16'b0001001000100000;
                14'h173 	:	o_val <= 16'b0001001000101100;
                14'h174 	:	o_val <= 16'b0001001000111001;
                14'h175 	:	o_val <= 16'b0001001001000101;
                14'h176 	:	o_val <= 16'b0001001001010001;
                14'h177 	:	o_val <= 16'b0001001001011110;
                14'h178 	:	o_val <= 16'b0001001001101010;
                14'h179 	:	o_val <= 16'b0001001001110111;
                14'h17a 	:	o_val <= 16'b0001001010000011;
                14'h17b 	:	o_val <= 16'b0001001010010000;
                14'h17c 	:	o_val <= 16'b0001001010011100;
                14'h17d 	:	o_val <= 16'b0001001010101000;
                14'h17e 	:	o_val <= 16'b0001001010110101;
                14'h17f 	:	o_val <= 16'b0001001011000001;
                14'h180 	:	o_val <= 16'b0001001011001110;
                14'h181 	:	o_val <= 16'b0001001011011010;
                14'h182 	:	o_val <= 16'b0001001011100111;
                14'h183 	:	o_val <= 16'b0001001011110011;
                14'h184 	:	o_val <= 16'b0001001011111111;
                14'h185 	:	o_val <= 16'b0001001100001100;
                14'h186 	:	o_val <= 16'b0001001100011000;
                14'h187 	:	o_val <= 16'b0001001100100101;
                14'h188 	:	o_val <= 16'b0001001100110001;
                14'h189 	:	o_val <= 16'b0001001100111110;
                14'h18a 	:	o_val <= 16'b0001001101001010;
                14'h18b 	:	o_val <= 16'b0001001101010110;
                14'h18c 	:	o_val <= 16'b0001001101100011;
                14'h18d 	:	o_val <= 16'b0001001101101111;
                14'h18e 	:	o_val <= 16'b0001001101111100;
                14'h18f 	:	o_val <= 16'b0001001110001000;
                14'h190 	:	o_val <= 16'b0001001110010101;
                14'h191 	:	o_val <= 16'b0001001110100001;
                14'h192 	:	o_val <= 16'b0001001110101101;
                14'h193 	:	o_val <= 16'b0001001110111010;
                14'h194 	:	o_val <= 16'b0001001111000110;
                14'h195 	:	o_val <= 16'b0001001111010011;
                14'h196 	:	o_val <= 16'b0001001111011111;
                14'h197 	:	o_val <= 16'b0001001111101011;
                14'h198 	:	o_val <= 16'b0001001111111000;
                14'h199 	:	o_val <= 16'b0001010000000100;
                14'h19a 	:	o_val <= 16'b0001010000010001;
                14'h19b 	:	o_val <= 16'b0001010000011101;
                14'h19c 	:	o_val <= 16'b0001010000101010;
                14'h19d 	:	o_val <= 16'b0001010000110110;
                14'h19e 	:	o_val <= 16'b0001010001000010;
                14'h19f 	:	o_val <= 16'b0001010001001111;
                14'h1a0 	:	o_val <= 16'b0001010001011011;
                14'h1a1 	:	o_val <= 16'b0001010001101000;
                14'h1a2 	:	o_val <= 16'b0001010001110100;
                14'h1a3 	:	o_val <= 16'b0001010010000000;
                14'h1a4 	:	o_val <= 16'b0001010010001101;
                14'h1a5 	:	o_val <= 16'b0001010010011001;
                14'h1a6 	:	o_val <= 16'b0001010010100110;
                14'h1a7 	:	o_val <= 16'b0001010010110010;
                14'h1a8 	:	o_val <= 16'b0001010010111110;
                14'h1a9 	:	o_val <= 16'b0001010011001011;
                14'h1aa 	:	o_val <= 16'b0001010011010111;
                14'h1ab 	:	o_val <= 16'b0001010011100100;
                14'h1ac 	:	o_val <= 16'b0001010011110000;
                14'h1ad 	:	o_val <= 16'b0001010011111100;
                14'h1ae 	:	o_val <= 16'b0001010100001001;
                14'h1af 	:	o_val <= 16'b0001010100010101;
                14'h1b0 	:	o_val <= 16'b0001010100100010;
                14'h1b1 	:	o_val <= 16'b0001010100101110;
                14'h1b2 	:	o_val <= 16'b0001010100111010;
                14'h1b3 	:	o_val <= 16'b0001010101000111;
                14'h1b4 	:	o_val <= 16'b0001010101010011;
                14'h1b5 	:	o_val <= 16'b0001010101100000;
                14'h1b6 	:	o_val <= 16'b0001010101101100;
                14'h1b7 	:	o_val <= 16'b0001010101111000;
                14'h1b8 	:	o_val <= 16'b0001010110000101;
                14'h1b9 	:	o_val <= 16'b0001010110010001;
                14'h1ba 	:	o_val <= 16'b0001010110011101;
                14'h1bb 	:	o_val <= 16'b0001010110101010;
                14'h1bc 	:	o_val <= 16'b0001010110110110;
                14'h1bd 	:	o_val <= 16'b0001010111000011;
                14'h1be 	:	o_val <= 16'b0001010111001111;
                14'h1bf 	:	o_val <= 16'b0001010111011011;
                14'h1c0 	:	o_val <= 16'b0001010111101000;
                14'h1c1 	:	o_val <= 16'b0001010111110100;
                14'h1c2 	:	o_val <= 16'b0001011000000001;
                14'h1c3 	:	o_val <= 16'b0001011000001101;
                14'h1c4 	:	o_val <= 16'b0001011000011001;
                14'h1c5 	:	o_val <= 16'b0001011000100110;
                14'h1c6 	:	o_val <= 16'b0001011000110010;
                14'h1c7 	:	o_val <= 16'b0001011000111110;
                14'h1c8 	:	o_val <= 16'b0001011001001011;
                14'h1c9 	:	o_val <= 16'b0001011001010111;
                14'h1ca 	:	o_val <= 16'b0001011001100100;
                14'h1cb 	:	o_val <= 16'b0001011001110000;
                14'h1cc 	:	o_val <= 16'b0001011001111100;
                14'h1cd 	:	o_val <= 16'b0001011010001001;
                14'h1ce 	:	o_val <= 16'b0001011010010101;
                14'h1cf 	:	o_val <= 16'b0001011010100001;
                14'h1d0 	:	o_val <= 16'b0001011010101110;
                14'h1d1 	:	o_val <= 16'b0001011010111010;
                14'h1d2 	:	o_val <= 16'b0001011011000110;
                14'h1d3 	:	o_val <= 16'b0001011011010011;
                14'h1d4 	:	o_val <= 16'b0001011011011111;
                14'h1d5 	:	o_val <= 16'b0001011011101100;
                14'h1d6 	:	o_val <= 16'b0001011011111000;
                14'h1d7 	:	o_val <= 16'b0001011100000100;
                14'h1d8 	:	o_val <= 16'b0001011100010001;
                14'h1d9 	:	o_val <= 16'b0001011100011101;
                14'h1da 	:	o_val <= 16'b0001011100101001;
                14'h1db 	:	o_val <= 16'b0001011100110110;
                14'h1dc 	:	o_val <= 16'b0001011101000010;
                14'h1dd 	:	o_val <= 16'b0001011101001110;
                14'h1de 	:	o_val <= 16'b0001011101011011;
                14'h1df 	:	o_val <= 16'b0001011101100111;
                14'h1e0 	:	o_val <= 16'b0001011101110100;
                14'h1e1 	:	o_val <= 16'b0001011110000000;
                14'h1e2 	:	o_val <= 16'b0001011110001100;
                14'h1e3 	:	o_val <= 16'b0001011110011001;
                14'h1e4 	:	o_val <= 16'b0001011110100101;
                14'h1e5 	:	o_val <= 16'b0001011110110001;
                14'h1e6 	:	o_val <= 16'b0001011110111110;
                14'h1e7 	:	o_val <= 16'b0001011111001010;
                14'h1e8 	:	o_val <= 16'b0001011111010110;
                14'h1e9 	:	o_val <= 16'b0001011111100011;
                14'h1ea 	:	o_val <= 16'b0001011111101111;
                14'h1eb 	:	o_val <= 16'b0001011111111011;
                14'h1ec 	:	o_val <= 16'b0001100000001000;
                14'h1ed 	:	o_val <= 16'b0001100000010100;
                14'h1ee 	:	o_val <= 16'b0001100000100000;
                14'h1ef 	:	o_val <= 16'b0001100000101101;
                14'h1f0 	:	o_val <= 16'b0001100000111001;
                14'h1f1 	:	o_val <= 16'b0001100001000101;
                14'h1f2 	:	o_val <= 16'b0001100001010010;
                14'h1f3 	:	o_val <= 16'b0001100001011110;
                14'h1f4 	:	o_val <= 16'b0001100001101010;
                14'h1f5 	:	o_val <= 16'b0001100001110111;
                14'h1f6 	:	o_val <= 16'b0001100010000011;
                14'h1f7 	:	o_val <= 16'b0001100010001111;
                14'h1f8 	:	o_val <= 16'b0001100010011100;
                14'h1f9 	:	o_val <= 16'b0001100010101000;
                14'h1fa 	:	o_val <= 16'b0001100010110100;
                14'h1fb 	:	o_val <= 16'b0001100011000001;
                14'h1fc 	:	o_val <= 16'b0001100011001101;
                14'h1fd 	:	o_val <= 16'b0001100011011001;
                14'h1fe 	:	o_val <= 16'b0001100011100110;
                14'h1ff 	:	o_val <= 16'b0001100011110010;
                14'h200 	:	o_val <= 16'b0001100011111110;
                14'h201 	:	o_val <= 16'b0001100100001011;
                14'h202 	:	o_val <= 16'b0001100100010111;
                14'h203 	:	o_val <= 16'b0001100100100011;
                14'h204 	:	o_val <= 16'b0001100100110000;
                14'h205 	:	o_val <= 16'b0001100100111100;
                14'h206 	:	o_val <= 16'b0001100101001000;
                14'h207 	:	o_val <= 16'b0001100101010101;
                14'h208 	:	o_val <= 16'b0001100101100001;
                14'h209 	:	o_val <= 16'b0001100101101101;
                14'h20a 	:	o_val <= 16'b0001100101111010;
                14'h20b 	:	o_val <= 16'b0001100110000110;
                14'h20c 	:	o_val <= 16'b0001100110010010;
                14'h20d 	:	o_val <= 16'b0001100110011111;
                14'h20e 	:	o_val <= 16'b0001100110101011;
                14'h20f 	:	o_val <= 16'b0001100110110111;
                14'h210 	:	o_val <= 16'b0001100111000011;
                14'h211 	:	o_val <= 16'b0001100111010000;
                14'h212 	:	o_val <= 16'b0001100111011100;
                14'h213 	:	o_val <= 16'b0001100111101000;
                14'h214 	:	o_val <= 16'b0001100111110101;
                14'h215 	:	o_val <= 16'b0001101000000001;
                14'h216 	:	o_val <= 16'b0001101000001101;
                14'h217 	:	o_val <= 16'b0001101000011010;
                14'h218 	:	o_val <= 16'b0001101000100110;
                14'h219 	:	o_val <= 16'b0001101000110010;
                14'h21a 	:	o_val <= 16'b0001101000111110;
                14'h21b 	:	o_val <= 16'b0001101001001011;
                14'h21c 	:	o_val <= 16'b0001101001010111;
                14'h21d 	:	o_val <= 16'b0001101001100011;
                14'h21e 	:	o_val <= 16'b0001101001110000;
                14'h21f 	:	o_val <= 16'b0001101001111100;
                14'h220 	:	o_val <= 16'b0001101010001000;
                14'h221 	:	o_val <= 16'b0001101010010101;
                14'h222 	:	o_val <= 16'b0001101010100001;
                14'h223 	:	o_val <= 16'b0001101010101101;
                14'h224 	:	o_val <= 16'b0001101010111001;
                14'h225 	:	o_val <= 16'b0001101011000110;
                14'h226 	:	o_val <= 16'b0001101011010010;
                14'h227 	:	o_val <= 16'b0001101011011110;
                14'h228 	:	o_val <= 16'b0001101011101011;
                14'h229 	:	o_val <= 16'b0001101011110111;
                14'h22a 	:	o_val <= 16'b0001101100000011;
                14'h22b 	:	o_val <= 16'b0001101100001111;
                14'h22c 	:	o_val <= 16'b0001101100011100;
                14'h22d 	:	o_val <= 16'b0001101100101000;
                14'h22e 	:	o_val <= 16'b0001101100110100;
                14'h22f 	:	o_val <= 16'b0001101101000001;
                14'h230 	:	o_val <= 16'b0001101101001101;
                14'h231 	:	o_val <= 16'b0001101101011001;
                14'h232 	:	o_val <= 16'b0001101101100101;
                14'h233 	:	o_val <= 16'b0001101101110010;
                14'h234 	:	o_val <= 16'b0001101101111110;
                14'h235 	:	o_val <= 16'b0001101110001010;
                14'h236 	:	o_val <= 16'b0001101110010110;
                14'h237 	:	o_val <= 16'b0001101110100011;
                14'h238 	:	o_val <= 16'b0001101110101111;
                14'h239 	:	o_val <= 16'b0001101110111011;
                14'h23a 	:	o_val <= 16'b0001101111001000;
                14'h23b 	:	o_val <= 16'b0001101111010100;
                14'h23c 	:	o_val <= 16'b0001101111100000;
                14'h23d 	:	o_val <= 16'b0001101111101100;
                14'h23e 	:	o_val <= 16'b0001101111111001;
                14'h23f 	:	o_val <= 16'b0001110000000101;
                14'h240 	:	o_val <= 16'b0001110000010001;
                14'h241 	:	o_val <= 16'b0001110000011101;
                14'h242 	:	o_val <= 16'b0001110000101010;
                14'h243 	:	o_val <= 16'b0001110000110110;
                14'h244 	:	o_val <= 16'b0001110001000010;
                14'h245 	:	o_val <= 16'b0001110001001110;
                14'h246 	:	o_val <= 16'b0001110001011011;
                14'h247 	:	o_val <= 16'b0001110001100111;
                14'h248 	:	o_val <= 16'b0001110001110011;
                14'h249 	:	o_val <= 16'b0001110001111111;
                14'h24a 	:	o_val <= 16'b0001110010001100;
                14'h24b 	:	o_val <= 16'b0001110010011000;
                14'h24c 	:	o_val <= 16'b0001110010100100;
                14'h24d 	:	o_val <= 16'b0001110010110000;
                14'h24e 	:	o_val <= 16'b0001110010111101;
                14'h24f 	:	o_val <= 16'b0001110011001001;
                14'h250 	:	o_val <= 16'b0001110011010101;
                14'h251 	:	o_val <= 16'b0001110011100001;
                14'h252 	:	o_val <= 16'b0001110011101110;
                14'h253 	:	o_val <= 16'b0001110011111010;
                14'h254 	:	o_val <= 16'b0001110100000110;
                14'h255 	:	o_val <= 16'b0001110100010010;
                14'h256 	:	o_val <= 16'b0001110100011111;
                14'h257 	:	o_val <= 16'b0001110100101011;
                14'h258 	:	o_val <= 16'b0001110100110111;
                14'h259 	:	o_val <= 16'b0001110101000011;
                14'h25a 	:	o_val <= 16'b0001110101010000;
                14'h25b 	:	o_val <= 16'b0001110101011100;
                14'h25c 	:	o_val <= 16'b0001110101101000;
                14'h25d 	:	o_val <= 16'b0001110101110100;
                14'h25e 	:	o_val <= 16'b0001110110000000;
                14'h25f 	:	o_val <= 16'b0001110110001101;
                14'h260 	:	o_val <= 16'b0001110110011001;
                14'h261 	:	o_val <= 16'b0001110110100101;
                14'h262 	:	o_val <= 16'b0001110110110001;
                14'h263 	:	o_val <= 16'b0001110110111110;
                14'h264 	:	o_val <= 16'b0001110111001010;
                14'h265 	:	o_val <= 16'b0001110111010110;
                14'h266 	:	o_val <= 16'b0001110111100010;
                14'h267 	:	o_val <= 16'b0001110111101110;
                14'h268 	:	o_val <= 16'b0001110111111011;
                14'h269 	:	o_val <= 16'b0001111000000111;
                14'h26a 	:	o_val <= 16'b0001111000010011;
                14'h26b 	:	o_val <= 16'b0001111000011111;
                14'h26c 	:	o_val <= 16'b0001111000101100;
                14'h26d 	:	o_val <= 16'b0001111000111000;
                14'h26e 	:	o_val <= 16'b0001111001000100;
                14'h26f 	:	o_val <= 16'b0001111001010000;
                14'h270 	:	o_val <= 16'b0001111001011100;
                14'h271 	:	o_val <= 16'b0001111001101001;
                14'h272 	:	o_val <= 16'b0001111001110101;
                14'h273 	:	o_val <= 16'b0001111010000001;
                14'h274 	:	o_val <= 16'b0001111010001101;
                14'h275 	:	o_val <= 16'b0001111010011001;
                14'h276 	:	o_val <= 16'b0001111010100110;
                14'h277 	:	o_val <= 16'b0001111010110010;
                14'h278 	:	o_val <= 16'b0001111010111110;
                14'h279 	:	o_val <= 16'b0001111011001010;
                14'h27a 	:	o_val <= 16'b0001111011010110;
                14'h27b 	:	o_val <= 16'b0001111011100011;
                14'h27c 	:	o_val <= 16'b0001111011101111;
                14'h27d 	:	o_val <= 16'b0001111011111011;
                14'h27e 	:	o_val <= 16'b0001111100000111;
                14'h27f 	:	o_val <= 16'b0001111100010011;
                14'h280 	:	o_val <= 16'b0001111100100000;
                14'h281 	:	o_val <= 16'b0001111100101100;
                14'h282 	:	o_val <= 16'b0001111100111000;
                14'h283 	:	o_val <= 16'b0001111101000100;
                14'h284 	:	o_val <= 16'b0001111101010000;
                14'h285 	:	o_val <= 16'b0001111101011101;
                14'h286 	:	o_val <= 16'b0001111101101001;
                14'h287 	:	o_val <= 16'b0001111101110101;
                14'h288 	:	o_val <= 16'b0001111110000001;
                14'h289 	:	o_val <= 16'b0001111110001101;
                14'h28a 	:	o_val <= 16'b0001111110011001;
                14'h28b 	:	o_val <= 16'b0001111110100110;
                14'h28c 	:	o_val <= 16'b0001111110110010;
                14'h28d 	:	o_val <= 16'b0001111110111110;
                14'h28e 	:	o_val <= 16'b0001111111001010;
                14'h28f 	:	o_val <= 16'b0001111111010110;
                14'h290 	:	o_val <= 16'b0001111111100010;
                14'h291 	:	o_val <= 16'b0001111111101111;
                14'h292 	:	o_val <= 16'b0001111111111011;
                14'h293 	:	o_val <= 16'b0010000000000111;
                14'h294 	:	o_val <= 16'b0010000000010011;
                14'h295 	:	o_val <= 16'b0010000000011111;
                14'h296 	:	o_val <= 16'b0010000000101011;
                14'h297 	:	o_val <= 16'b0010000000111000;
                14'h298 	:	o_val <= 16'b0010000001000100;
                14'h299 	:	o_val <= 16'b0010000001010000;
                14'h29a 	:	o_val <= 16'b0010000001011100;
                14'h29b 	:	o_val <= 16'b0010000001101000;
                14'h29c 	:	o_val <= 16'b0010000001110100;
                14'h29d 	:	o_val <= 16'b0010000010000001;
                14'h29e 	:	o_val <= 16'b0010000010001101;
                14'h29f 	:	o_val <= 16'b0010000010011001;
                14'h2a0 	:	o_val <= 16'b0010000010100101;
                14'h2a1 	:	o_val <= 16'b0010000010110001;
                14'h2a2 	:	o_val <= 16'b0010000010111101;
                14'h2a3 	:	o_val <= 16'b0010000011001001;
                14'h2a4 	:	o_val <= 16'b0010000011010110;
                14'h2a5 	:	o_val <= 16'b0010000011100010;
                14'h2a6 	:	o_val <= 16'b0010000011101110;
                14'h2a7 	:	o_val <= 16'b0010000011111010;
                14'h2a8 	:	o_val <= 16'b0010000100000110;
                14'h2a9 	:	o_val <= 16'b0010000100010010;
                14'h2aa 	:	o_val <= 16'b0010000100011110;
                14'h2ab 	:	o_val <= 16'b0010000100101011;
                14'h2ac 	:	o_val <= 16'b0010000100110111;
                14'h2ad 	:	o_val <= 16'b0010000101000011;
                14'h2ae 	:	o_val <= 16'b0010000101001111;
                14'h2af 	:	o_val <= 16'b0010000101011011;
                14'h2b0 	:	o_val <= 16'b0010000101100111;
                14'h2b1 	:	o_val <= 16'b0010000101110011;
                14'h2b2 	:	o_val <= 16'b0010000110000000;
                14'h2b3 	:	o_val <= 16'b0010000110001100;
                14'h2b4 	:	o_val <= 16'b0010000110011000;
                14'h2b5 	:	o_val <= 16'b0010000110100100;
                14'h2b6 	:	o_val <= 16'b0010000110110000;
                14'h2b7 	:	o_val <= 16'b0010000110111100;
                14'h2b8 	:	o_val <= 16'b0010000111001000;
                14'h2b9 	:	o_val <= 16'b0010000111010100;
                14'h2ba 	:	o_val <= 16'b0010000111100001;
                14'h2bb 	:	o_val <= 16'b0010000111101101;
                14'h2bc 	:	o_val <= 16'b0010000111111001;
                14'h2bd 	:	o_val <= 16'b0010001000000101;
                14'h2be 	:	o_val <= 16'b0010001000010001;
                14'h2bf 	:	o_val <= 16'b0010001000011101;
                14'h2c0 	:	o_val <= 16'b0010001000101001;
                14'h2c1 	:	o_val <= 16'b0010001000110101;
                14'h2c2 	:	o_val <= 16'b0010001001000001;
                14'h2c3 	:	o_val <= 16'b0010001001001110;
                14'h2c4 	:	o_val <= 16'b0010001001011010;
                14'h2c5 	:	o_val <= 16'b0010001001100110;
                14'h2c6 	:	o_val <= 16'b0010001001110010;
                14'h2c7 	:	o_val <= 16'b0010001001111110;
                14'h2c8 	:	o_val <= 16'b0010001010001010;
                14'h2c9 	:	o_val <= 16'b0010001010010110;
                14'h2ca 	:	o_val <= 16'b0010001010100010;
                14'h2cb 	:	o_val <= 16'b0010001010101110;
                14'h2cc 	:	o_val <= 16'b0010001010111010;
                14'h2cd 	:	o_val <= 16'b0010001011000111;
                14'h2ce 	:	o_val <= 16'b0010001011010011;
                14'h2cf 	:	o_val <= 16'b0010001011011111;
                14'h2d0 	:	o_val <= 16'b0010001011101011;
                14'h2d1 	:	o_val <= 16'b0010001011110111;
                14'h2d2 	:	o_val <= 16'b0010001100000011;
                14'h2d3 	:	o_val <= 16'b0010001100001111;
                14'h2d4 	:	o_val <= 16'b0010001100011011;
                14'h2d5 	:	o_val <= 16'b0010001100100111;
                14'h2d6 	:	o_val <= 16'b0010001100110011;
                14'h2d7 	:	o_val <= 16'b0010001100111111;
                14'h2d8 	:	o_val <= 16'b0010001101001011;
                14'h2d9 	:	o_val <= 16'b0010001101011000;
                14'h2da 	:	o_val <= 16'b0010001101100100;
                14'h2db 	:	o_val <= 16'b0010001101110000;
                14'h2dc 	:	o_val <= 16'b0010001101111100;
                14'h2dd 	:	o_val <= 16'b0010001110001000;
                14'h2de 	:	o_val <= 16'b0010001110010100;
                14'h2df 	:	o_val <= 16'b0010001110100000;
                14'h2e0 	:	o_val <= 16'b0010001110101100;
                14'h2e1 	:	o_val <= 16'b0010001110111000;
                14'h2e2 	:	o_val <= 16'b0010001111000100;
                14'h2e3 	:	o_val <= 16'b0010001111010000;
                14'h2e4 	:	o_val <= 16'b0010001111011100;
                14'h2e5 	:	o_val <= 16'b0010001111101000;
                14'h2e6 	:	o_val <= 16'b0010001111110100;
                14'h2e7 	:	o_val <= 16'b0010010000000001;
                14'h2e8 	:	o_val <= 16'b0010010000001101;
                14'h2e9 	:	o_val <= 16'b0010010000011001;
                14'h2ea 	:	o_val <= 16'b0010010000100101;
                14'h2eb 	:	o_val <= 16'b0010010000110001;
                14'h2ec 	:	o_val <= 16'b0010010000111101;
                14'h2ed 	:	o_val <= 16'b0010010001001001;
                14'h2ee 	:	o_val <= 16'b0010010001010101;
                14'h2ef 	:	o_val <= 16'b0010010001100001;
                14'h2f0 	:	o_val <= 16'b0010010001101101;
                14'h2f1 	:	o_val <= 16'b0010010001111001;
                14'h2f2 	:	o_val <= 16'b0010010010000101;
                14'h2f3 	:	o_val <= 16'b0010010010010001;
                14'h2f4 	:	o_val <= 16'b0010010010011101;
                14'h2f5 	:	o_val <= 16'b0010010010101001;
                14'h2f6 	:	o_val <= 16'b0010010010110101;
                14'h2f7 	:	o_val <= 16'b0010010011000001;
                14'h2f8 	:	o_val <= 16'b0010010011001101;
                14'h2f9 	:	o_val <= 16'b0010010011011001;
                14'h2fa 	:	o_val <= 16'b0010010011100101;
                14'h2fb 	:	o_val <= 16'b0010010011110001;
                14'h2fc 	:	o_val <= 16'b0010010011111101;
                14'h2fd 	:	o_val <= 16'b0010010100001001;
                14'h2fe 	:	o_val <= 16'b0010010100010110;
                14'h2ff 	:	o_val <= 16'b0010010100100010;
                14'h300 	:	o_val <= 16'b0010010100101110;
                14'h301 	:	o_val <= 16'b0010010100111010;
                14'h302 	:	o_val <= 16'b0010010101000110;
                14'h303 	:	o_val <= 16'b0010010101010010;
                14'h304 	:	o_val <= 16'b0010010101011110;
                14'h305 	:	o_val <= 16'b0010010101101010;
                14'h306 	:	o_val <= 16'b0010010101110110;
                14'h307 	:	o_val <= 16'b0010010110000010;
                14'h308 	:	o_val <= 16'b0010010110001110;
                14'h309 	:	o_val <= 16'b0010010110011010;
                14'h30a 	:	o_val <= 16'b0010010110100110;
                14'h30b 	:	o_val <= 16'b0010010110110010;
                14'h30c 	:	o_val <= 16'b0010010110111110;
                14'h30d 	:	o_val <= 16'b0010010111001010;
                14'h30e 	:	o_val <= 16'b0010010111010110;
                14'h30f 	:	o_val <= 16'b0010010111100010;
                14'h310 	:	o_val <= 16'b0010010111101110;
                14'h311 	:	o_val <= 16'b0010010111111010;
                14'h312 	:	o_val <= 16'b0010011000000110;
                14'h313 	:	o_val <= 16'b0010011000010010;
                14'h314 	:	o_val <= 16'b0010011000011110;
                14'h315 	:	o_val <= 16'b0010011000101010;
                14'h316 	:	o_val <= 16'b0010011000110110;
                14'h317 	:	o_val <= 16'b0010011001000010;
                14'h318 	:	o_val <= 16'b0010011001001110;
                14'h319 	:	o_val <= 16'b0010011001011010;
                14'h31a 	:	o_val <= 16'b0010011001100110;
                14'h31b 	:	o_val <= 16'b0010011001110010;
                14'h31c 	:	o_val <= 16'b0010011001111110;
                14'h31d 	:	o_val <= 16'b0010011010001010;
                14'h31e 	:	o_val <= 16'b0010011010010110;
                14'h31f 	:	o_val <= 16'b0010011010100010;
                14'h320 	:	o_val <= 16'b0010011010101110;
                14'h321 	:	o_val <= 16'b0010011010111010;
                14'h322 	:	o_val <= 16'b0010011011000110;
                14'h323 	:	o_val <= 16'b0010011011010010;
                14'h324 	:	o_val <= 16'b0010011011011110;
                14'h325 	:	o_val <= 16'b0010011011101001;
                14'h326 	:	o_val <= 16'b0010011011110101;
                14'h327 	:	o_val <= 16'b0010011100000001;
                14'h328 	:	o_val <= 16'b0010011100001101;
                14'h329 	:	o_val <= 16'b0010011100011001;
                14'h32a 	:	o_val <= 16'b0010011100100101;
                14'h32b 	:	o_val <= 16'b0010011100110001;
                14'h32c 	:	o_val <= 16'b0010011100111101;
                14'h32d 	:	o_val <= 16'b0010011101001001;
                14'h32e 	:	o_val <= 16'b0010011101010101;
                14'h32f 	:	o_val <= 16'b0010011101100001;
                14'h330 	:	o_val <= 16'b0010011101101101;
                14'h331 	:	o_val <= 16'b0010011101111001;
                14'h332 	:	o_val <= 16'b0010011110000101;
                14'h333 	:	o_val <= 16'b0010011110010001;
                14'h334 	:	o_val <= 16'b0010011110011101;
                14'h335 	:	o_val <= 16'b0010011110101001;
                14'h336 	:	o_val <= 16'b0010011110110101;
                14'h337 	:	o_val <= 16'b0010011111000001;
                14'h338 	:	o_val <= 16'b0010011111001101;
                14'h339 	:	o_val <= 16'b0010011111011001;
                14'h33a 	:	o_val <= 16'b0010011111100101;
                14'h33b 	:	o_val <= 16'b0010011111110001;
                14'h33c 	:	o_val <= 16'b0010011111111100;
                14'h33d 	:	o_val <= 16'b0010100000001000;
                14'h33e 	:	o_val <= 16'b0010100000010100;
                14'h33f 	:	o_val <= 16'b0010100000100000;
                14'h340 	:	o_val <= 16'b0010100000101100;
                14'h341 	:	o_val <= 16'b0010100000111000;
                14'h342 	:	o_val <= 16'b0010100001000100;
                14'h343 	:	o_val <= 16'b0010100001010000;
                14'h344 	:	o_val <= 16'b0010100001011100;
                14'h345 	:	o_val <= 16'b0010100001101000;
                14'h346 	:	o_val <= 16'b0010100001110100;
                14'h347 	:	o_val <= 16'b0010100010000000;
                14'h348 	:	o_val <= 16'b0010100010001100;
                14'h349 	:	o_val <= 16'b0010100010011000;
                14'h34a 	:	o_val <= 16'b0010100010100011;
                14'h34b 	:	o_val <= 16'b0010100010101111;
                14'h34c 	:	o_val <= 16'b0010100010111011;
                14'h34d 	:	o_val <= 16'b0010100011000111;
                14'h34e 	:	o_val <= 16'b0010100011010011;
                14'h34f 	:	o_val <= 16'b0010100011011111;
                14'h350 	:	o_val <= 16'b0010100011101011;
                14'h351 	:	o_val <= 16'b0010100011110111;
                14'h352 	:	o_val <= 16'b0010100100000011;
                14'h353 	:	o_val <= 16'b0010100100001111;
                14'h354 	:	o_val <= 16'b0010100100011011;
                14'h355 	:	o_val <= 16'b0010100100100110;
                14'h356 	:	o_val <= 16'b0010100100110010;
                14'h357 	:	o_val <= 16'b0010100100111110;
                14'h358 	:	o_val <= 16'b0010100101001010;
                14'h359 	:	o_val <= 16'b0010100101010110;
                14'h35a 	:	o_val <= 16'b0010100101100010;
                14'h35b 	:	o_val <= 16'b0010100101101110;
                14'h35c 	:	o_val <= 16'b0010100101111010;
                14'h35d 	:	o_val <= 16'b0010100110000110;
                14'h35e 	:	o_val <= 16'b0010100110010001;
                14'h35f 	:	o_val <= 16'b0010100110011101;
                14'h360 	:	o_val <= 16'b0010100110101001;
                14'h361 	:	o_val <= 16'b0010100110110101;
                14'h362 	:	o_val <= 16'b0010100111000001;
                14'h363 	:	o_val <= 16'b0010100111001101;
                14'h364 	:	o_val <= 16'b0010100111011001;
                14'h365 	:	o_val <= 16'b0010100111100101;
                14'h366 	:	o_val <= 16'b0010100111110000;
                14'h367 	:	o_val <= 16'b0010100111111100;
                14'h368 	:	o_val <= 16'b0010101000001000;
                14'h369 	:	o_val <= 16'b0010101000010100;
                14'h36a 	:	o_val <= 16'b0010101000100000;
                14'h36b 	:	o_val <= 16'b0010101000101100;
                14'h36c 	:	o_val <= 16'b0010101000111000;
                14'h36d 	:	o_val <= 16'b0010101001000100;
                14'h36e 	:	o_val <= 16'b0010101001001111;
                14'h36f 	:	o_val <= 16'b0010101001011011;
                14'h370 	:	o_val <= 16'b0010101001100111;
                14'h371 	:	o_val <= 16'b0010101001110011;
                14'h372 	:	o_val <= 16'b0010101001111111;
                14'h373 	:	o_val <= 16'b0010101010001011;
                14'h374 	:	o_val <= 16'b0010101010010111;
                14'h375 	:	o_val <= 16'b0010101010100010;
                14'h376 	:	o_val <= 16'b0010101010101110;
                14'h377 	:	o_val <= 16'b0010101010111010;
                14'h378 	:	o_val <= 16'b0010101011000110;
                14'h379 	:	o_val <= 16'b0010101011010010;
                14'h37a 	:	o_val <= 16'b0010101011011110;
                14'h37b 	:	o_val <= 16'b0010101011101001;
                14'h37c 	:	o_val <= 16'b0010101011110101;
                14'h37d 	:	o_val <= 16'b0010101100000001;
                14'h37e 	:	o_val <= 16'b0010101100001101;
                14'h37f 	:	o_val <= 16'b0010101100011001;
                14'h380 	:	o_val <= 16'b0010101100100101;
                14'h381 	:	o_val <= 16'b0010101100110000;
                14'h382 	:	o_val <= 16'b0010101100111100;
                14'h383 	:	o_val <= 16'b0010101101001000;
                14'h384 	:	o_val <= 16'b0010101101010100;
                14'h385 	:	o_val <= 16'b0010101101100000;
                14'h386 	:	o_val <= 16'b0010101101101100;
                14'h387 	:	o_val <= 16'b0010101101110111;
                14'h388 	:	o_val <= 16'b0010101110000011;
                14'h389 	:	o_val <= 16'b0010101110001111;
                14'h38a 	:	o_val <= 16'b0010101110011011;
                14'h38b 	:	o_val <= 16'b0010101110100111;
                14'h38c 	:	o_val <= 16'b0010101110110010;
                14'h38d 	:	o_val <= 16'b0010101110111110;
                14'h38e 	:	o_val <= 16'b0010101111001010;
                14'h38f 	:	o_val <= 16'b0010101111010110;
                14'h390 	:	o_val <= 16'b0010101111100010;
                14'h391 	:	o_val <= 16'b0010101111101110;
                14'h392 	:	o_val <= 16'b0010101111111001;
                14'h393 	:	o_val <= 16'b0010110000000101;
                14'h394 	:	o_val <= 16'b0010110000010001;
                14'h395 	:	o_val <= 16'b0010110000011101;
                14'h396 	:	o_val <= 16'b0010110000101001;
                14'h397 	:	o_val <= 16'b0010110000110100;
                14'h398 	:	o_val <= 16'b0010110001000000;
                14'h399 	:	o_val <= 16'b0010110001001100;
                14'h39a 	:	o_val <= 16'b0010110001011000;
                14'h39b 	:	o_val <= 16'b0010110001100011;
                14'h39c 	:	o_val <= 16'b0010110001101111;
                14'h39d 	:	o_val <= 16'b0010110001111011;
                14'h39e 	:	o_val <= 16'b0010110010000111;
                14'h39f 	:	o_val <= 16'b0010110010010011;
                14'h3a0 	:	o_val <= 16'b0010110010011110;
                14'h3a1 	:	o_val <= 16'b0010110010101010;
                14'h3a2 	:	o_val <= 16'b0010110010110110;
                14'h3a3 	:	o_val <= 16'b0010110011000010;
                14'h3a4 	:	o_val <= 16'b0010110011001101;
                14'h3a5 	:	o_val <= 16'b0010110011011001;
                14'h3a6 	:	o_val <= 16'b0010110011100101;
                14'h3a7 	:	o_val <= 16'b0010110011110001;
                14'h3a8 	:	o_val <= 16'b0010110011111101;
                14'h3a9 	:	o_val <= 16'b0010110100001000;
                14'h3aa 	:	o_val <= 16'b0010110100010100;
                14'h3ab 	:	o_val <= 16'b0010110100100000;
                14'h3ac 	:	o_val <= 16'b0010110100101100;
                14'h3ad 	:	o_val <= 16'b0010110100110111;
                14'h3ae 	:	o_val <= 16'b0010110101000011;
                14'h3af 	:	o_val <= 16'b0010110101001111;
                14'h3b0 	:	o_val <= 16'b0010110101011011;
                14'h3b1 	:	o_val <= 16'b0010110101100110;
                14'h3b2 	:	o_val <= 16'b0010110101110010;
                14'h3b3 	:	o_val <= 16'b0010110101111110;
                14'h3b4 	:	o_val <= 16'b0010110110001010;
                14'h3b5 	:	o_val <= 16'b0010110110010101;
                14'h3b6 	:	o_val <= 16'b0010110110100001;
                14'h3b7 	:	o_val <= 16'b0010110110101101;
                14'h3b8 	:	o_val <= 16'b0010110110111001;
                14'h3b9 	:	o_val <= 16'b0010110111000100;
                14'h3ba 	:	o_val <= 16'b0010110111010000;
                14'h3bb 	:	o_val <= 16'b0010110111011100;
                14'h3bc 	:	o_val <= 16'b0010110111100111;
                14'h3bd 	:	o_val <= 16'b0010110111110011;
                14'h3be 	:	o_val <= 16'b0010110111111111;
                14'h3bf 	:	o_val <= 16'b0010111000001011;
                14'h3c0 	:	o_val <= 16'b0010111000010110;
                14'h3c1 	:	o_val <= 16'b0010111000100010;
                14'h3c2 	:	o_val <= 16'b0010111000101110;
                14'h3c3 	:	o_val <= 16'b0010111000111010;
                14'h3c4 	:	o_val <= 16'b0010111001000101;
                14'h3c5 	:	o_val <= 16'b0010111001010001;
                14'h3c6 	:	o_val <= 16'b0010111001011101;
                14'h3c7 	:	o_val <= 16'b0010111001101000;
                14'h3c8 	:	o_val <= 16'b0010111001110100;
                14'h3c9 	:	o_val <= 16'b0010111010000000;
                14'h3ca 	:	o_val <= 16'b0010111010001100;
                14'h3cb 	:	o_val <= 16'b0010111010010111;
                14'h3cc 	:	o_val <= 16'b0010111010100011;
                14'h3cd 	:	o_val <= 16'b0010111010101111;
                14'h3ce 	:	o_val <= 16'b0010111010111010;
                14'h3cf 	:	o_val <= 16'b0010111011000110;
                14'h3d0 	:	o_val <= 16'b0010111011010010;
                14'h3d1 	:	o_val <= 16'b0010111011011101;
                14'h3d2 	:	o_val <= 16'b0010111011101001;
                14'h3d3 	:	o_val <= 16'b0010111011110101;
                14'h3d4 	:	o_val <= 16'b0010111100000001;
                14'h3d5 	:	o_val <= 16'b0010111100001100;
                14'h3d6 	:	o_val <= 16'b0010111100011000;
                14'h3d7 	:	o_val <= 16'b0010111100100100;
                14'h3d8 	:	o_val <= 16'b0010111100101111;
                14'h3d9 	:	o_val <= 16'b0010111100111011;
                14'h3da 	:	o_val <= 16'b0010111101000111;
                14'h3db 	:	o_val <= 16'b0010111101010010;
                14'h3dc 	:	o_val <= 16'b0010111101011110;
                14'h3dd 	:	o_val <= 16'b0010111101101010;
                14'h3de 	:	o_val <= 16'b0010111101110101;
                14'h3df 	:	o_val <= 16'b0010111110000001;
                14'h3e0 	:	o_val <= 16'b0010111110001101;
                14'h3e1 	:	o_val <= 16'b0010111110011000;
                14'h3e2 	:	o_val <= 16'b0010111110100100;
                14'h3e3 	:	o_val <= 16'b0010111110110000;
                14'h3e4 	:	o_val <= 16'b0010111110111011;
                14'h3e5 	:	o_val <= 16'b0010111111000111;
                14'h3e6 	:	o_val <= 16'b0010111111010011;
                14'h3e7 	:	o_val <= 16'b0010111111011110;
                14'h3e8 	:	o_val <= 16'b0010111111101010;
                14'h3e9 	:	o_val <= 16'b0010111111110110;
                14'h3ea 	:	o_val <= 16'b0011000000000001;
                14'h3eb 	:	o_val <= 16'b0011000000001101;
                14'h3ec 	:	o_val <= 16'b0011000000011001;
                14'h3ed 	:	o_val <= 16'b0011000000100100;
                14'h3ee 	:	o_val <= 16'b0011000000110000;
                14'h3ef 	:	o_val <= 16'b0011000000111011;
                14'h3f0 	:	o_val <= 16'b0011000001000111;
                14'h3f1 	:	o_val <= 16'b0011000001010011;
                14'h3f2 	:	o_val <= 16'b0011000001011110;
                14'h3f3 	:	o_val <= 16'b0011000001101010;
                14'h3f4 	:	o_val <= 16'b0011000001110110;
                14'h3f5 	:	o_val <= 16'b0011000010000001;
                14'h3f6 	:	o_val <= 16'b0011000010001101;
                14'h3f7 	:	o_val <= 16'b0011000010011001;
                14'h3f8 	:	o_val <= 16'b0011000010100100;
                14'h3f9 	:	o_val <= 16'b0011000010110000;
                14'h3fa 	:	o_val <= 16'b0011000010111011;
                14'h3fb 	:	o_val <= 16'b0011000011000111;
                14'h3fc 	:	o_val <= 16'b0011000011010011;
                14'h3fd 	:	o_val <= 16'b0011000011011110;
                14'h3fe 	:	o_val <= 16'b0011000011101010;
                14'h3ff 	:	o_val <= 16'b0011000011110101;
                14'h400 	:	o_val <= 16'b0011000100000001;
                14'h401 	:	o_val <= 16'b0011000100001101;
                14'h402 	:	o_val <= 16'b0011000100011000;
                14'h403 	:	o_val <= 16'b0011000100100100;
                14'h404 	:	o_val <= 16'b0011000100101111;
                14'h405 	:	o_val <= 16'b0011000100111011;
                14'h406 	:	o_val <= 16'b0011000101000111;
                14'h407 	:	o_val <= 16'b0011000101010010;
                14'h408 	:	o_val <= 16'b0011000101011110;
                14'h409 	:	o_val <= 16'b0011000101101001;
                14'h40a 	:	o_val <= 16'b0011000101110101;
                14'h40b 	:	o_val <= 16'b0011000110000001;
                14'h40c 	:	o_val <= 16'b0011000110001100;
                14'h40d 	:	o_val <= 16'b0011000110011000;
                14'h40e 	:	o_val <= 16'b0011000110100011;
                14'h40f 	:	o_val <= 16'b0011000110101111;
                14'h410 	:	o_val <= 16'b0011000110111011;
                14'h411 	:	o_val <= 16'b0011000111000110;
                14'h412 	:	o_val <= 16'b0011000111010010;
                14'h413 	:	o_val <= 16'b0011000111011101;
                14'h414 	:	o_val <= 16'b0011000111101001;
                14'h415 	:	o_val <= 16'b0011000111110100;
                14'h416 	:	o_val <= 16'b0011001000000000;
                14'h417 	:	o_val <= 16'b0011001000001100;
                14'h418 	:	o_val <= 16'b0011001000010111;
                14'h419 	:	o_val <= 16'b0011001000100011;
                14'h41a 	:	o_val <= 16'b0011001000101110;
                14'h41b 	:	o_val <= 16'b0011001000111010;
                14'h41c 	:	o_val <= 16'b0011001001000101;
                14'h41d 	:	o_val <= 16'b0011001001010001;
                14'h41e 	:	o_val <= 16'b0011001001011101;
                14'h41f 	:	o_val <= 16'b0011001001101000;
                14'h420 	:	o_val <= 16'b0011001001110100;
                14'h421 	:	o_val <= 16'b0011001001111111;
                14'h422 	:	o_val <= 16'b0011001010001011;
                14'h423 	:	o_val <= 16'b0011001010010110;
                14'h424 	:	o_val <= 16'b0011001010100010;
                14'h425 	:	o_val <= 16'b0011001010101101;
                14'h426 	:	o_val <= 16'b0011001010111001;
                14'h427 	:	o_val <= 16'b0011001011000100;
                14'h428 	:	o_val <= 16'b0011001011010000;
                14'h429 	:	o_val <= 16'b0011001011011011;
                14'h42a 	:	o_val <= 16'b0011001011100111;
                14'h42b 	:	o_val <= 16'b0011001011110011;
                14'h42c 	:	o_val <= 16'b0011001011111110;
                14'h42d 	:	o_val <= 16'b0011001100001010;
                14'h42e 	:	o_val <= 16'b0011001100010101;
                14'h42f 	:	o_val <= 16'b0011001100100001;
                14'h430 	:	o_val <= 16'b0011001100101100;
                14'h431 	:	o_val <= 16'b0011001100111000;
                14'h432 	:	o_val <= 16'b0011001101000011;
                14'h433 	:	o_val <= 16'b0011001101001111;
                14'h434 	:	o_val <= 16'b0011001101011010;
                14'h435 	:	o_val <= 16'b0011001101100110;
                14'h436 	:	o_val <= 16'b0011001101110001;
                14'h437 	:	o_val <= 16'b0011001101111101;
                14'h438 	:	o_val <= 16'b0011001110001000;
                14'h439 	:	o_val <= 16'b0011001110010100;
                14'h43a 	:	o_val <= 16'b0011001110011111;
                14'h43b 	:	o_val <= 16'b0011001110101011;
                14'h43c 	:	o_val <= 16'b0011001110110110;
                14'h43d 	:	o_val <= 16'b0011001111000010;
                14'h43e 	:	o_val <= 16'b0011001111001101;
                14'h43f 	:	o_val <= 16'b0011001111011001;
                14'h440 	:	o_val <= 16'b0011001111100100;
                14'h441 	:	o_val <= 16'b0011001111110000;
                14'h442 	:	o_val <= 16'b0011001111111011;
                14'h443 	:	o_val <= 16'b0011010000000111;
                14'h444 	:	o_val <= 16'b0011010000010010;
                14'h445 	:	o_val <= 16'b0011010000011110;
                14'h446 	:	o_val <= 16'b0011010000101001;
                14'h447 	:	o_val <= 16'b0011010000110101;
                14'h448 	:	o_val <= 16'b0011010001000000;
                14'h449 	:	o_val <= 16'b0011010001001011;
                14'h44a 	:	o_val <= 16'b0011010001010111;
                14'h44b 	:	o_val <= 16'b0011010001100010;
                14'h44c 	:	o_val <= 16'b0011010001101110;
                14'h44d 	:	o_val <= 16'b0011010001111001;
                14'h44e 	:	o_val <= 16'b0011010010000101;
                14'h44f 	:	o_val <= 16'b0011010010010000;
                14'h450 	:	o_val <= 16'b0011010010011100;
                14'h451 	:	o_val <= 16'b0011010010100111;
                14'h452 	:	o_val <= 16'b0011010010110011;
                14'h453 	:	o_val <= 16'b0011010010111110;
                14'h454 	:	o_val <= 16'b0011010011001010;
                14'h455 	:	o_val <= 16'b0011010011010101;
                14'h456 	:	o_val <= 16'b0011010011100000;
                14'h457 	:	o_val <= 16'b0011010011101100;
                14'h458 	:	o_val <= 16'b0011010011110111;
                14'h459 	:	o_val <= 16'b0011010100000011;
                14'h45a 	:	o_val <= 16'b0011010100001110;
                14'h45b 	:	o_val <= 16'b0011010100011010;
                14'h45c 	:	o_val <= 16'b0011010100100101;
                14'h45d 	:	o_val <= 16'b0011010100110000;
                14'h45e 	:	o_val <= 16'b0011010100111100;
                14'h45f 	:	o_val <= 16'b0011010101000111;
                14'h460 	:	o_val <= 16'b0011010101010011;
                14'h461 	:	o_val <= 16'b0011010101011110;
                14'h462 	:	o_val <= 16'b0011010101101010;
                14'h463 	:	o_val <= 16'b0011010101110101;
                14'h464 	:	o_val <= 16'b0011010110000000;
                14'h465 	:	o_val <= 16'b0011010110001100;
                14'h466 	:	o_val <= 16'b0011010110010111;
                14'h467 	:	o_val <= 16'b0011010110100011;
                14'h468 	:	o_val <= 16'b0011010110101110;
                14'h469 	:	o_val <= 16'b0011010110111010;
                14'h46a 	:	o_val <= 16'b0011010111000101;
                14'h46b 	:	o_val <= 16'b0011010111010000;
                14'h46c 	:	o_val <= 16'b0011010111011100;
                14'h46d 	:	o_val <= 16'b0011010111100111;
                14'h46e 	:	o_val <= 16'b0011010111110011;
                14'h46f 	:	o_val <= 16'b0011010111111110;
                14'h470 	:	o_val <= 16'b0011011000001001;
                14'h471 	:	o_val <= 16'b0011011000010101;
                14'h472 	:	o_val <= 16'b0011011000100000;
                14'h473 	:	o_val <= 16'b0011011000101011;
                14'h474 	:	o_val <= 16'b0011011000110111;
                14'h475 	:	o_val <= 16'b0011011001000010;
                14'h476 	:	o_val <= 16'b0011011001001110;
                14'h477 	:	o_val <= 16'b0011011001011001;
                14'h478 	:	o_val <= 16'b0011011001100100;
                14'h479 	:	o_val <= 16'b0011011001110000;
                14'h47a 	:	o_val <= 16'b0011011001111011;
                14'h47b 	:	o_val <= 16'b0011011010000110;
                14'h47c 	:	o_val <= 16'b0011011010010010;
                14'h47d 	:	o_val <= 16'b0011011010011101;
                14'h47e 	:	o_val <= 16'b0011011010101001;
                14'h47f 	:	o_val <= 16'b0011011010110100;
                14'h480 	:	o_val <= 16'b0011011010111111;
                14'h481 	:	o_val <= 16'b0011011011001011;
                14'h482 	:	o_val <= 16'b0011011011010110;
                14'h483 	:	o_val <= 16'b0011011011100001;
                14'h484 	:	o_val <= 16'b0011011011101101;
                14'h485 	:	o_val <= 16'b0011011011111000;
                14'h486 	:	o_val <= 16'b0011011100000011;
                14'h487 	:	o_val <= 16'b0011011100001111;
                14'h488 	:	o_val <= 16'b0011011100011010;
                14'h489 	:	o_val <= 16'b0011011100100101;
                14'h48a 	:	o_val <= 16'b0011011100110001;
                14'h48b 	:	o_val <= 16'b0011011100111100;
                14'h48c 	:	o_val <= 16'b0011011101000111;
                14'h48d 	:	o_val <= 16'b0011011101010011;
                14'h48e 	:	o_val <= 16'b0011011101011110;
                14'h48f 	:	o_val <= 16'b0011011101101001;
                14'h490 	:	o_val <= 16'b0011011101110101;
                14'h491 	:	o_val <= 16'b0011011110000000;
                14'h492 	:	o_val <= 16'b0011011110001011;
                14'h493 	:	o_val <= 16'b0011011110010111;
                14'h494 	:	o_val <= 16'b0011011110100010;
                14'h495 	:	o_val <= 16'b0011011110101101;
                14'h496 	:	o_val <= 16'b0011011110111001;
                14'h497 	:	o_val <= 16'b0011011111000100;
                14'h498 	:	o_val <= 16'b0011011111001111;
                14'h499 	:	o_val <= 16'b0011011111011011;
                14'h49a 	:	o_val <= 16'b0011011111100110;
                14'h49b 	:	o_val <= 16'b0011011111110001;
                14'h49c 	:	o_val <= 16'b0011011111111101;
                14'h49d 	:	o_val <= 16'b0011100000001000;
                14'h49e 	:	o_val <= 16'b0011100000010011;
                14'h49f 	:	o_val <= 16'b0011100000011110;
                14'h4a0 	:	o_val <= 16'b0011100000101010;
                14'h4a1 	:	o_val <= 16'b0011100000110101;
                14'h4a2 	:	o_val <= 16'b0011100001000000;
                14'h4a3 	:	o_val <= 16'b0011100001001100;
                14'h4a4 	:	o_val <= 16'b0011100001010111;
                14'h4a5 	:	o_val <= 16'b0011100001100010;
                14'h4a6 	:	o_val <= 16'b0011100001101101;
                14'h4a7 	:	o_val <= 16'b0011100001111001;
                14'h4a8 	:	o_val <= 16'b0011100010000100;
                14'h4a9 	:	o_val <= 16'b0011100010001111;
                14'h4aa 	:	o_val <= 16'b0011100010011011;
                14'h4ab 	:	o_val <= 16'b0011100010100110;
                14'h4ac 	:	o_val <= 16'b0011100010110001;
                14'h4ad 	:	o_val <= 16'b0011100010111100;
                14'h4ae 	:	o_val <= 16'b0011100011001000;
                14'h4af 	:	o_val <= 16'b0011100011010011;
                14'h4b0 	:	o_val <= 16'b0011100011011110;
                14'h4b1 	:	o_val <= 16'b0011100011101001;
                14'h4b2 	:	o_val <= 16'b0011100011110101;
                14'h4b3 	:	o_val <= 16'b0011100100000000;
                14'h4b4 	:	o_val <= 16'b0011100100001011;
                14'h4b5 	:	o_val <= 16'b0011100100010110;
                14'h4b6 	:	o_val <= 16'b0011100100100010;
                14'h4b7 	:	o_val <= 16'b0011100100101101;
                14'h4b8 	:	o_val <= 16'b0011100100111000;
                14'h4b9 	:	o_val <= 16'b0011100101000011;
                14'h4ba 	:	o_val <= 16'b0011100101001111;
                14'h4bb 	:	o_val <= 16'b0011100101011010;
                14'h4bc 	:	o_val <= 16'b0011100101100101;
                14'h4bd 	:	o_val <= 16'b0011100101110000;
                14'h4be 	:	o_val <= 16'b0011100101111100;
                14'h4bf 	:	o_val <= 16'b0011100110000111;
                14'h4c0 	:	o_val <= 16'b0011100110010010;
                14'h4c1 	:	o_val <= 16'b0011100110011101;
                14'h4c2 	:	o_val <= 16'b0011100110101000;
                14'h4c3 	:	o_val <= 16'b0011100110110100;
                14'h4c4 	:	o_val <= 16'b0011100110111111;
                14'h4c5 	:	o_val <= 16'b0011100111001010;
                14'h4c6 	:	o_val <= 16'b0011100111010101;
                14'h4c7 	:	o_val <= 16'b0011100111100000;
                14'h4c8 	:	o_val <= 16'b0011100111101100;
                14'h4c9 	:	o_val <= 16'b0011100111110111;
                14'h4ca 	:	o_val <= 16'b0011101000000010;
                14'h4cb 	:	o_val <= 16'b0011101000001101;
                14'h4cc 	:	o_val <= 16'b0011101000011001;
                14'h4cd 	:	o_val <= 16'b0011101000100100;
                14'h4ce 	:	o_val <= 16'b0011101000101111;
                14'h4cf 	:	o_val <= 16'b0011101000111010;
                14'h4d0 	:	o_val <= 16'b0011101001000101;
                14'h4d1 	:	o_val <= 16'b0011101001010000;
                14'h4d2 	:	o_val <= 16'b0011101001011100;
                14'h4d3 	:	o_val <= 16'b0011101001100111;
                14'h4d4 	:	o_val <= 16'b0011101001110010;
                14'h4d5 	:	o_val <= 16'b0011101001111101;
                14'h4d6 	:	o_val <= 16'b0011101010001000;
                14'h4d7 	:	o_val <= 16'b0011101010010100;
                14'h4d8 	:	o_val <= 16'b0011101010011111;
                14'h4d9 	:	o_val <= 16'b0011101010101010;
                14'h4da 	:	o_val <= 16'b0011101010110101;
                14'h4db 	:	o_val <= 16'b0011101011000000;
                14'h4dc 	:	o_val <= 16'b0011101011001011;
                14'h4dd 	:	o_val <= 16'b0011101011010111;
                14'h4de 	:	o_val <= 16'b0011101011100010;
                14'h4df 	:	o_val <= 16'b0011101011101101;
                14'h4e0 	:	o_val <= 16'b0011101011111000;
                14'h4e1 	:	o_val <= 16'b0011101100000011;
                14'h4e2 	:	o_val <= 16'b0011101100001110;
                14'h4e3 	:	o_val <= 16'b0011101100011001;
                14'h4e4 	:	o_val <= 16'b0011101100100101;
                14'h4e5 	:	o_val <= 16'b0011101100110000;
                14'h4e6 	:	o_val <= 16'b0011101100111011;
                14'h4e7 	:	o_val <= 16'b0011101101000110;
                14'h4e8 	:	o_val <= 16'b0011101101010001;
                14'h4e9 	:	o_val <= 16'b0011101101011100;
                14'h4ea 	:	o_val <= 16'b0011101101100111;
                14'h4eb 	:	o_val <= 16'b0011101101110011;
                14'h4ec 	:	o_val <= 16'b0011101101111110;
                14'h4ed 	:	o_val <= 16'b0011101110001001;
                14'h4ee 	:	o_val <= 16'b0011101110010100;
                14'h4ef 	:	o_val <= 16'b0011101110011111;
                14'h4f0 	:	o_val <= 16'b0011101110101010;
                14'h4f1 	:	o_val <= 16'b0011101110110101;
                14'h4f2 	:	o_val <= 16'b0011101111000000;
                14'h4f3 	:	o_val <= 16'b0011101111001100;
                14'h4f4 	:	o_val <= 16'b0011101111010111;
                14'h4f5 	:	o_val <= 16'b0011101111100010;
                14'h4f6 	:	o_val <= 16'b0011101111101101;
                14'h4f7 	:	o_val <= 16'b0011101111111000;
                14'h4f8 	:	o_val <= 16'b0011110000000011;
                14'h4f9 	:	o_val <= 16'b0011110000001110;
                14'h4fa 	:	o_val <= 16'b0011110000011001;
                14'h4fb 	:	o_val <= 16'b0011110000100100;
                14'h4fc 	:	o_val <= 16'b0011110000101111;
                14'h4fd 	:	o_val <= 16'b0011110000111011;
                14'h4fe 	:	o_val <= 16'b0011110001000110;
                14'h4ff 	:	o_val <= 16'b0011110001010001;
                14'h500 	:	o_val <= 16'b0011110001011100;
                14'h501 	:	o_val <= 16'b0011110001100111;
                14'h502 	:	o_val <= 16'b0011110001110010;
                14'h503 	:	o_val <= 16'b0011110001111101;
                14'h504 	:	o_val <= 16'b0011110010001000;
                14'h505 	:	o_val <= 16'b0011110010010011;
                14'h506 	:	o_val <= 16'b0011110010011110;
                14'h507 	:	o_val <= 16'b0011110010101001;
                14'h508 	:	o_val <= 16'b0011110010110100;
                14'h509 	:	o_val <= 16'b0011110010111111;
                14'h50a 	:	o_val <= 16'b0011110011001010;
                14'h50b 	:	o_val <= 16'b0011110011010110;
                14'h50c 	:	o_val <= 16'b0011110011100001;
                14'h50d 	:	o_val <= 16'b0011110011101100;
                14'h50e 	:	o_val <= 16'b0011110011110111;
                14'h50f 	:	o_val <= 16'b0011110100000010;
                14'h510 	:	o_val <= 16'b0011110100001101;
                14'h511 	:	o_val <= 16'b0011110100011000;
                14'h512 	:	o_val <= 16'b0011110100100011;
                14'h513 	:	o_val <= 16'b0011110100101110;
                14'h514 	:	o_val <= 16'b0011110100111001;
                14'h515 	:	o_val <= 16'b0011110101000100;
                14'h516 	:	o_val <= 16'b0011110101001111;
                14'h517 	:	o_val <= 16'b0011110101011010;
                14'h518 	:	o_val <= 16'b0011110101100101;
                14'h519 	:	o_val <= 16'b0011110101110000;
                14'h51a 	:	o_val <= 16'b0011110101111011;
                14'h51b 	:	o_val <= 16'b0011110110000110;
                14'h51c 	:	o_val <= 16'b0011110110010001;
                14'h51d 	:	o_val <= 16'b0011110110011100;
                14'h51e 	:	o_val <= 16'b0011110110100111;
                14'h51f 	:	o_val <= 16'b0011110110110010;
                14'h520 	:	o_val <= 16'b0011110110111101;
                14'h521 	:	o_val <= 16'b0011110111001000;
                14'h522 	:	o_val <= 16'b0011110111010011;
                14'h523 	:	o_val <= 16'b0011110111011110;
                14'h524 	:	o_val <= 16'b0011110111101001;
                14'h525 	:	o_val <= 16'b0011110111110100;
                14'h526 	:	o_val <= 16'b0011110111111111;
                14'h527 	:	o_val <= 16'b0011111000001010;
                14'h528 	:	o_val <= 16'b0011111000010101;
                14'h529 	:	o_val <= 16'b0011111000100000;
                14'h52a 	:	o_val <= 16'b0011111000101011;
                14'h52b 	:	o_val <= 16'b0011111000110110;
                14'h52c 	:	o_val <= 16'b0011111001000001;
                14'h52d 	:	o_val <= 16'b0011111001001100;
                14'h52e 	:	o_val <= 16'b0011111001010111;
                14'h52f 	:	o_val <= 16'b0011111001100010;
                14'h530 	:	o_val <= 16'b0011111001101101;
                14'h531 	:	o_val <= 16'b0011111001111000;
                14'h532 	:	o_val <= 16'b0011111010000011;
                14'h533 	:	o_val <= 16'b0011111010001110;
                14'h534 	:	o_val <= 16'b0011111010011001;
                14'h535 	:	o_val <= 16'b0011111010100100;
                14'h536 	:	o_val <= 16'b0011111010101111;
                14'h537 	:	o_val <= 16'b0011111010111010;
                14'h538 	:	o_val <= 16'b0011111011000101;
                14'h539 	:	o_val <= 16'b0011111011010000;
                14'h53a 	:	o_val <= 16'b0011111011011011;
                14'h53b 	:	o_val <= 16'b0011111011100110;
                14'h53c 	:	o_val <= 16'b0011111011110001;
                14'h53d 	:	o_val <= 16'b0011111011111011;
                14'h53e 	:	o_val <= 16'b0011111100000110;
                14'h53f 	:	o_val <= 16'b0011111100010001;
                14'h540 	:	o_val <= 16'b0011111100011100;
                14'h541 	:	o_val <= 16'b0011111100100111;
                14'h542 	:	o_val <= 16'b0011111100110010;
                14'h543 	:	o_val <= 16'b0011111100111101;
                14'h544 	:	o_val <= 16'b0011111101001000;
                14'h545 	:	o_val <= 16'b0011111101010011;
                14'h546 	:	o_val <= 16'b0011111101011110;
                14'h547 	:	o_val <= 16'b0011111101101001;
                14'h548 	:	o_val <= 16'b0011111101110100;
                14'h549 	:	o_val <= 16'b0011111101111111;
                14'h54a 	:	o_val <= 16'b0011111110001001;
                14'h54b 	:	o_val <= 16'b0011111110010100;
                14'h54c 	:	o_val <= 16'b0011111110011111;
                14'h54d 	:	o_val <= 16'b0011111110101010;
                14'h54e 	:	o_val <= 16'b0011111110110101;
                14'h54f 	:	o_val <= 16'b0011111111000000;
                14'h550 	:	o_val <= 16'b0011111111001011;
                14'h551 	:	o_val <= 16'b0011111111010110;
                14'h552 	:	o_val <= 16'b0011111111100001;
                14'h553 	:	o_val <= 16'b0011111111101100;
                14'h554 	:	o_val <= 16'b0011111111110110;
                14'h555 	:	o_val <= 16'b0100000000000001;
                14'h556 	:	o_val <= 16'b0100000000001100;
                14'h557 	:	o_val <= 16'b0100000000010111;
                14'h558 	:	o_val <= 16'b0100000000100010;
                14'h559 	:	o_val <= 16'b0100000000101101;
                14'h55a 	:	o_val <= 16'b0100000000111000;
                14'h55b 	:	o_val <= 16'b0100000001000011;
                14'h55c 	:	o_val <= 16'b0100000001001101;
                14'h55d 	:	o_val <= 16'b0100000001011000;
                14'h55e 	:	o_val <= 16'b0100000001100011;
                14'h55f 	:	o_val <= 16'b0100000001101110;
                14'h560 	:	o_val <= 16'b0100000001111001;
                14'h561 	:	o_val <= 16'b0100000010000100;
                14'h562 	:	o_val <= 16'b0100000010001111;
                14'h563 	:	o_val <= 16'b0100000010011001;
                14'h564 	:	o_val <= 16'b0100000010100100;
                14'h565 	:	o_val <= 16'b0100000010101111;
                14'h566 	:	o_val <= 16'b0100000010111010;
                14'h567 	:	o_val <= 16'b0100000011000101;
                14'h568 	:	o_val <= 16'b0100000011010000;
                14'h569 	:	o_val <= 16'b0100000011011010;
                14'h56a 	:	o_val <= 16'b0100000011100101;
                14'h56b 	:	o_val <= 16'b0100000011110000;
                14'h56c 	:	o_val <= 16'b0100000011111011;
                14'h56d 	:	o_val <= 16'b0100000100000110;
                14'h56e 	:	o_val <= 16'b0100000100010001;
                14'h56f 	:	o_val <= 16'b0100000100011011;
                14'h570 	:	o_val <= 16'b0100000100100110;
                14'h571 	:	o_val <= 16'b0100000100110001;
                14'h572 	:	o_val <= 16'b0100000100111100;
                14'h573 	:	o_val <= 16'b0100000101000111;
                14'h574 	:	o_val <= 16'b0100000101010010;
                14'h575 	:	o_val <= 16'b0100000101011100;
                14'h576 	:	o_val <= 16'b0100000101100111;
                14'h577 	:	o_val <= 16'b0100000101110010;
                14'h578 	:	o_val <= 16'b0100000101111101;
                14'h579 	:	o_val <= 16'b0100000110001000;
                14'h57a 	:	o_val <= 16'b0100000110010010;
                14'h57b 	:	o_val <= 16'b0100000110011101;
                14'h57c 	:	o_val <= 16'b0100000110101000;
                14'h57d 	:	o_val <= 16'b0100000110110011;
                14'h57e 	:	o_val <= 16'b0100000110111101;
                14'h57f 	:	o_val <= 16'b0100000111001000;
                14'h580 	:	o_val <= 16'b0100000111010011;
                14'h581 	:	o_val <= 16'b0100000111011110;
                14'h582 	:	o_val <= 16'b0100000111101001;
                14'h583 	:	o_val <= 16'b0100000111110011;
                14'h584 	:	o_val <= 16'b0100000111111110;
                14'h585 	:	o_val <= 16'b0100001000001001;
                14'h586 	:	o_val <= 16'b0100001000010100;
                14'h587 	:	o_val <= 16'b0100001000011110;
                14'h588 	:	o_val <= 16'b0100001000101001;
                14'h589 	:	o_val <= 16'b0100001000110100;
                14'h58a 	:	o_val <= 16'b0100001000111111;
                14'h58b 	:	o_val <= 16'b0100001001001001;
                14'h58c 	:	o_val <= 16'b0100001001010100;
                14'h58d 	:	o_val <= 16'b0100001001011111;
                14'h58e 	:	o_val <= 16'b0100001001101010;
                14'h58f 	:	o_val <= 16'b0100001001110100;
                14'h590 	:	o_val <= 16'b0100001001111111;
                14'h591 	:	o_val <= 16'b0100001010001010;
                14'h592 	:	o_val <= 16'b0100001010010101;
                14'h593 	:	o_val <= 16'b0100001010011111;
                14'h594 	:	o_val <= 16'b0100001010101010;
                14'h595 	:	o_val <= 16'b0100001010110101;
                14'h596 	:	o_val <= 16'b0100001011000000;
                14'h597 	:	o_val <= 16'b0100001011001010;
                14'h598 	:	o_val <= 16'b0100001011010101;
                14'h599 	:	o_val <= 16'b0100001011100000;
                14'h59a 	:	o_val <= 16'b0100001011101010;
                14'h59b 	:	o_val <= 16'b0100001011110101;
                14'h59c 	:	o_val <= 16'b0100001100000000;
                14'h59d 	:	o_val <= 16'b0100001100001011;
                14'h59e 	:	o_val <= 16'b0100001100010101;
                14'h59f 	:	o_val <= 16'b0100001100100000;
                14'h5a0 	:	o_val <= 16'b0100001100101011;
                14'h5a1 	:	o_val <= 16'b0100001100110101;
                14'h5a2 	:	o_val <= 16'b0100001101000000;
                14'h5a3 	:	o_val <= 16'b0100001101001011;
                14'h5a4 	:	o_val <= 16'b0100001101010101;
                14'h5a5 	:	o_val <= 16'b0100001101100000;
                14'h5a6 	:	o_val <= 16'b0100001101101011;
                14'h5a7 	:	o_val <= 16'b0100001101110101;
                14'h5a8 	:	o_val <= 16'b0100001110000000;
                14'h5a9 	:	o_val <= 16'b0100001110001011;
                14'h5aa 	:	o_val <= 16'b0100001110010101;
                14'h5ab 	:	o_val <= 16'b0100001110100000;
                14'h5ac 	:	o_val <= 16'b0100001110101011;
                14'h5ad 	:	o_val <= 16'b0100001110110101;
                14'h5ae 	:	o_val <= 16'b0100001111000000;
                14'h5af 	:	o_val <= 16'b0100001111001011;
                14'h5b0 	:	o_val <= 16'b0100001111010101;
                14'h5b1 	:	o_val <= 16'b0100001111100000;
                14'h5b2 	:	o_val <= 16'b0100001111101011;
                14'h5b3 	:	o_val <= 16'b0100001111110101;
                14'h5b4 	:	o_val <= 16'b0100010000000000;
                14'h5b5 	:	o_val <= 16'b0100010000001011;
                14'h5b6 	:	o_val <= 16'b0100010000010101;
                14'h5b7 	:	o_val <= 16'b0100010000100000;
                14'h5b8 	:	o_val <= 16'b0100010000101011;
                14'h5b9 	:	o_val <= 16'b0100010000110101;
                14'h5ba 	:	o_val <= 16'b0100010001000000;
                14'h5bb 	:	o_val <= 16'b0100010001001011;
                14'h5bc 	:	o_val <= 16'b0100010001010101;
                14'h5bd 	:	o_val <= 16'b0100010001100000;
                14'h5be 	:	o_val <= 16'b0100010001101010;
                14'h5bf 	:	o_val <= 16'b0100010001110101;
                14'h5c0 	:	o_val <= 16'b0100010010000000;
                14'h5c1 	:	o_val <= 16'b0100010010001010;
                14'h5c2 	:	o_val <= 16'b0100010010010101;
                14'h5c3 	:	o_val <= 16'b0100010010011111;
                14'h5c4 	:	o_val <= 16'b0100010010101010;
                14'h5c5 	:	o_val <= 16'b0100010010110101;
                14'h5c6 	:	o_val <= 16'b0100010010111111;
                14'h5c7 	:	o_val <= 16'b0100010011001010;
                14'h5c8 	:	o_val <= 16'b0100010011010100;
                14'h5c9 	:	o_val <= 16'b0100010011011111;
                14'h5ca 	:	o_val <= 16'b0100010011101010;
                14'h5cb 	:	o_val <= 16'b0100010011110100;
                14'h5cc 	:	o_val <= 16'b0100010011111111;
                14'h5cd 	:	o_val <= 16'b0100010100001001;
                14'h5ce 	:	o_val <= 16'b0100010100010100;
                14'h5cf 	:	o_val <= 16'b0100010100011111;
                14'h5d0 	:	o_val <= 16'b0100010100101001;
                14'h5d1 	:	o_val <= 16'b0100010100110100;
                14'h5d2 	:	o_val <= 16'b0100010100111110;
                14'h5d3 	:	o_val <= 16'b0100010101001001;
                14'h5d4 	:	o_val <= 16'b0100010101010011;
                14'h5d5 	:	o_val <= 16'b0100010101011110;
                14'h5d6 	:	o_val <= 16'b0100010101101001;
                14'h5d7 	:	o_val <= 16'b0100010101110011;
                14'h5d8 	:	o_val <= 16'b0100010101111110;
                14'h5d9 	:	o_val <= 16'b0100010110001000;
                14'h5da 	:	o_val <= 16'b0100010110010011;
                14'h5db 	:	o_val <= 16'b0100010110011101;
                14'h5dc 	:	o_val <= 16'b0100010110101000;
                14'h5dd 	:	o_val <= 16'b0100010110110010;
                14'h5de 	:	o_val <= 16'b0100010110111101;
                14'h5df 	:	o_val <= 16'b0100010111000111;
                14'h5e0 	:	o_val <= 16'b0100010111010010;
                14'h5e1 	:	o_val <= 16'b0100010111011101;
                14'h5e2 	:	o_val <= 16'b0100010111100111;
                14'h5e3 	:	o_val <= 16'b0100010111110010;
                14'h5e4 	:	o_val <= 16'b0100010111111100;
                14'h5e5 	:	o_val <= 16'b0100011000000111;
                14'h5e6 	:	o_val <= 16'b0100011000010001;
                14'h5e7 	:	o_val <= 16'b0100011000011100;
                14'h5e8 	:	o_val <= 16'b0100011000100110;
                14'h5e9 	:	o_val <= 16'b0100011000110001;
                14'h5ea 	:	o_val <= 16'b0100011000111011;
                14'h5eb 	:	o_val <= 16'b0100011001000110;
                14'h5ec 	:	o_val <= 16'b0100011001010000;
                14'h5ed 	:	o_val <= 16'b0100011001011011;
                14'h5ee 	:	o_val <= 16'b0100011001100101;
                14'h5ef 	:	o_val <= 16'b0100011001110000;
                14'h5f0 	:	o_val <= 16'b0100011001111010;
                14'h5f1 	:	o_val <= 16'b0100011010000101;
                14'h5f2 	:	o_val <= 16'b0100011010001111;
                14'h5f3 	:	o_val <= 16'b0100011010011010;
                14'h5f4 	:	o_val <= 16'b0100011010100100;
                14'h5f5 	:	o_val <= 16'b0100011010101111;
                14'h5f6 	:	o_val <= 16'b0100011010111001;
                14'h5f7 	:	o_val <= 16'b0100011011000100;
                14'h5f8 	:	o_val <= 16'b0100011011001110;
                14'h5f9 	:	o_val <= 16'b0100011011011000;
                14'h5fa 	:	o_val <= 16'b0100011011100011;
                14'h5fb 	:	o_val <= 16'b0100011011101101;
                14'h5fc 	:	o_val <= 16'b0100011011111000;
                14'h5fd 	:	o_val <= 16'b0100011100000010;
                14'h5fe 	:	o_val <= 16'b0100011100001101;
                14'h5ff 	:	o_val <= 16'b0100011100010111;
                14'h600 	:	o_val <= 16'b0100011100100010;
                14'h601 	:	o_val <= 16'b0100011100101100;
                14'h602 	:	o_val <= 16'b0100011100110111;
                14'h603 	:	o_val <= 16'b0100011101000001;
                14'h604 	:	o_val <= 16'b0100011101001011;
                14'h605 	:	o_val <= 16'b0100011101010110;
                14'h606 	:	o_val <= 16'b0100011101100000;
                14'h607 	:	o_val <= 16'b0100011101101011;
                14'h608 	:	o_val <= 16'b0100011101110101;
                14'h609 	:	o_val <= 16'b0100011110000000;
                14'h60a 	:	o_val <= 16'b0100011110001010;
                14'h60b 	:	o_val <= 16'b0100011110010100;
                14'h60c 	:	o_val <= 16'b0100011110011111;
                14'h60d 	:	o_val <= 16'b0100011110101001;
                14'h60e 	:	o_val <= 16'b0100011110110100;
                14'h60f 	:	o_val <= 16'b0100011110111110;
                14'h610 	:	o_val <= 16'b0100011111001000;
                14'h611 	:	o_val <= 16'b0100011111010011;
                14'h612 	:	o_val <= 16'b0100011111011101;
                14'h613 	:	o_val <= 16'b0100011111101000;
                14'h614 	:	o_val <= 16'b0100011111110010;
                14'h615 	:	o_val <= 16'b0100011111111100;
                14'h616 	:	o_val <= 16'b0100100000000111;
                14'h617 	:	o_val <= 16'b0100100000010001;
                14'h618 	:	o_val <= 16'b0100100000011100;
                14'h619 	:	o_val <= 16'b0100100000100110;
                14'h61a 	:	o_val <= 16'b0100100000110000;
                14'h61b 	:	o_val <= 16'b0100100000111011;
                14'h61c 	:	o_val <= 16'b0100100001000101;
                14'h61d 	:	o_val <= 16'b0100100001001111;
                14'h61e 	:	o_val <= 16'b0100100001011010;
                14'h61f 	:	o_val <= 16'b0100100001100100;
                14'h620 	:	o_val <= 16'b0100100001101111;
                14'h621 	:	o_val <= 16'b0100100001111001;
                14'h622 	:	o_val <= 16'b0100100010000011;
                14'h623 	:	o_val <= 16'b0100100010001110;
                14'h624 	:	o_val <= 16'b0100100010011000;
                14'h625 	:	o_val <= 16'b0100100010100010;
                14'h626 	:	o_val <= 16'b0100100010101101;
                14'h627 	:	o_val <= 16'b0100100010110111;
                14'h628 	:	o_val <= 16'b0100100011000001;
                14'h629 	:	o_val <= 16'b0100100011001100;
                14'h62a 	:	o_val <= 16'b0100100011010110;
                14'h62b 	:	o_val <= 16'b0100100011100000;
                14'h62c 	:	o_val <= 16'b0100100011101011;
                14'h62d 	:	o_val <= 16'b0100100011110101;
                14'h62e 	:	o_val <= 16'b0100100011111111;
                14'h62f 	:	o_val <= 16'b0100100100001010;
                14'h630 	:	o_val <= 16'b0100100100010100;
                14'h631 	:	o_val <= 16'b0100100100011110;
                14'h632 	:	o_val <= 16'b0100100100101001;
                14'h633 	:	o_val <= 16'b0100100100110011;
                14'h634 	:	o_val <= 16'b0100100100111101;
                14'h635 	:	o_val <= 16'b0100100101001000;
                14'h636 	:	o_val <= 16'b0100100101010010;
                14'h637 	:	o_val <= 16'b0100100101011100;
                14'h638 	:	o_val <= 16'b0100100101100110;
                14'h639 	:	o_val <= 16'b0100100101110001;
                14'h63a 	:	o_val <= 16'b0100100101111011;
                14'h63b 	:	o_val <= 16'b0100100110000101;
                14'h63c 	:	o_val <= 16'b0100100110010000;
                14'h63d 	:	o_val <= 16'b0100100110011010;
                14'h63e 	:	o_val <= 16'b0100100110100100;
                14'h63f 	:	o_val <= 16'b0100100110101110;
                14'h640 	:	o_val <= 16'b0100100110111001;
                14'h641 	:	o_val <= 16'b0100100111000011;
                14'h642 	:	o_val <= 16'b0100100111001101;
                14'h643 	:	o_val <= 16'b0100100111011000;
                14'h644 	:	o_val <= 16'b0100100111100010;
                14'h645 	:	o_val <= 16'b0100100111101100;
                14'h646 	:	o_val <= 16'b0100100111110110;
                14'h647 	:	o_val <= 16'b0100101000000001;
                14'h648 	:	o_val <= 16'b0100101000001011;
                14'h649 	:	o_val <= 16'b0100101000010101;
                14'h64a 	:	o_val <= 16'b0100101000011111;
                14'h64b 	:	o_val <= 16'b0100101000101010;
                14'h64c 	:	o_val <= 16'b0100101000110100;
                14'h64d 	:	o_val <= 16'b0100101000111110;
                14'h64e 	:	o_val <= 16'b0100101001001000;
                14'h64f 	:	o_val <= 16'b0100101001010010;
                14'h650 	:	o_val <= 16'b0100101001011101;
                14'h651 	:	o_val <= 16'b0100101001100111;
                14'h652 	:	o_val <= 16'b0100101001110001;
                14'h653 	:	o_val <= 16'b0100101001111011;
                14'h654 	:	o_val <= 16'b0100101010000110;
                14'h655 	:	o_val <= 16'b0100101010010000;
                14'h656 	:	o_val <= 16'b0100101010011010;
                14'h657 	:	o_val <= 16'b0100101010100100;
                14'h658 	:	o_val <= 16'b0100101010101110;
                14'h659 	:	o_val <= 16'b0100101010111001;
                14'h65a 	:	o_val <= 16'b0100101011000011;
                14'h65b 	:	o_val <= 16'b0100101011001101;
                14'h65c 	:	o_val <= 16'b0100101011010111;
                14'h65d 	:	o_val <= 16'b0100101011100001;
                14'h65e 	:	o_val <= 16'b0100101011101100;
                14'h65f 	:	o_val <= 16'b0100101011110110;
                14'h660 	:	o_val <= 16'b0100101100000000;
                14'h661 	:	o_val <= 16'b0100101100001010;
                14'h662 	:	o_val <= 16'b0100101100010100;
                14'h663 	:	o_val <= 16'b0100101100011111;
                14'h664 	:	o_val <= 16'b0100101100101001;
                14'h665 	:	o_val <= 16'b0100101100110011;
                14'h666 	:	o_val <= 16'b0100101100111101;
                14'h667 	:	o_val <= 16'b0100101101000111;
                14'h668 	:	o_val <= 16'b0100101101010001;
                14'h669 	:	o_val <= 16'b0100101101011100;
                14'h66a 	:	o_val <= 16'b0100101101100110;
                14'h66b 	:	o_val <= 16'b0100101101110000;
                14'h66c 	:	o_val <= 16'b0100101101111010;
                14'h66d 	:	o_val <= 16'b0100101110000100;
                14'h66e 	:	o_val <= 16'b0100101110001110;
                14'h66f 	:	o_val <= 16'b0100101110011000;
                14'h670 	:	o_val <= 16'b0100101110100011;
                14'h671 	:	o_val <= 16'b0100101110101101;
                14'h672 	:	o_val <= 16'b0100101110110111;
                14'h673 	:	o_val <= 16'b0100101111000001;
                14'h674 	:	o_val <= 16'b0100101111001011;
                14'h675 	:	o_val <= 16'b0100101111010101;
                14'h676 	:	o_val <= 16'b0100101111011111;
                14'h677 	:	o_val <= 16'b0100101111101001;
                14'h678 	:	o_val <= 16'b0100101111110100;
                14'h679 	:	o_val <= 16'b0100101111111110;
                14'h67a 	:	o_val <= 16'b0100110000001000;
                14'h67b 	:	o_val <= 16'b0100110000010010;
                14'h67c 	:	o_val <= 16'b0100110000011100;
                14'h67d 	:	o_val <= 16'b0100110000100110;
                14'h67e 	:	o_val <= 16'b0100110000110000;
                14'h67f 	:	o_val <= 16'b0100110000111010;
                14'h680 	:	o_val <= 16'b0100110001000100;
                14'h681 	:	o_val <= 16'b0100110001001111;
                14'h682 	:	o_val <= 16'b0100110001011001;
                14'h683 	:	o_val <= 16'b0100110001100011;
                14'h684 	:	o_val <= 16'b0100110001101101;
                14'h685 	:	o_val <= 16'b0100110001110111;
                14'h686 	:	o_val <= 16'b0100110010000001;
                14'h687 	:	o_val <= 16'b0100110010001011;
                14'h688 	:	o_val <= 16'b0100110010010101;
                14'h689 	:	o_val <= 16'b0100110010011111;
                14'h68a 	:	o_val <= 16'b0100110010101001;
                14'h68b 	:	o_val <= 16'b0100110010110011;
                14'h68c 	:	o_val <= 16'b0100110010111101;
                14'h68d 	:	o_val <= 16'b0100110011000111;
                14'h68e 	:	o_val <= 16'b0100110011010001;
                14'h68f 	:	o_val <= 16'b0100110011011011;
                14'h690 	:	o_val <= 16'b0100110011100110;
                14'h691 	:	o_val <= 16'b0100110011110000;
                14'h692 	:	o_val <= 16'b0100110011111010;
                14'h693 	:	o_val <= 16'b0100110100000100;
                14'h694 	:	o_val <= 16'b0100110100001110;
                14'h695 	:	o_val <= 16'b0100110100011000;
                14'h696 	:	o_val <= 16'b0100110100100010;
                14'h697 	:	o_val <= 16'b0100110100101100;
                14'h698 	:	o_val <= 16'b0100110100110110;
                14'h699 	:	o_val <= 16'b0100110101000000;
                14'h69a 	:	o_val <= 16'b0100110101001010;
                14'h69b 	:	o_val <= 16'b0100110101010100;
                14'h69c 	:	o_val <= 16'b0100110101011110;
                14'h69d 	:	o_val <= 16'b0100110101101000;
                14'h69e 	:	o_val <= 16'b0100110101110010;
                14'h69f 	:	o_val <= 16'b0100110101111100;
                14'h6a0 	:	o_val <= 16'b0100110110000110;
                14'h6a1 	:	o_val <= 16'b0100110110010000;
                14'h6a2 	:	o_val <= 16'b0100110110011010;
                14'h6a3 	:	o_val <= 16'b0100110110100100;
                14'h6a4 	:	o_val <= 16'b0100110110101110;
                14'h6a5 	:	o_val <= 16'b0100110110111000;
                14'h6a6 	:	o_val <= 16'b0100110111000010;
                14'h6a7 	:	o_val <= 16'b0100110111001100;
                14'h6a8 	:	o_val <= 16'b0100110111010110;
                14'h6a9 	:	o_val <= 16'b0100110111100000;
                14'h6aa 	:	o_val <= 16'b0100110111101010;
                14'h6ab 	:	o_val <= 16'b0100110111110100;
                14'h6ac 	:	o_val <= 16'b0100110111111110;
                14'h6ad 	:	o_val <= 16'b0100111000001000;
                14'h6ae 	:	o_val <= 16'b0100111000010010;
                14'h6af 	:	o_val <= 16'b0100111000011100;
                14'h6b0 	:	o_val <= 16'b0100111000100110;
                14'h6b1 	:	o_val <= 16'b0100111000101111;
                14'h6b2 	:	o_val <= 16'b0100111000111001;
                14'h6b3 	:	o_val <= 16'b0100111001000011;
                14'h6b4 	:	o_val <= 16'b0100111001001101;
                14'h6b5 	:	o_val <= 16'b0100111001010111;
                14'h6b6 	:	o_val <= 16'b0100111001100001;
                14'h6b7 	:	o_val <= 16'b0100111001101011;
                14'h6b8 	:	o_val <= 16'b0100111001110101;
                14'h6b9 	:	o_val <= 16'b0100111001111111;
                14'h6ba 	:	o_val <= 16'b0100111010001001;
                14'h6bb 	:	o_val <= 16'b0100111010010011;
                14'h6bc 	:	o_val <= 16'b0100111010011101;
                14'h6bd 	:	o_val <= 16'b0100111010100111;
                14'h6be 	:	o_val <= 16'b0100111010110001;
                14'h6bf 	:	o_val <= 16'b0100111010111010;
                14'h6c0 	:	o_val <= 16'b0100111011000100;
                14'h6c1 	:	o_val <= 16'b0100111011001110;
                14'h6c2 	:	o_val <= 16'b0100111011011000;
                14'h6c3 	:	o_val <= 16'b0100111011100010;
                14'h6c4 	:	o_val <= 16'b0100111011101100;
                14'h6c5 	:	o_val <= 16'b0100111011110110;
                14'h6c6 	:	o_val <= 16'b0100111100000000;
                14'h6c7 	:	o_val <= 16'b0100111100001010;
                14'h6c8 	:	o_val <= 16'b0100111100010100;
                14'h6c9 	:	o_val <= 16'b0100111100011101;
                14'h6ca 	:	o_val <= 16'b0100111100100111;
                14'h6cb 	:	o_val <= 16'b0100111100110001;
                14'h6cc 	:	o_val <= 16'b0100111100111011;
                14'h6cd 	:	o_val <= 16'b0100111101000101;
                14'h6ce 	:	o_val <= 16'b0100111101001111;
                14'h6cf 	:	o_val <= 16'b0100111101011001;
                14'h6d0 	:	o_val <= 16'b0100111101100010;
                14'h6d1 	:	o_val <= 16'b0100111101101100;
                14'h6d2 	:	o_val <= 16'b0100111101110110;
                14'h6d3 	:	o_val <= 16'b0100111110000000;
                14'h6d4 	:	o_val <= 16'b0100111110001010;
                14'h6d5 	:	o_val <= 16'b0100111110010100;
                14'h6d6 	:	o_val <= 16'b0100111110011110;
                14'h6d7 	:	o_val <= 16'b0100111110100111;
                14'h6d8 	:	o_val <= 16'b0100111110110001;
                14'h6d9 	:	o_val <= 16'b0100111110111011;
                14'h6da 	:	o_val <= 16'b0100111111000101;
                14'h6db 	:	o_val <= 16'b0100111111001111;
                14'h6dc 	:	o_val <= 16'b0100111111011001;
                14'h6dd 	:	o_val <= 16'b0100111111100010;
                14'h6de 	:	o_val <= 16'b0100111111101100;
                14'h6df 	:	o_val <= 16'b0100111111110110;
                14'h6e0 	:	o_val <= 16'b0101000000000000;
                14'h6e1 	:	o_val <= 16'b0101000000001010;
                14'h6e2 	:	o_val <= 16'b0101000000010011;
                14'h6e3 	:	o_val <= 16'b0101000000011101;
                14'h6e4 	:	o_val <= 16'b0101000000100111;
                14'h6e5 	:	o_val <= 16'b0101000000110001;
                14'h6e6 	:	o_val <= 16'b0101000000111011;
                14'h6e7 	:	o_val <= 16'b0101000001000100;
                14'h6e8 	:	o_val <= 16'b0101000001001110;
                14'h6e9 	:	o_val <= 16'b0101000001011000;
                14'h6ea 	:	o_val <= 16'b0101000001100010;
                14'h6eb 	:	o_val <= 16'b0101000001101100;
                14'h6ec 	:	o_val <= 16'b0101000001110101;
                14'h6ed 	:	o_val <= 16'b0101000001111111;
                14'h6ee 	:	o_val <= 16'b0101000010001001;
                14'h6ef 	:	o_val <= 16'b0101000010010011;
                14'h6f0 	:	o_val <= 16'b0101000010011100;
                14'h6f1 	:	o_val <= 16'b0101000010100110;
                14'h6f2 	:	o_val <= 16'b0101000010110000;
                14'h6f3 	:	o_val <= 16'b0101000010111010;
                14'h6f4 	:	o_val <= 16'b0101000011000011;
                14'h6f5 	:	o_val <= 16'b0101000011001101;
                14'h6f6 	:	o_val <= 16'b0101000011010111;
                14'h6f7 	:	o_val <= 16'b0101000011100001;
                14'h6f8 	:	o_val <= 16'b0101000011101010;
                14'h6f9 	:	o_val <= 16'b0101000011110100;
                14'h6fa 	:	o_val <= 16'b0101000011111110;
                14'h6fb 	:	o_val <= 16'b0101000100001000;
                14'h6fc 	:	o_val <= 16'b0101000100010001;
                14'h6fd 	:	o_val <= 16'b0101000100011011;
                14'h6fe 	:	o_val <= 16'b0101000100100101;
                14'h6ff 	:	o_val <= 16'b0101000100101110;
                14'h700 	:	o_val <= 16'b0101000100111000;
                14'h701 	:	o_val <= 16'b0101000101000010;
                14'h702 	:	o_val <= 16'b0101000101001100;
                14'h703 	:	o_val <= 16'b0101000101010101;
                14'h704 	:	o_val <= 16'b0101000101011111;
                14'h705 	:	o_val <= 16'b0101000101101001;
                14'h706 	:	o_val <= 16'b0101000101110010;
                14'h707 	:	o_val <= 16'b0101000101111100;
                14'h708 	:	o_val <= 16'b0101000110000110;
                14'h709 	:	o_val <= 16'b0101000110001111;
                14'h70a 	:	o_val <= 16'b0101000110011001;
                14'h70b 	:	o_val <= 16'b0101000110100011;
                14'h70c 	:	o_val <= 16'b0101000110101100;
                14'h70d 	:	o_val <= 16'b0101000110110110;
                14'h70e 	:	o_val <= 16'b0101000111000000;
                14'h70f 	:	o_val <= 16'b0101000111001001;
                14'h710 	:	o_val <= 16'b0101000111010011;
                14'h711 	:	o_val <= 16'b0101000111011101;
                14'h712 	:	o_val <= 16'b0101000111100110;
                14'h713 	:	o_val <= 16'b0101000111110000;
                14'h714 	:	o_val <= 16'b0101000111111010;
                14'h715 	:	o_val <= 16'b0101001000000011;
                14'h716 	:	o_val <= 16'b0101001000001101;
                14'h717 	:	o_val <= 16'b0101001000010111;
                14'h718 	:	o_val <= 16'b0101001000100000;
                14'h719 	:	o_val <= 16'b0101001000101010;
                14'h71a 	:	o_val <= 16'b0101001000110100;
                14'h71b 	:	o_val <= 16'b0101001000111101;
                14'h71c 	:	o_val <= 16'b0101001001000111;
                14'h71d 	:	o_val <= 16'b0101001001010001;
                14'h71e 	:	o_val <= 16'b0101001001011010;
                14'h71f 	:	o_val <= 16'b0101001001100100;
                14'h720 	:	o_val <= 16'b0101001001101101;
                14'h721 	:	o_val <= 16'b0101001001110111;
                14'h722 	:	o_val <= 16'b0101001010000001;
                14'h723 	:	o_val <= 16'b0101001010001010;
                14'h724 	:	o_val <= 16'b0101001010010100;
                14'h725 	:	o_val <= 16'b0101001010011101;
                14'h726 	:	o_val <= 16'b0101001010100111;
                14'h727 	:	o_val <= 16'b0101001010110001;
                14'h728 	:	o_val <= 16'b0101001010111010;
                14'h729 	:	o_val <= 16'b0101001011000100;
                14'h72a 	:	o_val <= 16'b0101001011001101;
                14'h72b 	:	o_val <= 16'b0101001011010111;
                14'h72c 	:	o_val <= 16'b0101001011100001;
                14'h72d 	:	o_val <= 16'b0101001011101010;
                14'h72e 	:	o_val <= 16'b0101001011110100;
                14'h72f 	:	o_val <= 16'b0101001011111101;
                14'h730 	:	o_val <= 16'b0101001100000111;
                14'h731 	:	o_val <= 16'b0101001100010000;
                14'h732 	:	o_val <= 16'b0101001100011010;
                14'h733 	:	o_val <= 16'b0101001100100011;
                14'h734 	:	o_val <= 16'b0101001100101101;
                14'h735 	:	o_val <= 16'b0101001100110111;
                14'h736 	:	o_val <= 16'b0101001101000000;
                14'h737 	:	o_val <= 16'b0101001101001010;
                14'h738 	:	o_val <= 16'b0101001101010011;
                14'h739 	:	o_val <= 16'b0101001101011101;
                14'h73a 	:	o_val <= 16'b0101001101100110;
                14'h73b 	:	o_val <= 16'b0101001101110000;
                14'h73c 	:	o_val <= 16'b0101001101111001;
                14'h73d 	:	o_val <= 16'b0101001110000011;
                14'h73e 	:	o_val <= 16'b0101001110001100;
                14'h73f 	:	o_val <= 16'b0101001110010110;
                14'h740 	:	o_val <= 16'b0101001110011111;
                14'h741 	:	o_val <= 16'b0101001110101001;
                14'h742 	:	o_val <= 16'b0101001110110010;
                14'h743 	:	o_val <= 16'b0101001110111100;
                14'h744 	:	o_val <= 16'b0101001111000101;
                14'h745 	:	o_val <= 16'b0101001111001111;
                14'h746 	:	o_val <= 16'b0101001111011000;
                14'h747 	:	o_val <= 16'b0101001111100010;
                14'h748 	:	o_val <= 16'b0101001111101011;
                14'h749 	:	o_val <= 16'b0101001111110101;
                14'h74a 	:	o_val <= 16'b0101001111111110;
                14'h74b 	:	o_val <= 16'b0101010000001000;
                14'h74c 	:	o_val <= 16'b0101010000010001;
                14'h74d 	:	o_val <= 16'b0101010000011011;
                14'h74e 	:	o_val <= 16'b0101010000100100;
                14'h74f 	:	o_val <= 16'b0101010000101110;
                14'h750 	:	o_val <= 16'b0101010000110111;
                14'h751 	:	o_val <= 16'b0101010001000001;
                14'h752 	:	o_val <= 16'b0101010001001010;
                14'h753 	:	o_val <= 16'b0101010001010100;
                14'h754 	:	o_val <= 16'b0101010001011101;
                14'h755 	:	o_val <= 16'b0101010001100111;
                14'h756 	:	o_val <= 16'b0101010001110000;
                14'h757 	:	o_val <= 16'b0101010001111001;
                14'h758 	:	o_val <= 16'b0101010010000011;
                14'h759 	:	o_val <= 16'b0101010010001100;
                14'h75a 	:	o_val <= 16'b0101010010010110;
                14'h75b 	:	o_val <= 16'b0101010010011111;
                14'h75c 	:	o_val <= 16'b0101010010101001;
                14'h75d 	:	o_val <= 16'b0101010010110010;
                14'h75e 	:	o_val <= 16'b0101010010111011;
                14'h75f 	:	o_val <= 16'b0101010011000101;
                14'h760 	:	o_val <= 16'b0101010011001110;
                14'h761 	:	o_val <= 16'b0101010011011000;
                14'h762 	:	o_val <= 16'b0101010011100001;
                14'h763 	:	o_val <= 16'b0101010011101010;
                14'h764 	:	o_val <= 16'b0101010011110100;
                14'h765 	:	o_val <= 16'b0101010011111101;
                14'h766 	:	o_val <= 16'b0101010100000111;
                14'h767 	:	o_val <= 16'b0101010100010000;
                14'h768 	:	o_val <= 16'b0101010100011001;
                14'h769 	:	o_val <= 16'b0101010100100011;
                14'h76a 	:	o_val <= 16'b0101010100101100;
                14'h76b 	:	o_val <= 16'b0101010100110110;
                14'h76c 	:	o_val <= 16'b0101010100111111;
                14'h76d 	:	o_val <= 16'b0101010101001000;
                14'h76e 	:	o_val <= 16'b0101010101010010;
                14'h76f 	:	o_val <= 16'b0101010101011011;
                14'h770 	:	o_val <= 16'b0101010101100100;
                14'h771 	:	o_val <= 16'b0101010101101110;
                14'h772 	:	o_val <= 16'b0101010101110111;
                14'h773 	:	o_val <= 16'b0101010110000001;
                14'h774 	:	o_val <= 16'b0101010110001010;
                14'h775 	:	o_val <= 16'b0101010110010011;
                14'h776 	:	o_val <= 16'b0101010110011101;
                14'h777 	:	o_val <= 16'b0101010110100110;
                14'h778 	:	o_val <= 16'b0101010110101111;
                14'h779 	:	o_val <= 16'b0101010110111001;
                14'h77a 	:	o_val <= 16'b0101010111000010;
                14'h77b 	:	o_val <= 16'b0101010111001011;
                14'h77c 	:	o_val <= 16'b0101010111010101;
                14'h77d 	:	o_val <= 16'b0101010111011110;
                14'h77e 	:	o_val <= 16'b0101010111100111;
                14'h77f 	:	o_val <= 16'b0101010111110000;
                14'h780 	:	o_val <= 16'b0101010111111010;
                14'h781 	:	o_val <= 16'b0101011000000011;
                14'h782 	:	o_val <= 16'b0101011000001100;
                14'h783 	:	o_val <= 16'b0101011000010110;
                14'h784 	:	o_val <= 16'b0101011000011111;
                14'h785 	:	o_val <= 16'b0101011000101000;
                14'h786 	:	o_val <= 16'b0101011000110010;
                14'h787 	:	o_val <= 16'b0101011000111011;
                14'h788 	:	o_val <= 16'b0101011001000100;
                14'h789 	:	o_val <= 16'b0101011001001101;
                14'h78a 	:	o_val <= 16'b0101011001010111;
                14'h78b 	:	o_val <= 16'b0101011001100000;
                14'h78c 	:	o_val <= 16'b0101011001101001;
                14'h78d 	:	o_val <= 16'b0101011001110011;
                14'h78e 	:	o_val <= 16'b0101011001111100;
                14'h78f 	:	o_val <= 16'b0101011010000101;
                14'h790 	:	o_val <= 16'b0101011010001110;
                14'h791 	:	o_val <= 16'b0101011010011000;
                14'h792 	:	o_val <= 16'b0101011010100001;
                14'h793 	:	o_val <= 16'b0101011010101010;
                14'h794 	:	o_val <= 16'b0101011010110011;
                14'h795 	:	o_val <= 16'b0101011010111101;
                14'h796 	:	o_val <= 16'b0101011011000110;
                14'h797 	:	o_val <= 16'b0101011011001111;
                14'h798 	:	o_val <= 16'b0101011011011000;
                14'h799 	:	o_val <= 16'b0101011011100010;
                14'h79a 	:	o_val <= 16'b0101011011101011;
                14'h79b 	:	o_val <= 16'b0101011011110100;
                14'h79c 	:	o_val <= 16'b0101011011111101;
                14'h79d 	:	o_val <= 16'b0101011100000110;
                14'h79e 	:	o_val <= 16'b0101011100010000;
                14'h79f 	:	o_val <= 16'b0101011100011001;
                14'h7a0 	:	o_val <= 16'b0101011100100010;
                14'h7a1 	:	o_val <= 16'b0101011100101011;
                14'h7a2 	:	o_val <= 16'b0101011100110100;
                14'h7a3 	:	o_val <= 16'b0101011100111110;
                14'h7a4 	:	o_val <= 16'b0101011101000111;
                14'h7a5 	:	o_val <= 16'b0101011101010000;
                14'h7a6 	:	o_val <= 16'b0101011101011001;
                14'h7a7 	:	o_val <= 16'b0101011101100010;
                14'h7a8 	:	o_val <= 16'b0101011101101100;
                14'h7a9 	:	o_val <= 16'b0101011101110101;
                14'h7aa 	:	o_val <= 16'b0101011101111110;
                14'h7ab 	:	o_val <= 16'b0101011110000111;
                14'h7ac 	:	o_val <= 16'b0101011110010000;
                14'h7ad 	:	o_val <= 16'b0101011110011001;
                14'h7ae 	:	o_val <= 16'b0101011110100011;
                14'h7af 	:	o_val <= 16'b0101011110101100;
                14'h7b0 	:	o_val <= 16'b0101011110110101;
                14'h7b1 	:	o_val <= 16'b0101011110111110;
                14'h7b2 	:	o_val <= 16'b0101011111000111;
                14'h7b3 	:	o_val <= 16'b0101011111010000;
                14'h7b4 	:	o_val <= 16'b0101011111011001;
                14'h7b5 	:	o_val <= 16'b0101011111100011;
                14'h7b6 	:	o_val <= 16'b0101011111101100;
                14'h7b7 	:	o_val <= 16'b0101011111110101;
                14'h7b8 	:	o_val <= 16'b0101011111111110;
                14'h7b9 	:	o_val <= 16'b0101100000000111;
                14'h7ba 	:	o_val <= 16'b0101100000010000;
                14'h7bb 	:	o_val <= 16'b0101100000011001;
                14'h7bc 	:	o_val <= 16'b0101100000100010;
                14'h7bd 	:	o_val <= 16'b0101100000101100;
                14'h7be 	:	o_val <= 16'b0101100000110101;
                14'h7bf 	:	o_val <= 16'b0101100000111110;
                14'h7c0 	:	o_val <= 16'b0101100001000111;
                14'h7c1 	:	o_val <= 16'b0101100001010000;
                14'h7c2 	:	o_val <= 16'b0101100001011001;
                14'h7c3 	:	o_val <= 16'b0101100001100010;
                14'h7c4 	:	o_val <= 16'b0101100001101011;
                14'h7c5 	:	o_val <= 16'b0101100001110100;
                14'h7c6 	:	o_val <= 16'b0101100001111101;
                14'h7c7 	:	o_val <= 16'b0101100010000111;
                14'h7c8 	:	o_val <= 16'b0101100010010000;
                14'h7c9 	:	o_val <= 16'b0101100010011001;
                14'h7ca 	:	o_val <= 16'b0101100010100010;
                14'h7cb 	:	o_val <= 16'b0101100010101011;
                14'h7cc 	:	o_val <= 16'b0101100010110100;
                14'h7cd 	:	o_val <= 16'b0101100010111101;
                14'h7ce 	:	o_val <= 16'b0101100011000110;
                14'h7cf 	:	o_val <= 16'b0101100011001111;
                14'h7d0 	:	o_val <= 16'b0101100011011000;
                14'h7d1 	:	o_val <= 16'b0101100011100001;
                14'h7d2 	:	o_val <= 16'b0101100011101010;
                14'h7d3 	:	o_val <= 16'b0101100011110011;
                14'h7d4 	:	o_val <= 16'b0101100011111100;
                14'h7d5 	:	o_val <= 16'b0101100100000101;
                14'h7d6 	:	o_val <= 16'b0101100100001110;
                14'h7d7 	:	o_val <= 16'b0101100100010111;
                14'h7d8 	:	o_val <= 16'b0101100100100000;
                14'h7d9 	:	o_val <= 16'b0101100100101001;
                14'h7da 	:	o_val <= 16'b0101100100110010;
                14'h7db 	:	o_val <= 16'b0101100100111011;
                14'h7dc 	:	o_val <= 16'b0101100101000100;
                14'h7dd 	:	o_val <= 16'b0101100101001101;
                14'h7de 	:	o_val <= 16'b0101100101010110;
                14'h7df 	:	o_val <= 16'b0101100101011111;
                14'h7e0 	:	o_val <= 16'b0101100101101000;
                14'h7e1 	:	o_val <= 16'b0101100101110001;
                14'h7e2 	:	o_val <= 16'b0101100101111010;
                14'h7e3 	:	o_val <= 16'b0101100110000011;
                14'h7e4 	:	o_val <= 16'b0101100110001100;
                14'h7e5 	:	o_val <= 16'b0101100110010101;
                14'h7e6 	:	o_val <= 16'b0101100110011110;
                14'h7e7 	:	o_val <= 16'b0101100110100111;
                14'h7e8 	:	o_val <= 16'b0101100110110000;
                14'h7e9 	:	o_val <= 16'b0101100110111001;
                14'h7ea 	:	o_val <= 16'b0101100111000010;
                14'h7eb 	:	o_val <= 16'b0101100111001011;
                14'h7ec 	:	o_val <= 16'b0101100111010100;
                14'h7ed 	:	o_val <= 16'b0101100111011101;
                14'h7ee 	:	o_val <= 16'b0101100111100110;
                14'h7ef 	:	o_val <= 16'b0101100111101111;
                14'h7f0 	:	o_val <= 16'b0101100111111000;
                14'h7f1 	:	o_val <= 16'b0101101000000001;
                14'h7f2 	:	o_val <= 16'b0101101000001010;
                14'h7f3 	:	o_val <= 16'b0101101000010011;
                14'h7f4 	:	o_val <= 16'b0101101000011100;
                14'h7f5 	:	o_val <= 16'b0101101000100100;
                14'h7f6 	:	o_val <= 16'b0101101000101101;
                14'h7f7 	:	o_val <= 16'b0101101000110110;
                14'h7f8 	:	o_val <= 16'b0101101000111111;
                14'h7f9 	:	o_val <= 16'b0101101001001000;
                14'h7fa 	:	o_val <= 16'b0101101001010001;
                14'h7fb 	:	o_val <= 16'b0101101001011010;
                14'h7fc 	:	o_val <= 16'b0101101001100011;
                14'h7fd 	:	o_val <= 16'b0101101001101100;
                14'h7fe 	:	o_val <= 16'b0101101001110101;
                14'h7ff 	:	o_val <= 16'b0101101001111110;
                14'h800 	:	o_val <= 16'b0101101010000110;
                14'h801 	:	o_val <= 16'b0101101010001111;
                14'h802 	:	o_val <= 16'b0101101010011000;
                14'h803 	:	o_val <= 16'b0101101010100001;
                14'h804 	:	o_val <= 16'b0101101010101010;
                14'h805 	:	o_val <= 16'b0101101010110011;
                14'h806 	:	o_val <= 16'b0101101010111100;
                14'h807 	:	o_val <= 16'b0101101011000101;
                14'h808 	:	o_val <= 16'b0101101011001101;
                14'h809 	:	o_val <= 16'b0101101011010110;
                14'h80a 	:	o_val <= 16'b0101101011011111;
                14'h80b 	:	o_val <= 16'b0101101011101000;
                14'h80c 	:	o_val <= 16'b0101101011110001;
                14'h80d 	:	o_val <= 16'b0101101011111010;
                14'h80e 	:	o_val <= 16'b0101101100000010;
                14'h80f 	:	o_val <= 16'b0101101100001011;
                14'h810 	:	o_val <= 16'b0101101100010100;
                14'h811 	:	o_val <= 16'b0101101100011101;
                14'h812 	:	o_val <= 16'b0101101100100110;
                14'h813 	:	o_val <= 16'b0101101100101111;
                14'h814 	:	o_val <= 16'b0101101100110111;
                14'h815 	:	o_val <= 16'b0101101101000000;
                14'h816 	:	o_val <= 16'b0101101101001001;
                14'h817 	:	o_val <= 16'b0101101101010010;
                14'h818 	:	o_val <= 16'b0101101101011011;
                14'h819 	:	o_val <= 16'b0101101101100011;
                14'h81a 	:	o_val <= 16'b0101101101101100;
                14'h81b 	:	o_val <= 16'b0101101101110101;
                14'h81c 	:	o_val <= 16'b0101101101111110;
                14'h81d 	:	o_val <= 16'b0101101110000111;
                14'h81e 	:	o_val <= 16'b0101101110001111;
                14'h81f 	:	o_val <= 16'b0101101110011000;
                14'h820 	:	o_val <= 16'b0101101110100001;
                14'h821 	:	o_val <= 16'b0101101110101010;
                14'h822 	:	o_val <= 16'b0101101110110010;
                14'h823 	:	o_val <= 16'b0101101110111011;
                14'h824 	:	o_val <= 16'b0101101111000100;
                14'h825 	:	o_val <= 16'b0101101111001101;
                14'h826 	:	o_val <= 16'b0101101111010110;
                14'h827 	:	o_val <= 16'b0101101111011110;
                14'h828 	:	o_val <= 16'b0101101111100111;
                14'h829 	:	o_val <= 16'b0101101111110000;
                14'h82a 	:	o_val <= 16'b0101101111111001;
                14'h82b 	:	o_val <= 16'b0101110000000001;
                14'h82c 	:	o_val <= 16'b0101110000001010;
                14'h82d 	:	o_val <= 16'b0101110000010011;
                14'h82e 	:	o_val <= 16'b0101110000011011;
                14'h82f 	:	o_val <= 16'b0101110000100100;
                14'h830 	:	o_val <= 16'b0101110000101101;
                14'h831 	:	o_val <= 16'b0101110000110110;
                14'h832 	:	o_val <= 16'b0101110000111110;
                14'h833 	:	o_val <= 16'b0101110001000111;
                14'h834 	:	o_val <= 16'b0101110001010000;
                14'h835 	:	o_val <= 16'b0101110001011000;
                14'h836 	:	o_val <= 16'b0101110001100001;
                14'h837 	:	o_val <= 16'b0101110001101010;
                14'h838 	:	o_val <= 16'b0101110001110011;
                14'h839 	:	o_val <= 16'b0101110001111011;
                14'h83a 	:	o_val <= 16'b0101110010000100;
                14'h83b 	:	o_val <= 16'b0101110010001101;
                14'h83c 	:	o_val <= 16'b0101110010010101;
                14'h83d 	:	o_val <= 16'b0101110010011110;
                14'h83e 	:	o_val <= 16'b0101110010100111;
                14'h83f 	:	o_val <= 16'b0101110010101111;
                14'h840 	:	o_val <= 16'b0101110010111000;
                14'h841 	:	o_val <= 16'b0101110011000001;
                14'h842 	:	o_val <= 16'b0101110011001001;
                14'h843 	:	o_val <= 16'b0101110011010010;
                14'h844 	:	o_val <= 16'b0101110011011011;
                14'h845 	:	o_val <= 16'b0101110011100011;
                14'h846 	:	o_val <= 16'b0101110011101100;
                14'h847 	:	o_val <= 16'b0101110011110101;
                14'h848 	:	o_val <= 16'b0101110011111101;
                14'h849 	:	o_val <= 16'b0101110100000110;
                14'h84a 	:	o_val <= 16'b0101110100001110;
                14'h84b 	:	o_val <= 16'b0101110100010111;
                14'h84c 	:	o_val <= 16'b0101110100100000;
                14'h84d 	:	o_val <= 16'b0101110100101000;
                14'h84e 	:	o_val <= 16'b0101110100110001;
                14'h84f 	:	o_val <= 16'b0101110100111010;
                14'h850 	:	o_val <= 16'b0101110101000010;
                14'h851 	:	o_val <= 16'b0101110101001011;
                14'h852 	:	o_val <= 16'b0101110101010011;
                14'h853 	:	o_val <= 16'b0101110101011100;
                14'h854 	:	o_val <= 16'b0101110101100101;
                14'h855 	:	o_val <= 16'b0101110101101101;
                14'h856 	:	o_val <= 16'b0101110101110110;
                14'h857 	:	o_val <= 16'b0101110101111110;
                14'h858 	:	o_val <= 16'b0101110110000111;
                14'h859 	:	o_val <= 16'b0101110110001111;
                14'h85a 	:	o_val <= 16'b0101110110011000;
                14'h85b 	:	o_val <= 16'b0101110110100001;
                14'h85c 	:	o_val <= 16'b0101110110101001;
                14'h85d 	:	o_val <= 16'b0101110110110010;
                14'h85e 	:	o_val <= 16'b0101110110111010;
                14'h85f 	:	o_val <= 16'b0101110111000011;
                14'h860 	:	o_val <= 16'b0101110111001011;
                14'h861 	:	o_val <= 16'b0101110111010100;
                14'h862 	:	o_val <= 16'b0101110111011100;
                14'h863 	:	o_val <= 16'b0101110111100101;
                14'h864 	:	o_val <= 16'b0101110111101110;
                14'h865 	:	o_val <= 16'b0101110111110110;
                14'h866 	:	o_val <= 16'b0101110111111111;
                14'h867 	:	o_val <= 16'b0101111000000111;
                14'h868 	:	o_val <= 16'b0101111000010000;
                14'h869 	:	o_val <= 16'b0101111000011000;
                14'h86a 	:	o_val <= 16'b0101111000100001;
                14'h86b 	:	o_val <= 16'b0101111000101001;
                14'h86c 	:	o_val <= 16'b0101111000110010;
                14'h86d 	:	o_val <= 16'b0101111000111010;
                14'h86e 	:	o_val <= 16'b0101111001000011;
                14'h86f 	:	o_val <= 16'b0101111001001011;
                14'h870 	:	o_val <= 16'b0101111001010100;
                14'h871 	:	o_val <= 16'b0101111001011100;
                14'h872 	:	o_val <= 16'b0101111001100101;
                14'h873 	:	o_val <= 16'b0101111001101101;
                14'h874 	:	o_val <= 16'b0101111001110110;
                14'h875 	:	o_val <= 16'b0101111001111110;
                14'h876 	:	o_val <= 16'b0101111010000111;
                14'h877 	:	o_val <= 16'b0101111010001111;
                14'h878 	:	o_val <= 16'b0101111010011000;
                14'h879 	:	o_val <= 16'b0101111010100000;
                14'h87a 	:	o_val <= 16'b0101111010101001;
                14'h87b 	:	o_val <= 16'b0101111010110001;
                14'h87c 	:	o_val <= 16'b0101111010111001;
                14'h87d 	:	o_val <= 16'b0101111011000010;
                14'h87e 	:	o_val <= 16'b0101111011001010;
                14'h87f 	:	o_val <= 16'b0101111011010011;
                14'h880 	:	o_val <= 16'b0101111011011011;
                14'h881 	:	o_val <= 16'b0101111011100100;
                14'h882 	:	o_val <= 16'b0101111011101100;
                14'h883 	:	o_val <= 16'b0101111011110101;
                14'h884 	:	o_val <= 16'b0101111011111101;
                14'h885 	:	o_val <= 16'b0101111100000101;
                14'h886 	:	o_val <= 16'b0101111100001110;
                14'h887 	:	o_val <= 16'b0101111100010110;
                14'h888 	:	o_val <= 16'b0101111100011111;
                14'h889 	:	o_val <= 16'b0101111100100111;
                14'h88a 	:	o_val <= 16'b0101111100101111;
                14'h88b 	:	o_val <= 16'b0101111100111000;
                14'h88c 	:	o_val <= 16'b0101111101000000;
                14'h88d 	:	o_val <= 16'b0101111101001001;
                14'h88e 	:	o_val <= 16'b0101111101010001;
                14'h88f 	:	o_val <= 16'b0101111101011001;
                14'h890 	:	o_val <= 16'b0101111101100010;
                14'h891 	:	o_val <= 16'b0101111101101010;
                14'h892 	:	o_val <= 16'b0101111101110010;
                14'h893 	:	o_val <= 16'b0101111101111011;
                14'h894 	:	o_val <= 16'b0101111110000011;
                14'h895 	:	o_val <= 16'b0101111110001100;
                14'h896 	:	o_val <= 16'b0101111110010100;
                14'h897 	:	o_val <= 16'b0101111110011100;
                14'h898 	:	o_val <= 16'b0101111110100101;
                14'h899 	:	o_val <= 16'b0101111110101101;
                14'h89a 	:	o_val <= 16'b0101111110110101;
                14'h89b 	:	o_val <= 16'b0101111110111110;
                14'h89c 	:	o_val <= 16'b0101111111000110;
                14'h89d 	:	o_val <= 16'b0101111111001110;
                14'h89e 	:	o_val <= 16'b0101111111010111;
                14'h89f 	:	o_val <= 16'b0101111111011111;
                14'h8a0 	:	o_val <= 16'b0101111111100111;
                14'h8a1 	:	o_val <= 16'b0101111111110000;
                14'h8a2 	:	o_val <= 16'b0101111111111000;
                14'h8a3 	:	o_val <= 16'b0110000000000000;
                14'h8a4 	:	o_val <= 16'b0110000000001001;
                14'h8a5 	:	o_val <= 16'b0110000000010001;
                14'h8a6 	:	o_val <= 16'b0110000000011001;
                14'h8a7 	:	o_val <= 16'b0110000000100010;
                14'h8a8 	:	o_val <= 16'b0110000000101010;
                14'h8a9 	:	o_val <= 16'b0110000000110010;
                14'h8aa 	:	o_val <= 16'b0110000000111010;
                14'h8ab 	:	o_val <= 16'b0110000001000011;
                14'h8ac 	:	o_val <= 16'b0110000001001011;
                14'h8ad 	:	o_val <= 16'b0110000001010011;
                14'h8ae 	:	o_val <= 16'b0110000001011100;
                14'h8af 	:	o_val <= 16'b0110000001100100;
                14'h8b0 	:	o_val <= 16'b0110000001101100;
                14'h8b1 	:	o_val <= 16'b0110000001110100;
                14'h8b2 	:	o_val <= 16'b0110000001111101;
                14'h8b3 	:	o_val <= 16'b0110000010000101;
                14'h8b4 	:	o_val <= 16'b0110000010001101;
                14'h8b5 	:	o_val <= 16'b0110000010010101;
                14'h8b6 	:	o_val <= 16'b0110000010011110;
                14'h8b7 	:	o_val <= 16'b0110000010100110;
                14'h8b8 	:	o_val <= 16'b0110000010101110;
                14'h8b9 	:	o_val <= 16'b0110000010110110;
                14'h8ba 	:	o_val <= 16'b0110000010111111;
                14'h8bb 	:	o_val <= 16'b0110000011000111;
                14'h8bc 	:	o_val <= 16'b0110000011001111;
                14'h8bd 	:	o_val <= 16'b0110000011010111;
                14'h8be 	:	o_val <= 16'b0110000011011111;
                14'h8bf 	:	o_val <= 16'b0110000011101000;
                14'h8c0 	:	o_val <= 16'b0110000011110000;
                14'h8c1 	:	o_val <= 16'b0110000011111000;
                14'h8c2 	:	o_val <= 16'b0110000100000000;
                14'h8c3 	:	o_val <= 16'b0110000100001000;
                14'h8c4 	:	o_val <= 16'b0110000100010001;
                14'h8c5 	:	o_val <= 16'b0110000100011001;
                14'h8c6 	:	o_val <= 16'b0110000100100001;
                14'h8c7 	:	o_val <= 16'b0110000100101001;
                14'h8c8 	:	o_val <= 16'b0110000100110001;
                14'h8c9 	:	o_val <= 16'b0110000100111010;
                14'h8ca 	:	o_val <= 16'b0110000101000010;
                14'h8cb 	:	o_val <= 16'b0110000101001010;
                14'h8cc 	:	o_val <= 16'b0110000101010010;
                14'h8cd 	:	o_val <= 16'b0110000101011010;
                14'h8ce 	:	o_val <= 16'b0110000101100010;
                14'h8cf 	:	o_val <= 16'b0110000101101011;
                14'h8d0 	:	o_val <= 16'b0110000101110011;
                14'h8d1 	:	o_val <= 16'b0110000101111011;
                14'h8d2 	:	o_val <= 16'b0110000110000011;
                14'h8d3 	:	o_val <= 16'b0110000110001011;
                14'h8d4 	:	o_val <= 16'b0110000110010011;
                14'h8d5 	:	o_val <= 16'b0110000110011011;
                14'h8d6 	:	o_val <= 16'b0110000110100011;
                14'h8d7 	:	o_val <= 16'b0110000110101100;
                14'h8d8 	:	o_val <= 16'b0110000110110100;
                14'h8d9 	:	o_val <= 16'b0110000110111100;
                14'h8da 	:	o_val <= 16'b0110000111000100;
                14'h8db 	:	o_val <= 16'b0110000111001100;
                14'h8dc 	:	o_val <= 16'b0110000111010100;
                14'h8dd 	:	o_val <= 16'b0110000111011100;
                14'h8de 	:	o_val <= 16'b0110000111100100;
                14'h8df 	:	o_val <= 16'b0110000111101100;
                14'h8e0 	:	o_val <= 16'b0110000111110101;
                14'h8e1 	:	o_val <= 16'b0110000111111101;
                14'h8e2 	:	o_val <= 16'b0110001000000101;
                14'h8e3 	:	o_val <= 16'b0110001000001101;
                14'h8e4 	:	o_val <= 16'b0110001000010101;
                14'h8e5 	:	o_val <= 16'b0110001000011101;
                14'h8e6 	:	o_val <= 16'b0110001000100101;
                14'h8e7 	:	o_val <= 16'b0110001000101101;
                14'h8e8 	:	o_val <= 16'b0110001000110101;
                14'h8e9 	:	o_val <= 16'b0110001000111101;
                14'h8ea 	:	o_val <= 16'b0110001001000101;
                14'h8eb 	:	o_val <= 16'b0110001001001101;
                14'h8ec 	:	o_val <= 16'b0110001001010101;
                14'h8ed 	:	o_val <= 16'b0110001001011101;
                14'h8ee 	:	o_val <= 16'b0110001001100101;
                14'h8ef 	:	o_val <= 16'b0110001001101101;
                14'h8f0 	:	o_val <= 16'b0110001001110101;
                14'h8f1 	:	o_val <= 16'b0110001001111110;
                14'h8f2 	:	o_val <= 16'b0110001010000110;
                14'h8f3 	:	o_val <= 16'b0110001010001110;
                14'h8f4 	:	o_val <= 16'b0110001010010110;
                14'h8f5 	:	o_val <= 16'b0110001010011110;
                14'h8f6 	:	o_val <= 16'b0110001010100110;
                14'h8f7 	:	o_val <= 16'b0110001010101110;
                14'h8f8 	:	o_val <= 16'b0110001010110110;
                14'h8f9 	:	o_val <= 16'b0110001010111110;
                14'h8fa 	:	o_val <= 16'b0110001011000110;
                14'h8fb 	:	o_val <= 16'b0110001011001110;
                14'h8fc 	:	o_val <= 16'b0110001011010110;
                14'h8fd 	:	o_val <= 16'b0110001011011110;
                14'h8fe 	:	o_val <= 16'b0110001011100110;
                14'h8ff 	:	o_val <= 16'b0110001011101110;
                14'h900 	:	o_val <= 16'b0110001011110101;
                14'h901 	:	o_val <= 16'b0110001011111101;
                14'h902 	:	o_val <= 16'b0110001100000101;
                14'h903 	:	o_val <= 16'b0110001100001101;
                14'h904 	:	o_val <= 16'b0110001100010101;
                14'h905 	:	o_val <= 16'b0110001100011101;
                14'h906 	:	o_val <= 16'b0110001100100101;
                14'h907 	:	o_val <= 16'b0110001100101101;
                14'h908 	:	o_val <= 16'b0110001100110101;
                14'h909 	:	o_val <= 16'b0110001100111101;
                14'h90a 	:	o_val <= 16'b0110001101000101;
                14'h90b 	:	o_val <= 16'b0110001101001101;
                14'h90c 	:	o_val <= 16'b0110001101010101;
                14'h90d 	:	o_val <= 16'b0110001101011101;
                14'h90e 	:	o_val <= 16'b0110001101100101;
                14'h90f 	:	o_val <= 16'b0110001101101101;
                14'h910 	:	o_val <= 16'b0110001101110101;
                14'h911 	:	o_val <= 16'b0110001101111100;
                14'h912 	:	o_val <= 16'b0110001110000100;
                14'h913 	:	o_val <= 16'b0110001110001100;
                14'h914 	:	o_val <= 16'b0110001110010100;
                14'h915 	:	o_val <= 16'b0110001110011100;
                14'h916 	:	o_val <= 16'b0110001110100100;
                14'h917 	:	o_val <= 16'b0110001110101100;
                14'h918 	:	o_val <= 16'b0110001110110100;
                14'h919 	:	o_val <= 16'b0110001110111100;
                14'h91a 	:	o_val <= 16'b0110001111000011;
                14'h91b 	:	o_val <= 16'b0110001111001011;
                14'h91c 	:	o_val <= 16'b0110001111010011;
                14'h91d 	:	o_val <= 16'b0110001111011011;
                14'h91e 	:	o_val <= 16'b0110001111100011;
                14'h91f 	:	o_val <= 16'b0110001111101011;
                14'h920 	:	o_val <= 16'b0110001111110011;
                14'h921 	:	o_val <= 16'b0110001111111010;
                14'h922 	:	o_val <= 16'b0110010000000010;
                14'h923 	:	o_val <= 16'b0110010000001010;
                14'h924 	:	o_val <= 16'b0110010000010010;
                14'h925 	:	o_val <= 16'b0110010000011010;
                14'h926 	:	o_val <= 16'b0110010000100010;
                14'h927 	:	o_val <= 16'b0110010000101001;
                14'h928 	:	o_val <= 16'b0110010000110001;
                14'h929 	:	o_val <= 16'b0110010000111001;
                14'h92a 	:	o_val <= 16'b0110010001000001;
                14'h92b 	:	o_val <= 16'b0110010001001001;
                14'h92c 	:	o_val <= 16'b0110010001010001;
                14'h92d 	:	o_val <= 16'b0110010001011000;
                14'h92e 	:	o_val <= 16'b0110010001100000;
                14'h92f 	:	o_val <= 16'b0110010001101000;
                14'h930 	:	o_val <= 16'b0110010001110000;
                14'h931 	:	o_val <= 16'b0110010001111000;
                14'h932 	:	o_val <= 16'b0110010001111111;
                14'h933 	:	o_val <= 16'b0110010010000111;
                14'h934 	:	o_val <= 16'b0110010010001111;
                14'h935 	:	o_val <= 16'b0110010010010111;
                14'h936 	:	o_val <= 16'b0110010010011110;
                14'h937 	:	o_val <= 16'b0110010010100110;
                14'h938 	:	o_val <= 16'b0110010010101110;
                14'h939 	:	o_val <= 16'b0110010010110110;
                14'h93a 	:	o_val <= 16'b0110010010111101;
                14'h93b 	:	o_val <= 16'b0110010011000101;
                14'h93c 	:	o_val <= 16'b0110010011001101;
                14'h93d 	:	o_val <= 16'b0110010011010101;
                14'h93e 	:	o_val <= 16'b0110010011011100;
                14'h93f 	:	o_val <= 16'b0110010011100100;
                14'h940 	:	o_val <= 16'b0110010011101100;
                14'h941 	:	o_val <= 16'b0110010011110100;
                14'h942 	:	o_val <= 16'b0110010011111011;
                14'h943 	:	o_val <= 16'b0110010100000011;
                14'h944 	:	o_val <= 16'b0110010100001011;
                14'h945 	:	o_val <= 16'b0110010100010011;
                14'h946 	:	o_val <= 16'b0110010100011010;
                14'h947 	:	o_val <= 16'b0110010100100010;
                14'h948 	:	o_val <= 16'b0110010100101010;
                14'h949 	:	o_val <= 16'b0110010100110001;
                14'h94a 	:	o_val <= 16'b0110010100111001;
                14'h94b 	:	o_val <= 16'b0110010101000001;
                14'h94c 	:	o_val <= 16'b0110010101001000;
                14'h94d 	:	o_val <= 16'b0110010101010000;
                14'h94e 	:	o_val <= 16'b0110010101011000;
                14'h94f 	:	o_val <= 16'b0110010101011111;
                14'h950 	:	o_val <= 16'b0110010101100111;
                14'h951 	:	o_val <= 16'b0110010101101111;
                14'h952 	:	o_val <= 16'b0110010101110110;
                14'h953 	:	o_val <= 16'b0110010101111110;
                14'h954 	:	o_val <= 16'b0110010110000110;
                14'h955 	:	o_val <= 16'b0110010110001101;
                14'h956 	:	o_val <= 16'b0110010110010101;
                14'h957 	:	o_val <= 16'b0110010110011101;
                14'h958 	:	o_val <= 16'b0110010110100100;
                14'h959 	:	o_val <= 16'b0110010110101100;
                14'h95a 	:	o_val <= 16'b0110010110110100;
                14'h95b 	:	o_val <= 16'b0110010110111011;
                14'h95c 	:	o_val <= 16'b0110010111000011;
                14'h95d 	:	o_val <= 16'b0110010111001010;
                14'h95e 	:	o_val <= 16'b0110010111010010;
                14'h95f 	:	o_val <= 16'b0110010111011010;
                14'h960 	:	o_val <= 16'b0110010111100001;
                14'h961 	:	o_val <= 16'b0110010111101001;
                14'h962 	:	o_val <= 16'b0110010111110000;
                14'h963 	:	o_val <= 16'b0110010111111000;
                14'h964 	:	o_val <= 16'b0110011000000000;
                14'h965 	:	o_val <= 16'b0110011000000111;
                14'h966 	:	o_val <= 16'b0110011000001111;
                14'h967 	:	o_val <= 16'b0110011000010110;
                14'h968 	:	o_val <= 16'b0110011000011110;
                14'h969 	:	o_val <= 16'b0110011000100110;
                14'h96a 	:	o_val <= 16'b0110011000101101;
                14'h96b 	:	o_val <= 16'b0110011000110101;
                14'h96c 	:	o_val <= 16'b0110011000111100;
                14'h96d 	:	o_val <= 16'b0110011001000100;
                14'h96e 	:	o_val <= 16'b0110011001001011;
                14'h96f 	:	o_val <= 16'b0110011001010011;
                14'h970 	:	o_val <= 16'b0110011001011011;
                14'h971 	:	o_val <= 16'b0110011001100010;
                14'h972 	:	o_val <= 16'b0110011001101010;
                14'h973 	:	o_val <= 16'b0110011001110001;
                14'h974 	:	o_val <= 16'b0110011001111001;
                14'h975 	:	o_val <= 16'b0110011010000000;
                14'h976 	:	o_val <= 16'b0110011010001000;
                14'h977 	:	o_val <= 16'b0110011010001111;
                14'h978 	:	o_val <= 16'b0110011010010111;
                14'h979 	:	o_val <= 16'b0110011010011110;
                14'h97a 	:	o_val <= 16'b0110011010100110;
                14'h97b 	:	o_val <= 16'b0110011010101101;
                14'h97c 	:	o_val <= 16'b0110011010110101;
                14'h97d 	:	o_val <= 16'b0110011010111100;
                14'h97e 	:	o_val <= 16'b0110011011000100;
                14'h97f 	:	o_val <= 16'b0110011011001011;
                14'h980 	:	o_val <= 16'b0110011011010011;
                14'h981 	:	o_val <= 16'b0110011011011010;
                14'h982 	:	o_val <= 16'b0110011011100010;
                14'h983 	:	o_val <= 16'b0110011011101001;
                14'h984 	:	o_val <= 16'b0110011011110001;
                14'h985 	:	o_val <= 16'b0110011011111000;
                14'h986 	:	o_val <= 16'b0110011100000000;
                14'h987 	:	o_val <= 16'b0110011100000111;
                14'h988 	:	o_val <= 16'b0110011100001110;
                14'h989 	:	o_val <= 16'b0110011100010110;
                14'h98a 	:	o_val <= 16'b0110011100011101;
                14'h98b 	:	o_val <= 16'b0110011100100101;
                14'h98c 	:	o_val <= 16'b0110011100101100;
                14'h98d 	:	o_val <= 16'b0110011100110100;
                14'h98e 	:	o_val <= 16'b0110011100111011;
                14'h98f 	:	o_val <= 16'b0110011101000011;
                14'h990 	:	o_val <= 16'b0110011101001010;
                14'h991 	:	o_val <= 16'b0110011101010001;
                14'h992 	:	o_val <= 16'b0110011101011001;
                14'h993 	:	o_val <= 16'b0110011101100000;
                14'h994 	:	o_val <= 16'b0110011101101000;
                14'h995 	:	o_val <= 16'b0110011101101111;
                14'h996 	:	o_val <= 16'b0110011101110110;
                14'h997 	:	o_val <= 16'b0110011101111110;
                14'h998 	:	o_val <= 16'b0110011110000101;
                14'h999 	:	o_val <= 16'b0110011110001101;
                14'h99a 	:	o_val <= 16'b0110011110010100;
                14'h99b 	:	o_val <= 16'b0110011110011011;
                14'h99c 	:	o_val <= 16'b0110011110100011;
                14'h99d 	:	o_val <= 16'b0110011110101010;
                14'h99e 	:	o_val <= 16'b0110011110110010;
                14'h99f 	:	o_val <= 16'b0110011110111001;
                14'h9a0 	:	o_val <= 16'b0110011111000000;
                14'h9a1 	:	o_val <= 16'b0110011111001000;
                14'h9a2 	:	o_val <= 16'b0110011111001111;
                14'h9a3 	:	o_val <= 16'b0110011111010110;
                14'h9a4 	:	o_val <= 16'b0110011111011110;
                14'h9a5 	:	o_val <= 16'b0110011111100101;
                14'h9a6 	:	o_val <= 16'b0110011111101100;
                14'h9a7 	:	o_val <= 16'b0110011111110100;
                14'h9a8 	:	o_val <= 16'b0110011111111011;
                14'h9a9 	:	o_val <= 16'b0110100000000010;
                14'h9aa 	:	o_val <= 16'b0110100000001010;
                14'h9ab 	:	o_val <= 16'b0110100000010001;
                14'h9ac 	:	o_val <= 16'b0110100000011000;
                14'h9ad 	:	o_val <= 16'b0110100000100000;
                14'h9ae 	:	o_val <= 16'b0110100000100111;
                14'h9af 	:	o_val <= 16'b0110100000101110;
                14'h9b0 	:	o_val <= 16'b0110100000110101;
                14'h9b1 	:	o_val <= 16'b0110100000111101;
                14'h9b2 	:	o_val <= 16'b0110100001000100;
                14'h9b3 	:	o_val <= 16'b0110100001001011;
                14'h9b4 	:	o_val <= 16'b0110100001010011;
                14'h9b5 	:	o_val <= 16'b0110100001011010;
                14'h9b6 	:	o_val <= 16'b0110100001100001;
                14'h9b7 	:	o_val <= 16'b0110100001101000;
                14'h9b8 	:	o_val <= 16'b0110100001110000;
                14'h9b9 	:	o_val <= 16'b0110100001110111;
                14'h9ba 	:	o_val <= 16'b0110100001111110;
                14'h9bb 	:	o_val <= 16'b0110100010000110;
                14'h9bc 	:	o_val <= 16'b0110100010001101;
                14'h9bd 	:	o_val <= 16'b0110100010010100;
                14'h9be 	:	o_val <= 16'b0110100010011011;
                14'h9bf 	:	o_val <= 16'b0110100010100011;
                14'h9c0 	:	o_val <= 16'b0110100010101010;
                14'h9c1 	:	o_val <= 16'b0110100010110001;
                14'h9c2 	:	o_val <= 16'b0110100010111000;
                14'h9c3 	:	o_val <= 16'b0110100010111111;
                14'h9c4 	:	o_val <= 16'b0110100011000111;
                14'h9c5 	:	o_val <= 16'b0110100011001110;
                14'h9c6 	:	o_val <= 16'b0110100011010101;
                14'h9c7 	:	o_val <= 16'b0110100011011100;
                14'h9c8 	:	o_val <= 16'b0110100011100011;
                14'h9c9 	:	o_val <= 16'b0110100011101011;
                14'h9ca 	:	o_val <= 16'b0110100011110010;
                14'h9cb 	:	o_val <= 16'b0110100011111001;
                14'h9cc 	:	o_val <= 16'b0110100100000000;
                14'h9cd 	:	o_val <= 16'b0110100100000111;
                14'h9ce 	:	o_val <= 16'b0110100100001111;
                14'h9cf 	:	o_val <= 16'b0110100100010110;
                14'h9d0 	:	o_val <= 16'b0110100100011101;
                14'h9d1 	:	o_val <= 16'b0110100100100100;
                14'h9d2 	:	o_val <= 16'b0110100100101011;
                14'h9d3 	:	o_val <= 16'b0110100100110010;
                14'h9d4 	:	o_val <= 16'b0110100100111010;
                14'h9d5 	:	o_val <= 16'b0110100101000001;
                14'h9d6 	:	o_val <= 16'b0110100101001000;
                14'h9d7 	:	o_val <= 16'b0110100101001111;
                14'h9d8 	:	o_val <= 16'b0110100101010110;
                14'h9d9 	:	o_val <= 16'b0110100101011101;
                14'h9da 	:	o_val <= 16'b0110100101100100;
                14'h9db 	:	o_val <= 16'b0110100101101100;
                14'h9dc 	:	o_val <= 16'b0110100101110011;
                14'h9dd 	:	o_val <= 16'b0110100101111010;
                14'h9de 	:	o_val <= 16'b0110100110000001;
                14'h9df 	:	o_val <= 16'b0110100110001000;
                14'h9e0 	:	o_val <= 16'b0110100110001111;
                14'h9e1 	:	o_val <= 16'b0110100110010110;
                14'h9e2 	:	o_val <= 16'b0110100110011101;
                14'h9e3 	:	o_val <= 16'b0110100110100101;
                14'h9e4 	:	o_val <= 16'b0110100110101100;
                14'h9e5 	:	o_val <= 16'b0110100110110011;
                14'h9e6 	:	o_val <= 16'b0110100110111010;
                14'h9e7 	:	o_val <= 16'b0110100111000001;
                14'h9e8 	:	o_val <= 16'b0110100111001000;
                14'h9e9 	:	o_val <= 16'b0110100111001111;
                14'h9ea 	:	o_val <= 16'b0110100111010110;
                14'h9eb 	:	o_val <= 16'b0110100111011101;
                14'h9ec 	:	o_val <= 16'b0110100111100100;
                14'h9ed 	:	o_val <= 16'b0110100111101011;
                14'h9ee 	:	o_val <= 16'b0110100111110010;
                14'h9ef 	:	o_val <= 16'b0110100111111001;
                14'h9f0 	:	o_val <= 16'b0110101000000000;
                14'h9f1 	:	o_val <= 16'b0110101000000111;
                14'h9f2 	:	o_val <= 16'b0110101000001110;
                14'h9f3 	:	o_val <= 16'b0110101000010110;
                14'h9f4 	:	o_val <= 16'b0110101000011101;
                14'h9f5 	:	o_val <= 16'b0110101000100100;
                14'h9f6 	:	o_val <= 16'b0110101000101011;
                14'h9f7 	:	o_val <= 16'b0110101000110010;
                14'h9f8 	:	o_val <= 16'b0110101000111001;
                14'h9f9 	:	o_val <= 16'b0110101001000000;
                14'h9fa 	:	o_val <= 16'b0110101001000111;
                14'h9fb 	:	o_val <= 16'b0110101001001110;
                14'h9fc 	:	o_val <= 16'b0110101001010101;
                14'h9fd 	:	o_val <= 16'b0110101001011100;
                14'h9fe 	:	o_val <= 16'b0110101001100011;
                14'h9ff 	:	o_val <= 16'b0110101001101010;
                14'ha00 	:	o_val <= 16'b0110101001110001;
                14'ha01 	:	o_val <= 16'b0110101001111000;
                14'ha02 	:	o_val <= 16'b0110101001111111;
                14'ha03 	:	o_val <= 16'b0110101010000110;
                14'ha04 	:	o_val <= 16'b0110101010001100;
                14'ha05 	:	o_val <= 16'b0110101010010011;
                14'ha06 	:	o_val <= 16'b0110101010011010;
                14'ha07 	:	o_val <= 16'b0110101010100001;
                14'ha08 	:	o_val <= 16'b0110101010101000;
                14'ha09 	:	o_val <= 16'b0110101010101111;
                14'ha0a 	:	o_val <= 16'b0110101010110110;
                14'ha0b 	:	o_val <= 16'b0110101010111101;
                14'ha0c 	:	o_val <= 16'b0110101011000100;
                14'ha0d 	:	o_val <= 16'b0110101011001011;
                14'ha0e 	:	o_val <= 16'b0110101011010010;
                14'ha0f 	:	o_val <= 16'b0110101011011001;
                14'ha10 	:	o_val <= 16'b0110101011100000;
                14'ha11 	:	o_val <= 16'b0110101011100111;
                14'ha12 	:	o_val <= 16'b0110101011101110;
                14'ha13 	:	o_val <= 16'b0110101011110100;
                14'ha14 	:	o_val <= 16'b0110101011111011;
                14'ha15 	:	o_val <= 16'b0110101100000010;
                14'ha16 	:	o_val <= 16'b0110101100001001;
                14'ha17 	:	o_val <= 16'b0110101100010000;
                14'ha18 	:	o_val <= 16'b0110101100010111;
                14'ha19 	:	o_val <= 16'b0110101100011110;
                14'ha1a 	:	o_val <= 16'b0110101100100101;
                14'ha1b 	:	o_val <= 16'b0110101100101100;
                14'ha1c 	:	o_val <= 16'b0110101100110010;
                14'ha1d 	:	o_val <= 16'b0110101100111001;
                14'ha1e 	:	o_val <= 16'b0110101101000000;
                14'ha1f 	:	o_val <= 16'b0110101101000111;
                14'ha20 	:	o_val <= 16'b0110101101001110;
                14'ha21 	:	o_val <= 16'b0110101101010101;
                14'ha22 	:	o_val <= 16'b0110101101011100;
                14'ha23 	:	o_val <= 16'b0110101101100010;
                14'ha24 	:	o_val <= 16'b0110101101101001;
                14'ha25 	:	o_val <= 16'b0110101101110000;
                14'ha26 	:	o_val <= 16'b0110101101110111;
                14'ha27 	:	o_val <= 16'b0110101101111110;
                14'ha28 	:	o_val <= 16'b0110101110000101;
                14'ha29 	:	o_val <= 16'b0110101110001011;
                14'ha2a 	:	o_val <= 16'b0110101110010010;
                14'ha2b 	:	o_val <= 16'b0110101110011001;
                14'ha2c 	:	o_val <= 16'b0110101110100000;
                14'ha2d 	:	o_val <= 16'b0110101110100111;
                14'ha2e 	:	o_val <= 16'b0110101110101101;
                14'ha2f 	:	o_val <= 16'b0110101110110100;
                14'ha30 	:	o_val <= 16'b0110101110111011;
                14'ha31 	:	o_val <= 16'b0110101111000010;
                14'ha32 	:	o_val <= 16'b0110101111001001;
                14'ha33 	:	o_val <= 16'b0110101111001111;
                14'ha34 	:	o_val <= 16'b0110101111010110;
                14'ha35 	:	o_val <= 16'b0110101111011101;
                14'ha36 	:	o_val <= 16'b0110101111100100;
                14'ha37 	:	o_val <= 16'b0110101111101010;
                14'ha38 	:	o_val <= 16'b0110101111110001;
                14'ha39 	:	o_val <= 16'b0110101111111000;
                14'ha3a 	:	o_val <= 16'b0110101111111111;
                14'ha3b 	:	o_val <= 16'b0110110000000101;
                14'ha3c 	:	o_val <= 16'b0110110000001100;
                14'ha3d 	:	o_val <= 16'b0110110000010011;
                14'ha3e 	:	o_val <= 16'b0110110000011010;
                14'ha3f 	:	o_val <= 16'b0110110000100000;
                14'ha40 	:	o_val <= 16'b0110110000100111;
                14'ha41 	:	o_val <= 16'b0110110000101110;
                14'ha42 	:	o_val <= 16'b0110110000110100;
                14'ha43 	:	o_val <= 16'b0110110000111011;
                14'ha44 	:	o_val <= 16'b0110110001000010;
                14'ha45 	:	o_val <= 16'b0110110001001001;
                14'ha46 	:	o_val <= 16'b0110110001001111;
                14'ha47 	:	o_val <= 16'b0110110001010110;
                14'ha48 	:	o_val <= 16'b0110110001011101;
                14'ha49 	:	o_val <= 16'b0110110001100011;
                14'ha4a 	:	o_val <= 16'b0110110001101010;
                14'ha4b 	:	o_val <= 16'b0110110001110001;
                14'ha4c 	:	o_val <= 16'b0110110001110111;
                14'ha4d 	:	o_val <= 16'b0110110001111110;
                14'ha4e 	:	o_val <= 16'b0110110010000101;
                14'ha4f 	:	o_val <= 16'b0110110010001011;
                14'ha50 	:	o_val <= 16'b0110110010010010;
                14'ha51 	:	o_val <= 16'b0110110010011001;
                14'ha52 	:	o_val <= 16'b0110110010011111;
                14'ha53 	:	o_val <= 16'b0110110010100110;
                14'ha54 	:	o_val <= 16'b0110110010101101;
                14'ha55 	:	o_val <= 16'b0110110010110011;
                14'ha56 	:	o_val <= 16'b0110110010111010;
                14'ha57 	:	o_val <= 16'b0110110011000001;
                14'ha58 	:	o_val <= 16'b0110110011000111;
                14'ha59 	:	o_val <= 16'b0110110011001110;
                14'ha5a 	:	o_val <= 16'b0110110011010100;
                14'ha5b 	:	o_val <= 16'b0110110011011011;
                14'ha5c 	:	o_val <= 16'b0110110011100010;
                14'ha5d 	:	o_val <= 16'b0110110011101000;
                14'ha5e 	:	o_val <= 16'b0110110011101111;
                14'ha5f 	:	o_val <= 16'b0110110011110101;
                14'ha60 	:	o_val <= 16'b0110110011111100;
                14'ha61 	:	o_val <= 16'b0110110100000011;
                14'ha62 	:	o_val <= 16'b0110110100001001;
                14'ha63 	:	o_val <= 16'b0110110100010000;
                14'ha64 	:	o_val <= 16'b0110110100010110;
                14'ha65 	:	o_val <= 16'b0110110100011101;
                14'ha66 	:	o_val <= 16'b0110110100100011;
                14'ha67 	:	o_val <= 16'b0110110100101010;
                14'ha68 	:	o_val <= 16'b0110110100110001;
                14'ha69 	:	o_val <= 16'b0110110100110111;
                14'ha6a 	:	o_val <= 16'b0110110100111110;
                14'ha6b 	:	o_val <= 16'b0110110101000100;
                14'ha6c 	:	o_val <= 16'b0110110101001011;
                14'ha6d 	:	o_val <= 16'b0110110101010001;
                14'ha6e 	:	o_val <= 16'b0110110101011000;
                14'ha6f 	:	o_val <= 16'b0110110101011110;
                14'ha70 	:	o_val <= 16'b0110110101100101;
                14'ha71 	:	o_val <= 16'b0110110101101011;
                14'ha72 	:	o_val <= 16'b0110110101110010;
                14'ha73 	:	o_val <= 16'b0110110101111000;
                14'ha74 	:	o_val <= 16'b0110110101111111;
                14'ha75 	:	o_val <= 16'b0110110110000101;
                14'ha76 	:	o_val <= 16'b0110110110001100;
                14'ha77 	:	o_val <= 16'b0110110110010010;
                14'ha78 	:	o_val <= 16'b0110110110011001;
                14'ha79 	:	o_val <= 16'b0110110110011111;
                14'ha7a 	:	o_val <= 16'b0110110110100110;
                14'ha7b 	:	o_val <= 16'b0110110110101100;
                14'ha7c 	:	o_val <= 16'b0110110110110011;
                14'ha7d 	:	o_val <= 16'b0110110110111001;
                14'ha7e 	:	o_val <= 16'b0110110111000000;
                14'ha7f 	:	o_val <= 16'b0110110111000110;
                14'ha80 	:	o_val <= 16'b0110110111001101;
                14'ha81 	:	o_val <= 16'b0110110111010011;
                14'ha82 	:	o_val <= 16'b0110110111011010;
                14'ha83 	:	o_val <= 16'b0110110111100000;
                14'ha84 	:	o_val <= 16'b0110110111100111;
                14'ha85 	:	o_val <= 16'b0110110111101101;
                14'ha86 	:	o_val <= 16'b0110110111110011;
                14'ha87 	:	o_val <= 16'b0110110111111010;
                14'ha88 	:	o_val <= 16'b0110111000000000;
                14'ha89 	:	o_val <= 16'b0110111000000111;
                14'ha8a 	:	o_val <= 16'b0110111000001101;
                14'ha8b 	:	o_val <= 16'b0110111000010100;
                14'ha8c 	:	o_val <= 16'b0110111000011010;
                14'ha8d 	:	o_val <= 16'b0110111000100000;
                14'ha8e 	:	o_val <= 16'b0110111000100111;
                14'ha8f 	:	o_val <= 16'b0110111000101101;
                14'ha90 	:	o_val <= 16'b0110111000110100;
                14'ha91 	:	o_val <= 16'b0110111000111010;
                14'ha92 	:	o_val <= 16'b0110111001000000;
                14'ha93 	:	o_val <= 16'b0110111001000111;
                14'ha94 	:	o_val <= 16'b0110111001001101;
                14'ha95 	:	o_val <= 16'b0110111001010011;
                14'ha96 	:	o_val <= 16'b0110111001011010;
                14'ha97 	:	o_val <= 16'b0110111001100000;
                14'ha98 	:	o_val <= 16'b0110111001100111;
                14'ha99 	:	o_val <= 16'b0110111001101101;
                14'ha9a 	:	o_val <= 16'b0110111001110011;
                14'ha9b 	:	o_val <= 16'b0110111001111010;
                14'ha9c 	:	o_val <= 16'b0110111010000000;
                14'ha9d 	:	o_val <= 16'b0110111010000110;
                14'ha9e 	:	o_val <= 16'b0110111010001101;
                14'ha9f 	:	o_val <= 16'b0110111010010011;
                14'haa0 	:	o_val <= 16'b0110111010011001;
                14'haa1 	:	o_val <= 16'b0110111010100000;
                14'haa2 	:	o_val <= 16'b0110111010100110;
                14'haa3 	:	o_val <= 16'b0110111010101100;
                14'haa4 	:	o_val <= 16'b0110111010110011;
                14'haa5 	:	o_val <= 16'b0110111010111001;
                14'haa6 	:	o_val <= 16'b0110111010111111;
                14'haa7 	:	o_val <= 16'b0110111011000110;
                14'haa8 	:	o_val <= 16'b0110111011001100;
                14'haa9 	:	o_val <= 16'b0110111011010010;
                14'haaa 	:	o_val <= 16'b0110111011011000;
                14'haab 	:	o_val <= 16'b0110111011011111;
                14'haac 	:	o_val <= 16'b0110111011100101;
                14'haad 	:	o_val <= 16'b0110111011101011;
                14'haae 	:	o_val <= 16'b0110111011110001;
                14'haaf 	:	o_val <= 16'b0110111011111000;
                14'hab0 	:	o_val <= 16'b0110111011111110;
                14'hab1 	:	o_val <= 16'b0110111100000100;
                14'hab2 	:	o_val <= 16'b0110111100001011;
                14'hab3 	:	o_val <= 16'b0110111100010001;
                14'hab4 	:	o_val <= 16'b0110111100010111;
                14'hab5 	:	o_val <= 16'b0110111100011101;
                14'hab6 	:	o_val <= 16'b0110111100100011;
                14'hab7 	:	o_val <= 16'b0110111100101010;
                14'hab8 	:	o_val <= 16'b0110111100110000;
                14'hab9 	:	o_val <= 16'b0110111100110110;
                14'haba 	:	o_val <= 16'b0110111100111100;
                14'habb 	:	o_val <= 16'b0110111101000011;
                14'habc 	:	o_val <= 16'b0110111101001001;
                14'habd 	:	o_val <= 16'b0110111101001111;
                14'habe 	:	o_val <= 16'b0110111101010101;
                14'habf 	:	o_val <= 16'b0110111101011011;
                14'hac0 	:	o_val <= 16'b0110111101100010;
                14'hac1 	:	o_val <= 16'b0110111101101000;
                14'hac2 	:	o_val <= 16'b0110111101101110;
                14'hac3 	:	o_val <= 16'b0110111101110100;
                14'hac4 	:	o_val <= 16'b0110111101111010;
                14'hac5 	:	o_val <= 16'b0110111110000001;
                14'hac6 	:	o_val <= 16'b0110111110000111;
                14'hac7 	:	o_val <= 16'b0110111110001101;
                14'hac8 	:	o_val <= 16'b0110111110010011;
                14'hac9 	:	o_val <= 16'b0110111110011001;
                14'haca 	:	o_val <= 16'b0110111110011111;
                14'hacb 	:	o_val <= 16'b0110111110100101;
                14'hacc 	:	o_val <= 16'b0110111110101100;
                14'hacd 	:	o_val <= 16'b0110111110110010;
                14'hace 	:	o_val <= 16'b0110111110111000;
                14'hacf 	:	o_val <= 16'b0110111110111110;
                14'had0 	:	o_val <= 16'b0110111111000100;
                14'had1 	:	o_val <= 16'b0110111111001010;
                14'had2 	:	o_val <= 16'b0110111111010000;
                14'had3 	:	o_val <= 16'b0110111111010110;
                14'had4 	:	o_val <= 16'b0110111111011101;
                14'had5 	:	o_val <= 16'b0110111111100011;
                14'had6 	:	o_val <= 16'b0110111111101001;
                14'had7 	:	o_val <= 16'b0110111111101111;
                14'had8 	:	o_val <= 16'b0110111111110101;
                14'had9 	:	o_val <= 16'b0110111111111011;
                14'hada 	:	o_val <= 16'b0111000000000001;
                14'hadb 	:	o_val <= 16'b0111000000000111;
                14'hadc 	:	o_val <= 16'b0111000000001101;
                14'hadd 	:	o_val <= 16'b0111000000010011;
                14'hade 	:	o_val <= 16'b0111000000011001;
                14'hadf 	:	o_val <= 16'b0111000000100000;
                14'hae0 	:	o_val <= 16'b0111000000100110;
                14'hae1 	:	o_val <= 16'b0111000000101100;
                14'hae2 	:	o_val <= 16'b0111000000110010;
                14'hae3 	:	o_val <= 16'b0111000000111000;
                14'hae4 	:	o_val <= 16'b0111000000111110;
                14'hae5 	:	o_val <= 16'b0111000001000100;
                14'hae6 	:	o_val <= 16'b0111000001001010;
                14'hae7 	:	o_val <= 16'b0111000001010000;
                14'hae8 	:	o_val <= 16'b0111000001010110;
                14'hae9 	:	o_val <= 16'b0111000001011100;
                14'haea 	:	o_val <= 16'b0111000001100010;
                14'haeb 	:	o_val <= 16'b0111000001101000;
                14'haec 	:	o_val <= 16'b0111000001101110;
                14'haed 	:	o_val <= 16'b0111000001110100;
                14'haee 	:	o_val <= 16'b0111000001111010;
                14'haef 	:	o_val <= 16'b0111000010000000;
                14'haf0 	:	o_val <= 16'b0111000010000110;
                14'haf1 	:	o_val <= 16'b0111000010001100;
                14'haf2 	:	o_val <= 16'b0111000010010010;
                14'haf3 	:	o_val <= 16'b0111000010011000;
                14'haf4 	:	o_val <= 16'b0111000010011110;
                14'haf5 	:	o_val <= 16'b0111000010100100;
                14'haf6 	:	o_val <= 16'b0111000010101010;
                14'haf7 	:	o_val <= 16'b0111000010110000;
                14'haf8 	:	o_val <= 16'b0111000010110110;
                14'haf9 	:	o_val <= 16'b0111000010111100;
                14'hafa 	:	o_val <= 16'b0111000011000010;
                14'hafb 	:	o_val <= 16'b0111000011001000;
                14'hafc 	:	o_val <= 16'b0111000011001110;
                14'hafd 	:	o_val <= 16'b0111000011010011;
                14'hafe 	:	o_val <= 16'b0111000011011001;
                14'haff 	:	o_val <= 16'b0111000011011111;
                14'hb00 	:	o_val <= 16'b0111000011100101;
                14'hb01 	:	o_val <= 16'b0111000011101011;
                14'hb02 	:	o_val <= 16'b0111000011110001;
                14'hb03 	:	o_val <= 16'b0111000011110111;
                14'hb04 	:	o_val <= 16'b0111000011111101;
                14'hb05 	:	o_val <= 16'b0111000100000011;
                14'hb06 	:	o_val <= 16'b0111000100001001;
                14'hb07 	:	o_val <= 16'b0111000100001111;
                14'hb08 	:	o_val <= 16'b0111000100010100;
                14'hb09 	:	o_val <= 16'b0111000100011010;
                14'hb0a 	:	o_val <= 16'b0111000100100000;
                14'hb0b 	:	o_val <= 16'b0111000100100110;
                14'hb0c 	:	o_val <= 16'b0111000100101100;
                14'hb0d 	:	o_val <= 16'b0111000100110010;
                14'hb0e 	:	o_val <= 16'b0111000100111000;
                14'hb0f 	:	o_val <= 16'b0111000100111110;
                14'hb10 	:	o_val <= 16'b0111000101000011;
                14'hb11 	:	o_val <= 16'b0111000101001001;
                14'hb12 	:	o_val <= 16'b0111000101001111;
                14'hb13 	:	o_val <= 16'b0111000101010101;
                14'hb14 	:	o_val <= 16'b0111000101011011;
                14'hb15 	:	o_val <= 16'b0111000101100001;
                14'hb16 	:	o_val <= 16'b0111000101100111;
                14'hb17 	:	o_val <= 16'b0111000101101100;
                14'hb18 	:	o_val <= 16'b0111000101110010;
                14'hb19 	:	o_val <= 16'b0111000101111000;
                14'hb1a 	:	o_val <= 16'b0111000101111110;
                14'hb1b 	:	o_val <= 16'b0111000110000100;
                14'hb1c 	:	o_val <= 16'b0111000110001001;
                14'hb1d 	:	o_val <= 16'b0111000110001111;
                14'hb1e 	:	o_val <= 16'b0111000110010101;
                14'hb1f 	:	o_val <= 16'b0111000110011011;
                14'hb20 	:	o_val <= 16'b0111000110100001;
                14'hb21 	:	o_val <= 16'b0111000110100110;
                14'hb22 	:	o_val <= 16'b0111000110101100;
                14'hb23 	:	o_val <= 16'b0111000110110010;
                14'hb24 	:	o_val <= 16'b0111000110111000;
                14'hb25 	:	o_val <= 16'b0111000110111101;
                14'hb26 	:	o_val <= 16'b0111000111000011;
                14'hb27 	:	o_val <= 16'b0111000111001001;
                14'hb28 	:	o_val <= 16'b0111000111001111;
                14'hb29 	:	o_val <= 16'b0111000111010100;
                14'hb2a 	:	o_val <= 16'b0111000111011010;
                14'hb2b 	:	o_val <= 16'b0111000111100000;
                14'hb2c 	:	o_val <= 16'b0111000111100110;
                14'hb2d 	:	o_val <= 16'b0111000111101011;
                14'hb2e 	:	o_val <= 16'b0111000111110001;
                14'hb2f 	:	o_val <= 16'b0111000111110111;
                14'hb30 	:	o_val <= 16'b0111000111111101;
                14'hb31 	:	o_val <= 16'b0111001000000010;
                14'hb32 	:	o_val <= 16'b0111001000001000;
                14'hb33 	:	o_val <= 16'b0111001000001110;
                14'hb34 	:	o_val <= 16'b0111001000010011;
                14'hb35 	:	o_val <= 16'b0111001000011001;
                14'hb36 	:	o_val <= 16'b0111001000011111;
                14'hb37 	:	o_val <= 16'b0111001000100100;
                14'hb38 	:	o_val <= 16'b0111001000101010;
                14'hb39 	:	o_val <= 16'b0111001000110000;
                14'hb3a 	:	o_val <= 16'b0111001000110110;
                14'hb3b 	:	o_val <= 16'b0111001000111011;
                14'hb3c 	:	o_val <= 16'b0111001001000001;
                14'hb3d 	:	o_val <= 16'b0111001001000111;
                14'hb3e 	:	o_val <= 16'b0111001001001100;
                14'hb3f 	:	o_val <= 16'b0111001001010010;
                14'hb40 	:	o_val <= 16'b0111001001010111;
                14'hb41 	:	o_val <= 16'b0111001001011101;
                14'hb42 	:	o_val <= 16'b0111001001100011;
                14'hb43 	:	o_val <= 16'b0111001001101000;
                14'hb44 	:	o_val <= 16'b0111001001101110;
                14'hb45 	:	o_val <= 16'b0111001001110100;
                14'hb46 	:	o_val <= 16'b0111001001111001;
                14'hb47 	:	o_val <= 16'b0111001001111111;
                14'hb48 	:	o_val <= 16'b0111001010000101;
                14'hb49 	:	o_val <= 16'b0111001010001010;
                14'hb4a 	:	o_val <= 16'b0111001010010000;
                14'hb4b 	:	o_val <= 16'b0111001010010101;
                14'hb4c 	:	o_val <= 16'b0111001010011011;
                14'hb4d 	:	o_val <= 16'b0111001010100001;
                14'hb4e 	:	o_val <= 16'b0111001010100110;
                14'hb4f 	:	o_val <= 16'b0111001010101100;
                14'hb50 	:	o_val <= 16'b0111001010110001;
                14'hb51 	:	o_val <= 16'b0111001010110111;
                14'hb52 	:	o_val <= 16'b0111001010111100;
                14'hb53 	:	o_val <= 16'b0111001011000010;
                14'hb54 	:	o_val <= 16'b0111001011001000;
                14'hb55 	:	o_val <= 16'b0111001011001101;
                14'hb56 	:	o_val <= 16'b0111001011010011;
                14'hb57 	:	o_val <= 16'b0111001011011000;
                14'hb58 	:	o_val <= 16'b0111001011011110;
                14'hb59 	:	o_val <= 16'b0111001011100011;
                14'hb5a 	:	o_val <= 16'b0111001011101001;
                14'hb5b 	:	o_val <= 16'b0111001011101110;
                14'hb5c 	:	o_val <= 16'b0111001011110100;
                14'hb5d 	:	o_val <= 16'b0111001011111001;
                14'hb5e 	:	o_val <= 16'b0111001011111111;
                14'hb5f 	:	o_val <= 16'b0111001100000101;
                14'hb60 	:	o_val <= 16'b0111001100001010;
                14'hb61 	:	o_val <= 16'b0111001100010000;
                14'hb62 	:	o_val <= 16'b0111001100010101;
                14'hb63 	:	o_val <= 16'b0111001100011011;
                14'hb64 	:	o_val <= 16'b0111001100100000;
                14'hb65 	:	o_val <= 16'b0111001100100110;
                14'hb66 	:	o_val <= 16'b0111001100101011;
                14'hb67 	:	o_val <= 16'b0111001100110000;
                14'hb68 	:	o_val <= 16'b0111001100110110;
                14'hb69 	:	o_val <= 16'b0111001100111011;
                14'hb6a 	:	o_val <= 16'b0111001101000001;
                14'hb6b 	:	o_val <= 16'b0111001101000110;
                14'hb6c 	:	o_val <= 16'b0111001101001100;
                14'hb6d 	:	o_val <= 16'b0111001101010001;
                14'hb6e 	:	o_val <= 16'b0111001101010111;
                14'hb6f 	:	o_val <= 16'b0111001101011100;
                14'hb70 	:	o_val <= 16'b0111001101100010;
                14'hb71 	:	o_val <= 16'b0111001101100111;
                14'hb72 	:	o_val <= 16'b0111001101101100;
                14'hb73 	:	o_val <= 16'b0111001101110010;
                14'hb74 	:	o_val <= 16'b0111001101110111;
                14'hb75 	:	o_val <= 16'b0111001101111101;
                14'hb76 	:	o_val <= 16'b0111001110000010;
                14'hb77 	:	o_val <= 16'b0111001110001000;
                14'hb78 	:	o_val <= 16'b0111001110001101;
                14'hb79 	:	o_val <= 16'b0111001110010010;
                14'hb7a 	:	o_val <= 16'b0111001110011000;
                14'hb7b 	:	o_val <= 16'b0111001110011101;
                14'hb7c 	:	o_val <= 16'b0111001110100011;
                14'hb7d 	:	o_val <= 16'b0111001110101000;
                14'hb7e 	:	o_val <= 16'b0111001110101101;
                14'hb7f 	:	o_val <= 16'b0111001110110011;
                14'hb80 	:	o_val <= 16'b0111001110111000;
                14'hb81 	:	o_val <= 16'b0111001110111101;
                14'hb82 	:	o_val <= 16'b0111001111000011;
                14'hb83 	:	o_val <= 16'b0111001111001000;
                14'hb84 	:	o_val <= 16'b0111001111001110;
                14'hb85 	:	o_val <= 16'b0111001111010011;
                14'hb86 	:	o_val <= 16'b0111001111011000;
                14'hb87 	:	o_val <= 16'b0111001111011110;
                14'hb88 	:	o_val <= 16'b0111001111100011;
                14'hb89 	:	o_val <= 16'b0111001111101000;
                14'hb8a 	:	o_val <= 16'b0111001111101110;
                14'hb8b 	:	o_val <= 16'b0111001111110011;
                14'hb8c 	:	o_val <= 16'b0111001111111000;
                14'hb8d 	:	o_val <= 16'b0111001111111110;
                14'hb8e 	:	o_val <= 16'b0111010000000011;
                14'hb8f 	:	o_val <= 16'b0111010000001000;
                14'hb90 	:	o_val <= 16'b0111010000001101;
                14'hb91 	:	o_val <= 16'b0111010000010011;
                14'hb92 	:	o_val <= 16'b0111010000011000;
                14'hb93 	:	o_val <= 16'b0111010000011101;
                14'hb94 	:	o_val <= 16'b0111010000100011;
                14'hb95 	:	o_val <= 16'b0111010000101000;
                14'hb96 	:	o_val <= 16'b0111010000101101;
                14'hb97 	:	o_val <= 16'b0111010000110010;
                14'hb98 	:	o_val <= 16'b0111010000111000;
                14'hb99 	:	o_val <= 16'b0111010000111101;
                14'hb9a 	:	o_val <= 16'b0111010001000010;
                14'hb9b 	:	o_val <= 16'b0111010001001000;
                14'hb9c 	:	o_val <= 16'b0111010001001101;
                14'hb9d 	:	o_val <= 16'b0111010001010010;
                14'hb9e 	:	o_val <= 16'b0111010001010111;
                14'hb9f 	:	o_val <= 16'b0111010001011100;
                14'hba0 	:	o_val <= 16'b0111010001100010;
                14'hba1 	:	o_val <= 16'b0111010001100111;
                14'hba2 	:	o_val <= 16'b0111010001101100;
                14'hba3 	:	o_val <= 16'b0111010001110001;
                14'hba4 	:	o_val <= 16'b0111010001110111;
                14'hba5 	:	o_val <= 16'b0111010001111100;
                14'hba6 	:	o_val <= 16'b0111010010000001;
                14'hba7 	:	o_val <= 16'b0111010010000110;
                14'hba8 	:	o_val <= 16'b0111010010001011;
                14'hba9 	:	o_val <= 16'b0111010010010001;
                14'hbaa 	:	o_val <= 16'b0111010010010110;
                14'hbab 	:	o_val <= 16'b0111010010011011;
                14'hbac 	:	o_val <= 16'b0111010010100000;
                14'hbad 	:	o_val <= 16'b0111010010100101;
                14'hbae 	:	o_val <= 16'b0111010010101011;
                14'hbaf 	:	o_val <= 16'b0111010010110000;
                14'hbb0 	:	o_val <= 16'b0111010010110101;
                14'hbb1 	:	o_val <= 16'b0111010010111010;
                14'hbb2 	:	o_val <= 16'b0111010010111111;
                14'hbb3 	:	o_val <= 16'b0111010011000100;
                14'hbb4 	:	o_val <= 16'b0111010011001001;
                14'hbb5 	:	o_val <= 16'b0111010011001111;
                14'hbb6 	:	o_val <= 16'b0111010011010100;
                14'hbb7 	:	o_val <= 16'b0111010011011001;
                14'hbb8 	:	o_val <= 16'b0111010011011110;
                14'hbb9 	:	o_val <= 16'b0111010011100011;
                14'hbba 	:	o_val <= 16'b0111010011101000;
                14'hbbb 	:	o_val <= 16'b0111010011101101;
                14'hbbc 	:	o_val <= 16'b0111010011110010;
                14'hbbd 	:	o_val <= 16'b0111010011111000;
                14'hbbe 	:	o_val <= 16'b0111010011111101;
                14'hbbf 	:	o_val <= 16'b0111010100000010;
                14'hbc0 	:	o_val <= 16'b0111010100000111;
                14'hbc1 	:	o_val <= 16'b0111010100001100;
                14'hbc2 	:	o_val <= 16'b0111010100010001;
                14'hbc3 	:	o_val <= 16'b0111010100010110;
                14'hbc4 	:	o_val <= 16'b0111010100011011;
                14'hbc5 	:	o_val <= 16'b0111010100100000;
                14'hbc6 	:	o_val <= 16'b0111010100100101;
                14'hbc7 	:	o_val <= 16'b0111010100101010;
                14'hbc8 	:	o_val <= 16'b0111010100101111;
                14'hbc9 	:	o_val <= 16'b0111010100110101;
                14'hbca 	:	o_val <= 16'b0111010100111010;
                14'hbcb 	:	o_val <= 16'b0111010100111111;
                14'hbcc 	:	o_val <= 16'b0111010101000100;
                14'hbcd 	:	o_val <= 16'b0111010101001001;
                14'hbce 	:	o_val <= 16'b0111010101001110;
                14'hbcf 	:	o_val <= 16'b0111010101010011;
                14'hbd0 	:	o_val <= 16'b0111010101011000;
                14'hbd1 	:	o_val <= 16'b0111010101011101;
                14'hbd2 	:	o_val <= 16'b0111010101100010;
                14'hbd3 	:	o_val <= 16'b0111010101100111;
                14'hbd4 	:	o_val <= 16'b0111010101101100;
                14'hbd5 	:	o_val <= 16'b0111010101110001;
                14'hbd6 	:	o_val <= 16'b0111010101110110;
                14'hbd7 	:	o_val <= 16'b0111010101111011;
                14'hbd8 	:	o_val <= 16'b0111010110000000;
                14'hbd9 	:	o_val <= 16'b0111010110000101;
                14'hbda 	:	o_val <= 16'b0111010110001010;
                14'hbdb 	:	o_val <= 16'b0111010110001111;
                14'hbdc 	:	o_val <= 16'b0111010110010100;
                14'hbdd 	:	o_val <= 16'b0111010110011001;
                14'hbde 	:	o_val <= 16'b0111010110011110;
                14'hbdf 	:	o_val <= 16'b0111010110100011;
                14'hbe0 	:	o_val <= 16'b0111010110100111;
                14'hbe1 	:	o_val <= 16'b0111010110101100;
                14'hbe2 	:	o_val <= 16'b0111010110110001;
                14'hbe3 	:	o_val <= 16'b0111010110110110;
                14'hbe4 	:	o_val <= 16'b0111010110111011;
                14'hbe5 	:	o_val <= 16'b0111010111000000;
                14'hbe6 	:	o_val <= 16'b0111010111000101;
                14'hbe7 	:	o_val <= 16'b0111010111001010;
                14'hbe8 	:	o_val <= 16'b0111010111001111;
                14'hbe9 	:	o_val <= 16'b0111010111010100;
                14'hbea 	:	o_val <= 16'b0111010111011001;
                14'hbeb 	:	o_val <= 16'b0111010111011110;
                14'hbec 	:	o_val <= 16'b0111010111100011;
                14'hbed 	:	o_val <= 16'b0111010111100111;
                14'hbee 	:	o_val <= 16'b0111010111101100;
                14'hbef 	:	o_val <= 16'b0111010111110001;
                14'hbf0 	:	o_val <= 16'b0111010111110110;
                14'hbf1 	:	o_val <= 16'b0111010111111011;
                14'hbf2 	:	o_val <= 16'b0111011000000000;
                14'hbf3 	:	o_val <= 16'b0111011000000101;
                14'hbf4 	:	o_val <= 16'b0111011000001010;
                14'hbf5 	:	o_val <= 16'b0111011000001110;
                14'hbf6 	:	o_val <= 16'b0111011000010011;
                14'hbf7 	:	o_val <= 16'b0111011000011000;
                14'hbf8 	:	o_val <= 16'b0111011000011101;
                14'hbf9 	:	o_val <= 16'b0111011000100010;
                14'hbfa 	:	o_val <= 16'b0111011000100111;
                14'hbfb 	:	o_val <= 16'b0111011000101011;
                14'hbfc 	:	o_val <= 16'b0111011000110000;
                14'hbfd 	:	o_val <= 16'b0111011000110101;
                14'hbfe 	:	o_val <= 16'b0111011000111010;
                14'hbff 	:	o_val <= 16'b0111011000111111;
                14'hc00 	:	o_val <= 16'b0111011001000100;
                14'hc01 	:	o_val <= 16'b0111011001001000;
                14'hc02 	:	o_val <= 16'b0111011001001101;
                14'hc03 	:	o_val <= 16'b0111011001010010;
                14'hc04 	:	o_val <= 16'b0111011001010111;
                14'hc05 	:	o_val <= 16'b0111011001011100;
                14'hc06 	:	o_val <= 16'b0111011001100000;
                14'hc07 	:	o_val <= 16'b0111011001100101;
                14'hc08 	:	o_val <= 16'b0111011001101010;
                14'hc09 	:	o_val <= 16'b0111011001101111;
                14'hc0a 	:	o_val <= 16'b0111011001110011;
                14'hc0b 	:	o_val <= 16'b0111011001111000;
                14'hc0c 	:	o_val <= 16'b0111011001111101;
                14'hc0d 	:	o_val <= 16'b0111011010000010;
                14'hc0e 	:	o_val <= 16'b0111011010000110;
                14'hc0f 	:	o_val <= 16'b0111011010001011;
                14'hc10 	:	o_val <= 16'b0111011010010000;
                14'hc11 	:	o_val <= 16'b0111011010010101;
                14'hc12 	:	o_val <= 16'b0111011010011001;
                14'hc13 	:	o_val <= 16'b0111011010011110;
                14'hc14 	:	o_val <= 16'b0111011010100011;
                14'hc15 	:	o_val <= 16'b0111011010101000;
                14'hc16 	:	o_val <= 16'b0111011010101100;
                14'hc17 	:	o_val <= 16'b0111011010110001;
                14'hc18 	:	o_val <= 16'b0111011010110110;
                14'hc19 	:	o_val <= 16'b0111011010111010;
                14'hc1a 	:	o_val <= 16'b0111011010111111;
                14'hc1b 	:	o_val <= 16'b0111011011000100;
                14'hc1c 	:	o_val <= 16'b0111011011001000;
                14'hc1d 	:	o_val <= 16'b0111011011001101;
                14'hc1e 	:	o_val <= 16'b0111011011010010;
                14'hc1f 	:	o_val <= 16'b0111011011010110;
                14'hc20 	:	o_val <= 16'b0111011011011011;
                14'hc21 	:	o_val <= 16'b0111011011100000;
                14'hc22 	:	o_val <= 16'b0111011011100100;
                14'hc23 	:	o_val <= 16'b0111011011101001;
                14'hc24 	:	o_val <= 16'b0111011011101110;
                14'hc25 	:	o_val <= 16'b0111011011110010;
                14'hc26 	:	o_val <= 16'b0111011011110111;
                14'hc27 	:	o_val <= 16'b0111011011111100;
                14'hc28 	:	o_val <= 16'b0111011100000000;
                14'hc29 	:	o_val <= 16'b0111011100000101;
                14'hc2a 	:	o_val <= 16'b0111011100001010;
                14'hc2b 	:	o_val <= 16'b0111011100001110;
                14'hc2c 	:	o_val <= 16'b0111011100010011;
                14'hc2d 	:	o_val <= 16'b0111011100010111;
                14'hc2e 	:	o_val <= 16'b0111011100011100;
                14'hc2f 	:	o_val <= 16'b0111011100100001;
                14'hc30 	:	o_val <= 16'b0111011100100101;
                14'hc31 	:	o_val <= 16'b0111011100101010;
                14'hc32 	:	o_val <= 16'b0111011100101110;
                14'hc33 	:	o_val <= 16'b0111011100110011;
                14'hc34 	:	o_val <= 16'b0111011100111000;
                14'hc35 	:	o_val <= 16'b0111011100111100;
                14'hc36 	:	o_val <= 16'b0111011101000001;
                14'hc37 	:	o_val <= 16'b0111011101000101;
                14'hc38 	:	o_val <= 16'b0111011101001010;
                14'hc39 	:	o_val <= 16'b0111011101001110;
                14'hc3a 	:	o_val <= 16'b0111011101010011;
                14'hc3b 	:	o_val <= 16'b0111011101010111;
                14'hc3c 	:	o_val <= 16'b0111011101011100;
                14'hc3d 	:	o_val <= 16'b0111011101100000;
                14'hc3e 	:	o_val <= 16'b0111011101100101;
                14'hc3f 	:	o_val <= 16'b0111011101101010;
                14'hc40 	:	o_val <= 16'b0111011101101110;
                14'hc41 	:	o_val <= 16'b0111011101110011;
                14'hc42 	:	o_val <= 16'b0111011101110111;
                14'hc43 	:	o_val <= 16'b0111011101111100;
                14'hc44 	:	o_val <= 16'b0111011110000000;
                14'hc45 	:	o_val <= 16'b0111011110000101;
                14'hc46 	:	o_val <= 16'b0111011110001001;
                14'hc47 	:	o_val <= 16'b0111011110001110;
                14'hc48 	:	o_val <= 16'b0111011110010010;
                14'hc49 	:	o_val <= 16'b0111011110010111;
                14'hc4a 	:	o_val <= 16'b0111011110011011;
                14'hc4b 	:	o_val <= 16'b0111011110100000;
                14'hc4c 	:	o_val <= 16'b0111011110100100;
                14'hc4d 	:	o_val <= 16'b0111011110101000;
                14'hc4e 	:	o_val <= 16'b0111011110101101;
                14'hc4f 	:	o_val <= 16'b0111011110110001;
                14'hc50 	:	o_val <= 16'b0111011110110110;
                14'hc51 	:	o_val <= 16'b0111011110111010;
                14'hc52 	:	o_val <= 16'b0111011110111111;
                14'hc53 	:	o_val <= 16'b0111011111000011;
                14'hc54 	:	o_val <= 16'b0111011111001000;
                14'hc55 	:	o_val <= 16'b0111011111001100;
                14'hc56 	:	o_val <= 16'b0111011111010000;
                14'hc57 	:	o_val <= 16'b0111011111010101;
                14'hc58 	:	o_val <= 16'b0111011111011001;
                14'hc59 	:	o_val <= 16'b0111011111011110;
                14'hc5a 	:	o_val <= 16'b0111011111100010;
                14'hc5b 	:	o_val <= 16'b0111011111100110;
                14'hc5c 	:	o_val <= 16'b0111011111101011;
                14'hc5d 	:	o_val <= 16'b0111011111101111;
                14'hc5e 	:	o_val <= 16'b0111011111110100;
                14'hc5f 	:	o_val <= 16'b0111011111111000;
                14'hc60 	:	o_val <= 16'b0111011111111100;
                14'hc61 	:	o_val <= 16'b0111100000000001;
                14'hc62 	:	o_val <= 16'b0111100000000101;
                14'hc63 	:	o_val <= 16'b0111100000001010;
                14'hc64 	:	o_val <= 16'b0111100000001110;
                14'hc65 	:	o_val <= 16'b0111100000010010;
                14'hc66 	:	o_val <= 16'b0111100000010111;
                14'hc67 	:	o_val <= 16'b0111100000011011;
                14'hc68 	:	o_val <= 16'b0111100000011111;
                14'hc69 	:	o_val <= 16'b0111100000100100;
                14'hc6a 	:	o_val <= 16'b0111100000101000;
                14'hc6b 	:	o_val <= 16'b0111100000101100;
                14'hc6c 	:	o_val <= 16'b0111100000110001;
                14'hc6d 	:	o_val <= 16'b0111100000110101;
                14'hc6e 	:	o_val <= 16'b0111100000111001;
                14'hc6f 	:	o_val <= 16'b0111100000111110;
                14'hc70 	:	o_val <= 16'b0111100001000010;
                14'hc71 	:	o_val <= 16'b0111100001000110;
                14'hc72 	:	o_val <= 16'b0111100001001010;
                14'hc73 	:	o_val <= 16'b0111100001001111;
                14'hc74 	:	o_val <= 16'b0111100001010011;
                14'hc75 	:	o_val <= 16'b0111100001010111;
                14'hc76 	:	o_val <= 16'b0111100001011100;
                14'hc77 	:	o_val <= 16'b0111100001100000;
                14'hc78 	:	o_val <= 16'b0111100001100100;
                14'hc79 	:	o_val <= 16'b0111100001101000;
                14'hc7a 	:	o_val <= 16'b0111100001101101;
                14'hc7b 	:	o_val <= 16'b0111100001110001;
                14'hc7c 	:	o_val <= 16'b0111100001110101;
                14'hc7d 	:	o_val <= 16'b0111100001111001;
                14'hc7e 	:	o_val <= 16'b0111100001111110;
                14'hc7f 	:	o_val <= 16'b0111100010000010;
                14'hc80 	:	o_val <= 16'b0111100010000110;
                14'hc81 	:	o_val <= 16'b0111100010001010;
                14'hc82 	:	o_val <= 16'b0111100010001111;
                14'hc83 	:	o_val <= 16'b0111100010010011;
                14'hc84 	:	o_val <= 16'b0111100010010111;
                14'hc85 	:	o_val <= 16'b0111100010011011;
                14'hc86 	:	o_val <= 16'b0111100010011111;
                14'hc87 	:	o_val <= 16'b0111100010100100;
                14'hc88 	:	o_val <= 16'b0111100010101000;
                14'hc89 	:	o_val <= 16'b0111100010101100;
                14'hc8a 	:	o_val <= 16'b0111100010110000;
                14'hc8b 	:	o_val <= 16'b0111100010110100;
                14'hc8c 	:	o_val <= 16'b0111100010111001;
                14'hc8d 	:	o_val <= 16'b0111100010111101;
                14'hc8e 	:	o_val <= 16'b0111100011000001;
                14'hc8f 	:	o_val <= 16'b0111100011000101;
                14'hc90 	:	o_val <= 16'b0111100011001001;
                14'hc91 	:	o_val <= 16'b0111100011001101;
                14'hc92 	:	o_val <= 16'b0111100011010010;
                14'hc93 	:	o_val <= 16'b0111100011010110;
                14'hc94 	:	o_val <= 16'b0111100011011010;
                14'hc95 	:	o_val <= 16'b0111100011011110;
                14'hc96 	:	o_val <= 16'b0111100011100010;
                14'hc97 	:	o_val <= 16'b0111100011100110;
                14'hc98 	:	o_val <= 16'b0111100011101010;
                14'hc99 	:	o_val <= 16'b0111100011101110;
                14'hc9a 	:	o_val <= 16'b0111100011110011;
                14'hc9b 	:	o_val <= 16'b0111100011110111;
                14'hc9c 	:	o_val <= 16'b0111100011111011;
                14'hc9d 	:	o_val <= 16'b0111100011111111;
                14'hc9e 	:	o_val <= 16'b0111100100000011;
                14'hc9f 	:	o_val <= 16'b0111100100000111;
                14'hca0 	:	o_val <= 16'b0111100100001011;
                14'hca1 	:	o_val <= 16'b0111100100001111;
                14'hca2 	:	o_val <= 16'b0111100100010011;
                14'hca3 	:	o_val <= 16'b0111100100010111;
                14'hca4 	:	o_val <= 16'b0111100100011100;
                14'hca5 	:	o_val <= 16'b0111100100100000;
                14'hca6 	:	o_val <= 16'b0111100100100100;
                14'hca7 	:	o_val <= 16'b0111100100101000;
                14'hca8 	:	o_val <= 16'b0111100100101100;
                14'hca9 	:	o_val <= 16'b0111100100110000;
                14'hcaa 	:	o_val <= 16'b0111100100110100;
                14'hcab 	:	o_val <= 16'b0111100100111000;
                14'hcac 	:	o_val <= 16'b0111100100111100;
                14'hcad 	:	o_val <= 16'b0111100101000000;
                14'hcae 	:	o_val <= 16'b0111100101000100;
                14'hcaf 	:	o_val <= 16'b0111100101001000;
                14'hcb0 	:	o_val <= 16'b0111100101001100;
                14'hcb1 	:	o_val <= 16'b0111100101010000;
                14'hcb2 	:	o_val <= 16'b0111100101010100;
                14'hcb3 	:	o_val <= 16'b0111100101011000;
                14'hcb4 	:	o_val <= 16'b0111100101011100;
                14'hcb5 	:	o_val <= 16'b0111100101100000;
                14'hcb6 	:	o_val <= 16'b0111100101100100;
                14'hcb7 	:	o_val <= 16'b0111100101101000;
                14'hcb8 	:	o_val <= 16'b0111100101101100;
                14'hcb9 	:	o_val <= 16'b0111100101110000;
                14'hcba 	:	o_val <= 16'b0111100101110100;
                14'hcbb 	:	o_val <= 16'b0111100101111000;
                14'hcbc 	:	o_val <= 16'b0111100101111100;
                14'hcbd 	:	o_val <= 16'b0111100110000000;
                14'hcbe 	:	o_val <= 16'b0111100110000100;
                14'hcbf 	:	o_val <= 16'b0111100110001000;
                14'hcc0 	:	o_val <= 16'b0111100110001100;
                14'hcc1 	:	o_val <= 16'b0111100110010000;
                14'hcc2 	:	o_val <= 16'b0111100110010011;
                14'hcc3 	:	o_val <= 16'b0111100110010111;
                14'hcc4 	:	o_val <= 16'b0111100110011011;
                14'hcc5 	:	o_val <= 16'b0111100110011111;
                14'hcc6 	:	o_val <= 16'b0111100110100011;
                14'hcc7 	:	o_val <= 16'b0111100110100111;
                14'hcc8 	:	o_val <= 16'b0111100110101011;
                14'hcc9 	:	o_val <= 16'b0111100110101111;
                14'hcca 	:	o_val <= 16'b0111100110110011;
                14'hccb 	:	o_val <= 16'b0111100110110111;
                14'hccc 	:	o_val <= 16'b0111100110111011;
                14'hccd 	:	o_val <= 16'b0111100110111110;
                14'hcce 	:	o_val <= 16'b0111100111000010;
                14'hccf 	:	o_val <= 16'b0111100111000110;
                14'hcd0 	:	o_val <= 16'b0111100111001010;
                14'hcd1 	:	o_val <= 16'b0111100111001110;
                14'hcd2 	:	o_val <= 16'b0111100111010010;
                14'hcd3 	:	o_val <= 16'b0111100111010110;
                14'hcd4 	:	o_val <= 16'b0111100111011001;
                14'hcd5 	:	o_val <= 16'b0111100111011101;
                14'hcd6 	:	o_val <= 16'b0111100111100001;
                14'hcd7 	:	o_val <= 16'b0111100111100101;
                14'hcd8 	:	o_val <= 16'b0111100111101001;
                14'hcd9 	:	o_val <= 16'b0111100111101101;
                14'hcda 	:	o_val <= 16'b0111100111110000;
                14'hcdb 	:	o_val <= 16'b0111100111110100;
                14'hcdc 	:	o_val <= 16'b0111100111111000;
                14'hcdd 	:	o_val <= 16'b0111100111111100;
                14'hcde 	:	o_val <= 16'b0111101000000000;
                14'hcdf 	:	o_val <= 16'b0111101000000100;
                14'hce0 	:	o_val <= 16'b0111101000000111;
                14'hce1 	:	o_val <= 16'b0111101000001011;
                14'hce2 	:	o_val <= 16'b0111101000001111;
                14'hce3 	:	o_val <= 16'b0111101000010011;
                14'hce4 	:	o_val <= 16'b0111101000010110;
                14'hce5 	:	o_val <= 16'b0111101000011010;
                14'hce6 	:	o_val <= 16'b0111101000011110;
                14'hce7 	:	o_val <= 16'b0111101000100010;
                14'hce8 	:	o_val <= 16'b0111101000100110;
                14'hce9 	:	o_val <= 16'b0111101000101001;
                14'hcea 	:	o_val <= 16'b0111101000101101;
                14'hceb 	:	o_val <= 16'b0111101000110001;
                14'hcec 	:	o_val <= 16'b0111101000110101;
                14'hced 	:	o_val <= 16'b0111101000111000;
                14'hcee 	:	o_val <= 16'b0111101000111100;
                14'hcef 	:	o_val <= 16'b0111101001000000;
                14'hcf0 	:	o_val <= 16'b0111101001000011;
                14'hcf1 	:	o_val <= 16'b0111101001000111;
                14'hcf2 	:	o_val <= 16'b0111101001001011;
                14'hcf3 	:	o_val <= 16'b0111101001001111;
                14'hcf4 	:	o_val <= 16'b0111101001010010;
                14'hcf5 	:	o_val <= 16'b0111101001010110;
                14'hcf6 	:	o_val <= 16'b0111101001011010;
                14'hcf7 	:	o_val <= 16'b0111101001011101;
                14'hcf8 	:	o_val <= 16'b0111101001100001;
                14'hcf9 	:	o_val <= 16'b0111101001100101;
                14'hcfa 	:	o_val <= 16'b0111101001101000;
                14'hcfb 	:	o_val <= 16'b0111101001101100;
                14'hcfc 	:	o_val <= 16'b0111101001110000;
                14'hcfd 	:	o_val <= 16'b0111101001110011;
                14'hcfe 	:	o_val <= 16'b0111101001110111;
                14'hcff 	:	o_val <= 16'b0111101001111011;
                14'hd00 	:	o_val <= 16'b0111101001111110;
                14'hd01 	:	o_val <= 16'b0111101010000010;
                14'hd02 	:	o_val <= 16'b0111101010000110;
                14'hd03 	:	o_val <= 16'b0111101010001001;
                14'hd04 	:	o_val <= 16'b0111101010001101;
                14'hd05 	:	o_val <= 16'b0111101010010001;
                14'hd06 	:	o_val <= 16'b0111101010010100;
                14'hd07 	:	o_val <= 16'b0111101010011000;
                14'hd08 	:	o_val <= 16'b0111101010011011;
                14'hd09 	:	o_val <= 16'b0111101010011111;
                14'hd0a 	:	o_val <= 16'b0111101010100011;
                14'hd0b 	:	o_val <= 16'b0111101010100110;
                14'hd0c 	:	o_val <= 16'b0111101010101010;
                14'hd0d 	:	o_val <= 16'b0111101010101101;
                14'hd0e 	:	o_val <= 16'b0111101010110001;
                14'hd0f 	:	o_val <= 16'b0111101010110101;
                14'hd10 	:	o_val <= 16'b0111101010111000;
                14'hd11 	:	o_val <= 16'b0111101010111100;
                14'hd12 	:	o_val <= 16'b0111101010111111;
                14'hd13 	:	o_val <= 16'b0111101011000011;
                14'hd14 	:	o_val <= 16'b0111101011000110;
                14'hd15 	:	o_val <= 16'b0111101011001010;
                14'hd16 	:	o_val <= 16'b0111101011001101;
                14'hd17 	:	o_val <= 16'b0111101011010001;
                14'hd18 	:	o_val <= 16'b0111101011010101;
                14'hd19 	:	o_val <= 16'b0111101011011000;
                14'hd1a 	:	o_val <= 16'b0111101011011100;
                14'hd1b 	:	o_val <= 16'b0111101011011111;
                14'hd1c 	:	o_val <= 16'b0111101011100011;
                14'hd1d 	:	o_val <= 16'b0111101011100110;
                14'hd1e 	:	o_val <= 16'b0111101011101010;
                14'hd1f 	:	o_val <= 16'b0111101011101101;
                14'hd20 	:	o_val <= 16'b0111101011110001;
                14'hd21 	:	o_val <= 16'b0111101011110100;
                14'hd22 	:	o_val <= 16'b0111101011111000;
                14'hd23 	:	o_val <= 16'b0111101011111011;
                14'hd24 	:	o_val <= 16'b0111101011111111;
                14'hd25 	:	o_val <= 16'b0111101100000010;
                14'hd26 	:	o_val <= 16'b0111101100000110;
                14'hd27 	:	o_val <= 16'b0111101100001001;
                14'hd28 	:	o_val <= 16'b0111101100001100;
                14'hd29 	:	o_val <= 16'b0111101100010000;
                14'hd2a 	:	o_val <= 16'b0111101100010011;
                14'hd2b 	:	o_val <= 16'b0111101100010111;
                14'hd2c 	:	o_val <= 16'b0111101100011010;
                14'hd2d 	:	o_val <= 16'b0111101100011110;
                14'hd2e 	:	o_val <= 16'b0111101100100001;
                14'hd2f 	:	o_val <= 16'b0111101100100101;
                14'hd30 	:	o_val <= 16'b0111101100101000;
                14'hd31 	:	o_val <= 16'b0111101100101011;
                14'hd32 	:	o_val <= 16'b0111101100101111;
                14'hd33 	:	o_val <= 16'b0111101100110010;
                14'hd34 	:	o_val <= 16'b0111101100110110;
                14'hd35 	:	o_val <= 16'b0111101100111001;
                14'hd36 	:	o_val <= 16'b0111101100111100;
                14'hd37 	:	o_val <= 16'b0111101101000000;
                14'hd38 	:	o_val <= 16'b0111101101000011;
                14'hd39 	:	o_val <= 16'b0111101101000111;
                14'hd3a 	:	o_val <= 16'b0111101101001010;
                14'hd3b 	:	o_val <= 16'b0111101101001101;
                14'hd3c 	:	o_val <= 16'b0111101101010001;
                14'hd3d 	:	o_val <= 16'b0111101101010100;
                14'hd3e 	:	o_val <= 16'b0111101101010111;
                14'hd3f 	:	o_val <= 16'b0111101101011011;
                14'hd40 	:	o_val <= 16'b0111101101011110;
                14'hd41 	:	o_val <= 16'b0111101101100010;
                14'hd42 	:	o_val <= 16'b0111101101100101;
                14'hd43 	:	o_val <= 16'b0111101101101000;
                14'hd44 	:	o_val <= 16'b0111101101101100;
                14'hd45 	:	o_val <= 16'b0111101101101111;
                14'hd46 	:	o_val <= 16'b0111101101110010;
                14'hd47 	:	o_val <= 16'b0111101101110110;
                14'hd48 	:	o_val <= 16'b0111101101111001;
                14'hd49 	:	o_val <= 16'b0111101101111100;
                14'hd4a 	:	o_val <= 16'b0111101101111111;
                14'hd4b 	:	o_val <= 16'b0111101110000011;
                14'hd4c 	:	o_val <= 16'b0111101110000110;
                14'hd4d 	:	o_val <= 16'b0111101110001001;
                14'hd4e 	:	o_val <= 16'b0111101110001101;
                14'hd4f 	:	o_val <= 16'b0111101110010000;
                14'hd50 	:	o_val <= 16'b0111101110010011;
                14'hd51 	:	o_val <= 16'b0111101110010110;
                14'hd52 	:	o_val <= 16'b0111101110011010;
                14'hd53 	:	o_val <= 16'b0111101110011101;
                14'hd54 	:	o_val <= 16'b0111101110100000;
                14'hd55 	:	o_val <= 16'b0111101110100011;
                14'hd56 	:	o_val <= 16'b0111101110100111;
                14'hd57 	:	o_val <= 16'b0111101110101010;
                14'hd58 	:	o_val <= 16'b0111101110101101;
                14'hd59 	:	o_val <= 16'b0111101110110000;
                14'hd5a 	:	o_val <= 16'b0111101110110100;
                14'hd5b 	:	o_val <= 16'b0111101110110111;
                14'hd5c 	:	o_val <= 16'b0111101110111010;
                14'hd5d 	:	o_val <= 16'b0111101110111101;
                14'hd5e 	:	o_val <= 16'b0111101111000001;
                14'hd5f 	:	o_val <= 16'b0111101111000100;
                14'hd60 	:	o_val <= 16'b0111101111000111;
                14'hd61 	:	o_val <= 16'b0111101111001010;
                14'hd62 	:	o_val <= 16'b0111101111001101;
                14'hd63 	:	o_val <= 16'b0111101111010001;
                14'hd64 	:	o_val <= 16'b0111101111010100;
                14'hd65 	:	o_val <= 16'b0111101111010111;
                14'hd66 	:	o_val <= 16'b0111101111011010;
                14'hd67 	:	o_val <= 16'b0111101111011101;
                14'hd68 	:	o_val <= 16'b0111101111100000;
                14'hd69 	:	o_val <= 16'b0111101111100100;
                14'hd6a 	:	o_val <= 16'b0111101111100111;
                14'hd6b 	:	o_val <= 16'b0111101111101010;
                14'hd6c 	:	o_val <= 16'b0111101111101101;
                14'hd6d 	:	o_val <= 16'b0111101111110000;
                14'hd6e 	:	o_val <= 16'b0111101111110011;
                14'hd6f 	:	o_val <= 16'b0111101111110110;
                14'hd70 	:	o_val <= 16'b0111101111111010;
                14'hd71 	:	o_val <= 16'b0111101111111101;
                14'hd72 	:	o_val <= 16'b0111110000000000;
                14'hd73 	:	o_val <= 16'b0111110000000011;
                14'hd74 	:	o_val <= 16'b0111110000000110;
                14'hd75 	:	o_val <= 16'b0111110000001001;
                14'hd76 	:	o_val <= 16'b0111110000001100;
                14'hd77 	:	o_val <= 16'b0111110000001111;
                14'hd78 	:	o_val <= 16'b0111110000010010;
                14'hd79 	:	o_val <= 16'b0111110000010110;
                14'hd7a 	:	o_val <= 16'b0111110000011001;
                14'hd7b 	:	o_val <= 16'b0111110000011100;
                14'hd7c 	:	o_val <= 16'b0111110000011111;
                14'hd7d 	:	o_val <= 16'b0111110000100010;
                14'hd7e 	:	o_val <= 16'b0111110000100101;
                14'hd7f 	:	o_val <= 16'b0111110000101000;
                14'hd80 	:	o_val <= 16'b0111110000101011;
                14'hd81 	:	o_val <= 16'b0111110000101110;
                14'hd82 	:	o_val <= 16'b0111110000110001;
                14'hd83 	:	o_val <= 16'b0111110000110100;
                14'hd84 	:	o_val <= 16'b0111110000110111;
                14'hd85 	:	o_val <= 16'b0111110000111010;
                14'hd86 	:	o_val <= 16'b0111110000111101;
                14'hd87 	:	o_val <= 16'b0111110001000000;
                14'hd88 	:	o_val <= 16'b0111110001000011;
                14'hd89 	:	o_val <= 16'b0111110001000110;
                14'hd8a 	:	o_val <= 16'b0111110001001001;
                14'hd8b 	:	o_val <= 16'b0111110001001100;
                14'hd8c 	:	o_val <= 16'b0111110001001111;
                14'hd8d 	:	o_val <= 16'b0111110001010010;
                14'hd8e 	:	o_val <= 16'b0111110001010101;
                14'hd8f 	:	o_val <= 16'b0111110001011000;
                14'hd90 	:	o_val <= 16'b0111110001011011;
                14'hd91 	:	o_val <= 16'b0111110001011110;
                14'hd92 	:	o_val <= 16'b0111110001100001;
                14'hd93 	:	o_val <= 16'b0111110001100100;
                14'hd94 	:	o_val <= 16'b0111110001100111;
                14'hd95 	:	o_val <= 16'b0111110001101010;
                14'hd96 	:	o_val <= 16'b0111110001101101;
                14'hd97 	:	o_val <= 16'b0111110001110000;
                14'hd98 	:	o_val <= 16'b0111110001110011;
                14'hd99 	:	o_val <= 16'b0111110001110110;
                14'hd9a 	:	o_val <= 16'b0111110001111001;
                14'hd9b 	:	o_val <= 16'b0111110001111100;
                14'hd9c 	:	o_val <= 16'b0111110001111111;
                14'hd9d 	:	o_val <= 16'b0111110010000010;
                14'hd9e 	:	o_val <= 16'b0111110010000100;
                14'hd9f 	:	o_val <= 16'b0111110010000111;
                14'hda0 	:	o_val <= 16'b0111110010001010;
                14'hda1 	:	o_val <= 16'b0111110010001101;
                14'hda2 	:	o_val <= 16'b0111110010010000;
                14'hda3 	:	o_val <= 16'b0111110010010011;
                14'hda4 	:	o_val <= 16'b0111110010010110;
                14'hda5 	:	o_val <= 16'b0111110010011001;
                14'hda6 	:	o_val <= 16'b0111110010011100;
                14'hda7 	:	o_val <= 16'b0111110010011110;
                14'hda8 	:	o_val <= 16'b0111110010100001;
                14'hda9 	:	o_val <= 16'b0111110010100100;
                14'hdaa 	:	o_val <= 16'b0111110010100111;
                14'hdab 	:	o_val <= 16'b0111110010101010;
                14'hdac 	:	o_val <= 16'b0111110010101101;
                14'hdad 	:	o_val <= 16'b0111110010110000;
                14'hdae 	:	o_val <= 16'b0111110010110010;
                14'hdaf 	:	o_val <= 16'b0111110010110101;
                14'hdb0 	:	o_val <= 16'b0111110010111000;
                14'hdb1 	:	o_val <= 16'b0111110010111011;
                14'hdb2 	:	o_val <= 16'b0111110010111110;
                14'hdb3 	:	o_val <= 16'b0111110011000001;
                14'hdb4 	:	o_val <= 16'b0111110011000011;
                14'hdb5 	:	o_val <= 16'b0111110011000110;
                14'hdb6 	:	o_val <= 16'b0111110011001001;
                14'hdb7 	:	o_val <= 16'b0111110011001100;
                14'hdb8 	:	o_val <= 16'b0111110011001111;
                14'hdb9 	:	o_val <= 16'b0111110011010001;
                14'hdba 	:	o_val <= 16'b0111110011010100;
                14'hdbb 	:	o_val <= 16'b0111110011010111;
                14'hdbc 	:	o_val <= 16'b0111110011011010;
                14'hdbd 	:	o_val <= 16'b0111110011011100;
                14'hdbe 	:	o_val <= 16'b0111110011011111;
                14'hdbf 	:	o_val <= 16'b0111110011100010;
                14'hdc0 	:	o_val <= 16'b0111110011100101;
                14'hdc1 	:	o_val <= 16'b0111110011100111;
                14'hdc2 	:	o_val <= 16'b0111110011101010;
                14'hdc3 	:	o_val <= 16'b0111110011101101;
                14'hdc4 	:	o_val <= 16'b0111110011110000;
                14'hdc5 	:	o_val <= 16'b0111110011110010;
                14'hdc6 	:	o_val <= 16'b0111110011110101;
                14'hdc7 	:	o_val <= 16'b0111110011111000;
                14'hdc8 	:	o_val <= 16'b0111110011111011;
                14'hdc9 	:	o_val <= 16'b0111110011111101;
                14'hdca 	:	o_val <= 16'b0111110100000000;
                14'hdcb 	:	o_val <= 16'b0111110100000011;
                14'hdcc 	:	o_val <= 16'b0111110100000101;
                14'hdcd 	:	o_val <= 16'b0111110100001000;
                14'hdce 	:	o_val <= 16'b0111110100001011;
                14'hdcf 	:	o_val <= 16'b0111110100001101;
                14'hdd0 	:	o_val <= 16'b0111110100010000;
                14'hdd1 	:	o_val <= 16'b0111110100010011;
                14'hdd2 	:	o_val <= 16'b0111110100010101;
                14'hdd3 	:	o_val <= 16'b0111110100011000;
                14'hdd4 	:	o_val <= 16'b0111110100011011;
                14'hdd5 	:	o_val <= 16'b0111110100011101;
                14'hdd6 	:	o_val <= 16'b0111110100100000;
                14'hdd7 	:	o_val <= 16'b0111110100100011;
                14'hdd8 	:	o_val <= 16'b0111110100100101;
                14'hdd9 	:	o_val <= 16'b0111110100101000;
                14'hdda 	:	o_val <= 16'b0111110100101011;
                14'hddb 	:	o_val <= 16'b0111110100101101;
                14'hddc 	:	o_val <= 16'b0111110100110000;
                14'hddd 	:	o_val <= 16'b0111110100110010;
                14'hdde 	:	o_val <= 16'b0111110100110101;
                14'hddf 	:	o_val <= 16'b0111110100111000;
                14'hde0 	:	o_val <= 16'b0111110100111010;
                14'hde1 	:	o_val <= 16'b0111110100111101;
                14'hde2 	:	o_val <= 16'b0111110100111111;
                14'hde3 	:	o_val <= 16'b0111110101000010;
                14'hde4 	:	o_val <= 16'b0111110101000101;
                14'hde5 	:	o_val <= 16'b0111110101000111;
                14'hde6 	:	o_val <= 16'b0111110101001010;
                14'hde7 	:	o_val <= 16'b0111110101001100;
                14'hde8 	:	o_val <= 16'b0111110101001111;
                14'hde9 	:	o_val <= 16'b0111110101010010;
                14'hdea 	:	o_val <= 16'b0111110101010100;
                14'hdeb 	:	o_val <= 16'b0111110101010111;
                14'hdec 	:	o_val <= 16'b0111110101011001;
                14'hded 	:	o_val <= 16'b0111110101011100;
                14'hdee 	:	o_val <= 16'b0111110101011110;
                14'hdef 	:	o_val <= 16'b0111110101100001;
                14'hdf0 	:	o_val <= 16'b0111110101100011;
                14'hdf1 	:	o_val <= 16'b0111110101100110;
                14'hdf2 	:	o_val <= 16'b0111110101101000;
                14'hdf3 	:	o_val <= 16'b0111110101101011;
                14'hdf4 	:	o_val <= 16'b0111110101101101;
                14'hdf5 	:	o_val <= 16'b0111110101110000;
                14'hdf6 	:	o_val <= 16'b0111110101110010;
                14'hdf7 	:	o_val <= 16'b0111110101110101;
                14'hdf8 	:	o_val <= 16'b0111110101110111;
                14'hdf9 	:	o_val <= 16'b0111110101111010;
                14'hdfa 	:	o_val <= 16'b0111110101111100;
                14'hdfb 	:	o_val <= 16'b0111110101111111;
                14'hdfc 	:	o_val <= 16'b0111110110000001;
                14'hdfd 	:	o_val <= 16'b0111110110000100;
                14'hdfe 	:	o_val <= 16'b0111110110000110;
                14'hdff 	:	o_val <= 16'b0111110110001001;
                14'he00 	:	o_val <= 16'b0111110110001011;
                14'he01 	:	o_val <= 16'b0111110110001110;
                14'he02 	:	o_val <= 16'b0111110110010000;
                14'he03 	:	o_val <= 16'b0111110110010010;
                14'he04 	:	o_val <= 16'b0111110110010101;
                14'he05 	:	o_val <= 16'b0111110110010111;
                14'he06 	:	o_val <= 16'b0111110110011010;
                14'he07 	:	o_val <= 16'b0111110110011100;
                14'he08 	:	o_val <= 16'b0111110110011111;
                14'he09 	:	o_val <= 16'b0111110110100001;
                14'he0a 	:	o_val <= 16'b0111110110100011;
                14'he0b 	:	o_val <= 16'b0111110110100110;
                14'he0c 	:	o_val <= 16'b0111110110101000;
                14'he0d 	:	o_val <= 16'b0111110110101011;
                14'he0e 	:	o_val <= 16'b0111110110101101;
                14'he0f 	:	o_val <= 16'b0111110110101111;
                14'he10 	:	o_val <= 16'b0111110110110010;
                14'he11 	:	o_val <= 16'b0111110110110100;
                14'he12 	:	o_val <= 16'b0111110110110110;
                14'he13 	:	o_val <= 16'b0111110110111001;
                14'he14 	:	o_val <= 16'b0111110110111011;
                14'he15 	:	o_val <= 16'b0111110110111101;
                14'he16 	:	o_val <= 16'b0111110111000000;
                14'he17 	:	o_val <= 16'b0111110111000010;
                14'he18 	:	o_val <= 16'b0111110111000101;
                14'he19 	:	o_val <= 16'b0111110111000111;
                14'he1a 	:	o_val <= 16'b0111110111001001;
                14'he1b 	:	o_val <= 16'b0111110111001100;
                14'he1c 	:	o_val <= 16'b0111110111001110;
                14'he1d 	:	o_val <= 16'b0111110111010000;
                14'he1e 	:	o_val <= 16'b0111110111010010;
                14'he1f 	:	o_val <= 16'b0111110111010101;
                14'he20 	:	o_val <= 16'b0111110111010111;
                14'he21 	:	o_val <= 16'b0111110111011001;
                14'he22 	:	o_val <= 16'b0111110111011100;
                14'he23 	:	o_val <= 16'b0111110111011110;
                14'he24 	:	o_val <= 16'b0111110111100000;
                14'he25 	:	o_val <= 16'b0111110111100010;
                14'he26 	:	o_val <= 16'b0111110111100101;
                14'he27 	:	o_val <= 16'b0111110111100111;
                14'he28 	:	o_val <= 16'b0111110111101001;
                14'he29 	:	o_val <= 16'b0111110111101100;
                14'he2a 	:	o_val <= 16'b0111110111101110;
                14'he2b 	:	o_val <= 16'b0111110111110000;
                14'he2c 	:	o_val <= 16'b0111110111110010;
                14'he2d 	:	o_val <= 16'b0111110111110101;
                14'he2e 	:	o_val <= 16'b0111110111110111;
                14'he2f 	:	o_val <= 16'b0111110111111001;
                14'he30 	:	o_val <= 16'b0111110111111011;
                14'he31 	:	o_val <= 16'b0111110111111101;
                14'he32 	:	o_val <= 16'b0111111000000000;
                14'he33 	:	o_val <= 16'b0111111000000010;
                14'he34 	:	o_val <= 16'b0111111000000100;
                14'he35 	:	o_val <= 16'b0111111000000110;
                14'he36 	:	o_val <= 16'b0111111000001000;
                14'he37 	:	o_val <= 16'b0111111000001011;
                14'he38 	:	o_val <= 16'b0111111000001101;
                14'he39 	:	o_val <= 16'b0111111000001111;
                14'he3a 	:	o_val <= 16'b0111111000010001;
                14'he3b 	:	o_val <= 16'b0111111000010011;
                14'he3c 	:	o_val <= 16'b0111111000010110;
                14'he3d 	:	o_val <= 16'b0111111000011000;
                14'he3e 	:	o_val <= 16'b0111111000011010;
                14'he3f 	:	o_val <= 16'b0111111000011100;
                14'he40 	:	o_val <= 16'b0111111000011110;
                14'he41 	:	o_val <= 16'b0111111000100000;
                14'he42 	:	o_val <= 16'b0111111000100010;
                14'he43 	:	o_val <= 16'b0111111000100101;
                14'he44 	:	o_val <= 16'b0111111000100111;
                14'he45 	:	o_val <= 16'b0111111000101001;
                14'he46 	:	o_val <= 16'b0111111000101011;
                14'he47 	:	o_val <= 16'b0111111000101101;
                14'he48 	:	o_val <= 16'b0111111000101111;
                14'he49 	:	o_val <= 16'b0111111000110001;
                14'he4a 	:	o_val <= 16'b0111111000110011;
                14'he4b 	:	o_val <= 16'b0111111000110101;
                14'he4c 	:	o_val <= 16'b0111111000111000;
                14'he4d 	:	o_val <= 16'b0111111000111010;
                14'he4e 	:	o_val <= 16'b0111111000111100;
                14'he4f 	:	o_val <= 16'b0111111000111110;
                14'he50 	:	o_val <= 16'b0111111001000000;
                14'he51 	:	o_val <= 16'b0111111001000010;
                14'he52 	:	o_val <= 16'b0111111001000100;
                14'he53 	:	o_val <= 16'b0111111001000110;
                14'he54 	:	o_val <= 16'b0111111001001000;
                14'he55 	:	o_val <= 16'b0111111001001010;
                14'he56 	:	o_val <= 16'b0111111001001100;
                14'he57 	:	o_val <= 16'b0111111001001110;
                14'he58 	:	o_val <= 16'b0111111001010000;
                14'he59 	:	o_val <= 16'b0111111001010010;
                14'he5a 	:	o_val <= 16'b0111111001010100;
                14'he5b 	:	o_val <= 16'b0111111001010110;
                14'he5c 	:	o_val <= 16'b0111111001011000;
                14'he5d 	:	o_val <= 16'b0111111001011010;
                14'he5e 	:	o_val <= 16'b0111111001011100;
                14'he5f 	:	o_val <= 16'b0111111001011110;
                14'he60 	:	o_val <= 16'b0111111001100000;
                14'he61 	:	o_val <= 16'b0111111001100010;
                14'he62 	:	o_val <= 16'b0111111001100100;
                14'he63 	:	o_val <= 16'b0111111001100110;
                14'he64 	:	o_val <= 16'b0111111001101000;
                14'he65 	:	o_val <= 16'b0111111001101010;
                14'he66 	:	o_val <= 16'b0111111001101100;
                14'he67 	:	o_val <= 16'b0111111001101110;
                14'he68 	:	o_val <= 16'b0111111001110000;
                14'he69 	:	o_val <= 16'b0111111001110010;
                14'he6a 	:	o_val <= 16'b0111111001110100;
                14'he6b 	:	o_val <= 16'b0111111001110110;
                14'he6c 	:	o_val <= 16'b0111111001111000;
                14'he6d 	:	o_val <= 16'b0111111001111010;
                14'he6e 	:	o_val <= 16'b0111111001111100;
                14'he6f 	:	o_val <= 16'b0111111001111110;
                14'he70 	:	o_val <= 16'b0111111010000000;
                14'he71 	:	o_val <= 16'b0111111010000010;
                14'he72 	:	o_val <= 16'b0111111010000100;
                14'he73 	:	o_val <= 16'b0111111010000101;
                14'he74 	:	o_val <= 16'b0111111010000111;
                14'he75 	:	o_val <= 16'b0111111010001001;
                14'he76 	:	o_val <= 16'b0111111010001011;
                14'he77 	:	o_val <= 16'b0111111010001101;
                14'he78 	:	o_val <= 16'b0111111010001111;
                14'he79 	:	o_val <= 16'b0111111010010001;
                14'he7a 	:	o_val <= 16'b0111111010010011;
                14'he7b 	:	o_val <= 16'b0111111010010100;
                14'he7c 	:	o_val <= 16'b0111111010010110;
                14'he7d 	:	o_val <= 16'b0111111010011000;
                14'he7e 	:	o_val <= 16'b0111111010011010;
                14'he7f 	:	o_val <= 16'b0111111010011100;
                14'he80 	:	o_val <= 16'b0111111010011110;
                14'he81 	:	o_val <= 16'b0111111010100000;
                14'he82 	:	o_val <= 16'b0111111010100001;
                14'he83 	:	o_val <= 16'b0111111010100011;
                14'he84 	:	o_val <= 16'b0111111010100101;
                14'he85 	:	o_val <= 16'b0111111010100111;
                14'he86 	:	o_val <= 16'b0111111010101001;
                14'he87 	:	o_val <= 16'b0111111010101011;
                14'he88 	:	o_val <= 16'b0111111010101100;
                14'he89 	:	o_val <= 16'b0111111010101110;
                14'he8a 	:	o_val <= 16'b0111111010110000;
                14'he8b 	:	o_val <= 16'b0111111010110010;
                14'he8c 	:	o_val <= 16'b0111111010110100;
                14'he8d 	:	o_val <= 16'b0111111010110101;
                14'he8e 	:	o_val <= 16'b0111111010110111;
                14'he8f 	:	o_val <= 16'b0111111010111001;
                14'he90 	:	o_val <= 16'b0111111010111011;
                14'he91 	:	o_val <= 16'b0111111010111100;
                14'he92 	:	o_val <= 16'b0111111010111110;
                14'he93 	:	o_val <= 16'b0111111011000000;
                14'he94 	:	o_val <= 16'b0111111011000010;
                14'he95 	:	o_val <= 16'b0111111011000011;
                14'he96 	:	o_val <= 16'b0111111011000101;
                14'he97 	:	o_val <= 16'b0111111011000111;
                14'he98 	:	o_val <= 16'b0111111011001001;
                14'he99 	:	o_val <= 16'b0111111011001010;
                14'he9a 	:	o_val <= 16'b0111111011001100;
                14'he9b 	:	o_val <= 16'b0111111011001110;
                14'he9c 	:	o_val <= 16'b0111111011001111;
                14'he9d 	:	o_val <= 16'b0111111011010001;
                14'he9e 	:	o_val <= 16'b0111111011010011;
                14'he9f 	:	o_val <= 16'b0111111011010101;
                14'hea0 	:	o_val <= 16'b0111111011010110;
                14'hea1 	:	o_val <= 16'b0111111011011000;
                14'hea2 	:	o_val <= 16'b0111111011011010;
                14'hea3 	:	o_val <= 16'b0111111011011011;
                14'hea4 	:	o_val <= 16'b0111111011011101;
                14'hea5 	:	o_val <= 16'b0111111011011111;
                14'hea6 	:	o_val <= 16'b0111111011100000;
                14'hea7 	:	o_val <= 16'b0111111011100010;
                14'hea8 	:	o_val <= 16'b0111111011100100;
                14'hea9 	:	o_val <= 16'b0111111011100101;
                14'heaa 	:	o_val <= 16'b0111111011100111;
                14'heab 	:	o_val <= 16'b0111111011101001;
                14'heac 	:	o_val <= 16'b0111111011101010;
                14'head 	:	o_val <= 16'b0111111011101100;
                14'heae 	:	o_val <= 16'b0111111011101101;
                14'heaf 	:	o_val <= 16'b0111111011101111;
                14'heb0 	:	o_val <= 16'b0111111011110001;
                14'heb1 	:	o_val <= 16'b0111111011110010;
                14'heb2 	:	o_val <= 16'b0111111011110100;
                14'heb3 	:	o_val <= 16'b0111111011110101;
                14'heb4 	:	o_val <= 16'b0111111011110111;
                14'heb5 	:	o_val <= 16'b0111111011111001;
                14'heb6 	:	o_val <= 16'b0111111011111010;
                14'heb7 	:	o_val <= 16'b0111111011111100;
                14'heb8 	:	o_val <= 16'b0111111011111101;
                14'heb9 	:	o_val <= 16'b0111111011111111;
                14'heba 	:	o_val <= 16'b0111111100000001;
                14'hebb 	:	o_val <= 16'b0111111100000010;
                14'hebc 	:	o_val <= 16'b0111111100000100;
                14'hebd 	:	o_val <= 16'b0111111100000101;
                14'hebe 	:	o_val <= 16'b0111111100000111;
                14'hebf 	:	o_val <= 16'b0111111100001000;
                14'hec0 	:	o_val <= 16'b0111111100001010;
                14'hec1 	:	o_val <= 16'b0111111100001011;
                14'hec2 	:	o_val <= 16'b0111111100001101;
                14'hec3 	:	o_val <= 16'b0111111100001110;
                14'hec4 	:	o_val <= 16'b0111111100010000;
                14'hec5 	:	o_val <= 16'b0111111100010001;
                14'hec6 	:	o_val <= 16'b0111111100010011;
                14'hec7 	:	o_val <= 16'b0111111100010100;
                14'hec8 	:	o_val <= 16'b0111111100010110;
                14'hec9 	:	o_val <= 16'b0111111100010111;
                14'heca 	:	o_val <= 16'b0111111100011001;
                14'hecb 	:	o_val <= 16'b0111111100011010;
                14'hecc 	:	o_val <= 16'b0111111100011100;
                14'hecd 	:	o_val <= 16'b0111111100011101;
                14'hece 	:	o_val <= 16'b0111111100011111;
                14'hecf 	:	o_val <= 16'b0111111100100000;
                14'hed0 	:	o_val <= 16'b0111111100100010;
                14'hed1 	:	o_val <= 16'b0111111100100011;
                14'hed2 	:	o_val <= 16'b0111111100100101;
                14'hed3 	:	o_val <= 16'b0111111100100110;
                14'hed4 	:	o_val <= 16'b0111111100101000;
                14'hed5 	:	o_val <= 16'b0111111100101001;
                14'hed6 	:	o_val <= 16'b0111111100101010;
                14'hed7 	:	o_val <= 16'b0111111100101100;
                14'hed8 	:	o_val <= 16'b0111111100101101;
                14'hed9 	:	o_val <= 16'b0111111100101111;
                14'heda 	:	o_val <= 16'b0111111100110000;
                14'hedb 	:	o_val <= 16'b0111111100110010;
                14'hedc 	:	o_val <= 16'b0111111100110011;
                14'hedd 	:	o_val <= 16'b0111111100110100;
                14'hede 	:	o_val <= 16'b0111111100110110;
                14'hedf 	:	o_val <= 16'b0111111100110111;
                14'hee0 	:	o_val <= 16'b0111111100111001;
                14'hee1 	:	o_val <= 16'b0111111100111010;
                14'hee2 	:	o_val <= 16'b0111111100111011;
                14'hee3 	:	o_val <= 16'b0111111100111101;
                14'hee4 	:	o_val <= 16'b0111111100111110;
                14'hee5 	:	o_val <= 16'b0111111100111111;
                14'hee6 	:	o_val <= 16'b0111111101000001;
                14'hee7 	:	o_val <= 16'b0111111101000010;
                14'hee8 	:	o_val <= 16'b0111111101000011;
                14'hee9 	:	o_val <= 16'b0111111101000101;
                14'heea 	:	o_val <= 16'b0111111101000110;
                14'heeb 	:	o_val <= 16'b0111111101000111;
                14'heec 	:	o_val <= 16'b0111111101001001;
                14'heed 	:	o_val <= 16'b0111111101001010;
                14'heee 	:	o_val <= 16'b0111111101001011;
                14'heef 	:	o_val <= 16'b0111111101001101;
                14'hef0 	:	o_val <= 16'b0111111101001110;
                14'hef1 	:	o_val <= 16'b0111111101001111;
                14'hef2 	:	o_val <= 16'b0111111101010001;
                14'hef3 	:	o_val <= 16'b0111111101010010;
                14'hef4 	:	o_val <= 16'b0111111101010011;
                14'hef5 	:	o_val <= 16'b0111111101010101;
                14'hef6 	:	o_val <= 16'b0111111101010110;
                14'hef7 	:	o_val <= 16'b0111111101010111;
                14'hef8 	:	o_val <= 16'b0111111101011000;
                14'hef9 	:	o_val <= 16'b0111111101011010;
                14'hefa 	:	o_val <= 16'b0111111101011011;
                14'hefb 	:	o_val <= 16'b0111111101011100;
                14'hefc 	:	o_val <= 16'b0111111101011101;
                14'hefd 	:	o_val <= 16'b0111111101011111;
                14'hefe 	:	o_val <= 16'b0111111101100000;
                14'heff 	:	o_val <= 16'b0111111101100001;
                14'hf00 	:	o_val <= 16'b0111111101100010;
                14'hf01 	:	o_val <= 16'b0111111101100100;
                14'hf02 	:	o_val <= 16'b0111111101100101;
                14'hf03 	:	o_val <= 16'b0111111101100110;
                14'hf04 	:	o_val <= 16'b0111111101100111;
                14'hf05 	:	o_val <= 16'b0111111101101000;
                14'hf06 	:	o_val <= 16'b0111111101101010;
                14'hf07 	:	o_val <= 16'b0111111101101011;
                14'hf08 	:	o_val <= 16'b0111111101101100;
                14'hf09 	:	o_val <= 16'b0111111101101101;
                14'hf0a 	:	o_val <= 16'b0111111101101110;
                14'hf0b 	:	o_val <= 16'b0111111101110000;
                14'hf0c 	:	o_val <= 16'b0111111101110001;
                14'hf0d 	:	o_val <= 16'b0111111101110010;
                14'hf0e 	:	o_val <= 16'b0111111101110011;
                14'hf0f 	:	o_val <= 16'b0111111101110100;
                14'hf10 	:	o_val <= 16'b0111111101110101;
                14'hf11 	:	o_val <= 16'b0111111101110111;
                14'hf12 	:	o_val <= 16'b0111111101111000;
                14'hf13 	:	o_val <= 16'b0111111101111001;
                14'hf14 	:	o_val <= 16'b0111111101111010;
                14'hf15 	:	o_val <= 16'b0111111101111011;
                14'hf16 	:	o_val <= 16'b0111111101111100;
                14'hf17 	:	o_val <= 16'b0111111101111101;
                14'hf18 	:	o_val <= 16'b0111111101111110;
                14'hf19 	:	o_val <= 16'b0111111110000000;
                14'hf1a 	:	o_val <= 16'b0111111110000001;
                14'hf1b 	:	o_val <= 16'b0111111110000010;
                14'hf1c 	:	o_val <= 16'b0111111110000011;
                14'hf1d 	:	o_val <= 16'b0111111110000100;
                14'hf1e 	:	o_val <= 16'b0111111110000101;
                14'hf1f 	:	o_val <= 16'b0111111110000110;
                14'hf20 	:	o_val <= 16'b0111111110000111;
                14'hf21 	:	o_val <= 16'b0111111110001000;
                14'hf22 	:	o_val <= 16'b0111111110001001;
                14'hf23 	:	o_val <= 16'b0111111110001010;
                14'hf24 	:	o_val <= 16'b0111111110001011;
                14'hf25 	:	o_val <= 16'b0111111110001101;
                14'hf26 	:	o_val <= 16'b0111111110001110;
                14'hf27 	:	o_val <= 16'b0111111110001111;
                14'hf28 	:	o_val <= 16'b0111111110010000;
                14'hf29 	:	o_val <= 16'b0111111110010001;
                14'hf2a 	:	o_val <= 16'b0111111110010010;
                14'hf2b 	:	o_val <= 16'b0111111110010011;
                14'hf2c 	:	o_val <= 16'b0111111110010100;
                14'hf2d 	:	o_val <= 16'b0111111110010101;
                14'hf2e 	:	o_val <= 16'b0111111110010110;
                14'hf2f 	:	o_val <= 16'b0111111110010111;
                14'hf30 	:	o_val <= 16'b0111111110011000;
                14'hf31 	:	o_val <= 16'b0111111110011001;
                14'hf32 	:	o_val <= 16'b0111111110011010;
                14'hf33 	:	o_val <= 16'b0111111110011011;
                14'hf34 	:	o_val <= 16'b0111111110011100;
                14'hf35 	:	o_val <= 16'b0111111110011101;
                14'hf36 	:	o_val <= 16'b0111111110011110;
                14'hf37 	:	o_val <= 16'b0111111110011111;
                14'hf38 	:	o_val <= 16'b0111111110100000;
                14'hf39 	:	o_val <= 16'b0111111110100001;
                14'hf3a 	:	o_val <= 16'b0111111110100010;
                14'hf3b 	:	o_val <= 16'b0111111110100011;
                14'hf3c 	:	o_val <= 16'b0111111110100011;
                14'hf3d 	:	o_val <= 16'b0111111110100100;
                14'hf3e 	:	o_val <= 16'b0111111110100101;
                14'hf3f 	:	o_val <= 16'b0111111110100110;
                14'hf40 	:	o_val <= 16'b0111111110100111;
                14'hf41 	:	o_val <= 16'b0111111110101000;
                14'hf42 	:	o_val <= 16'b0111111110101001;
                14'hf43 	:	o_val <= 16'b0111111110101010;
                14'hf44 	:	o_val <= 16'b0111111110101011;
                14'hf45 	:	o_val <= 16'b0111111110101100;
                14'hf46 	:	o_val <= 16'b0111111110101101;
                14'hf47 	:	o_val <= 16'b0111111110101110;
                14'hf48 	:	o_val <= 16'b0111111110101110;
                14'hf49 	:	o_val <= 16'b0111111110101111;
                14'hf4a 	:	o_val <= 16'b0111111110110000;
                14'hf4b 	:	o_val <= 16'b0111111110110001;
                14'hf4c 	:	o_val <= 16'b0111111110110010;
                14'hf4d 	:	o_val <= 16'b0111111110110011;
                14'hf4e 	:	o_val <= 16'b0111111110110100;
                14'hf4f 	:	o_val <= 16'b0111111110110100;
                14'hf50 	:	o_val <= 16'b0111111110110101;
                14'hf51 	:	o_val <= 16'b0111111110110110;
                14'hf52 	:	o_val <= 16'b0111111110110111;
                14'hf53 	:	o_val <= 16'b0111111110111000;
                14'hf54 	:	o_val <= 16'b0111111110111001;
                14'hf55 	:	o_val <= 16'b0111111110111001;
                14'hf56 	:	o_val <= 16'b0111111110111010;
                14'hf57 	:	o_val <= 16'b0111111110111011;
                14'hf58 	:	o_val <= 16'b0111111110111100;
                14'hf59 	:	o_val <= 16'b0111111110111101;
                14'hf5a 	:	o_val <= 16'b0111111110111110;
                14'hf5b 	:	o_val <= 16'b0111111110111110;
                14'hf5c 	:	o_val <= 16'b0111111110111111;
                14'hf5d 	:	o_val <= 16'b0111111111000000;
                14'hf5e 	:	o_val <= 16'b0111111111000001;
                14'hf5f 	:	o_val <= 16'b0111111111000001;
                14'hf60 	:	o_val <= 16'b0111111111000010;
                14'hf61 	:	o_val <= 16'b0111111111000011;
                14'hf62 	:	o_val <= 16'b0111111111000100;
                14'hf63 	:	o_val <= 16'b0111111111000101;
                14'hf64 	:	o_val <= 16'b0111111111000101;
                14'hf65 	:	o_val <= 16'b0111111111000110;
                14'hf66 	:	o_val <= 16'b0111111111000111;
                14'hf67 	:	o_val <= 16'b0111111111000111;
                14'hf68 	:	o_val <= 16'b0111111111001000;
                14'hf69 	:	o_val <= 16'b0111111111001001;
                14'hf6a 	:	o_val <= 16'b0111111111001010;
                14'hf6b 	:	o_val <= 16'b0111111111001010;
                14'hf6c 	:	o_val <= 16'b0111111111001011;
                14'hf6d 	:	o_val <= 16'b0111111111001100;
                14'hf6e 	:	o_val <= 16'b0111111111001101;
                14'hf6f 	:	o_val <= 16'b0111111111001101;
                14'hf70 	:	o_val <= 16'b0111111111001110;
                14'hf71 	:	o_val <= 16'b0111111111001111;
                14'hf72 	:	o_val <= 16'b0111111111001111;
                14'hf73 	:	o_val <= 16'b0111111111010000;
                14'hf74 	:	o_val <= 16'b0111111111010001;
                14'hf75 	:	o_val <= 16'b0111111111010001;
                14'hf76 	:	o_val <= 16'b0111111111010010;
                14'hf77 	:	o_val <= 16'b0111111111010011;
                14'hf78 	:	o_val <= 16'b0111111111010011;
                14'hf79 	:	o_val <= 16'b0111111111010100;
                14'hf7a 	:	o_val <= 16'b0111111111010101;
                14'hf7b 	:	o_val <= 16'b0111111111010101;
                14'hf7c 	:	o_val <= 16'b0111111111010110;
                14'hf7d 	:	o_val <= 16'b0111111111010110;
                14'hf7e 	:	o_val <= 16'b0111111111010111;
                14'hf7f 	:	o_val <= 16'b0111111111011000;
                14'hf80 	:	o_val <= 16'b0111111111011000;
                14'hf81 	:	o_val <= 16'b0111111111011001;
                14'hf82 	:	o_val <= 16'b0111111111011010;
                14'hf83 	:	o_val <= 16'b0111111111011010;
                14'hf84 	:	o_val <= 16'b0111111111011011;
                14'hf85 	:	o_val <= 16'b0111111111011011;
                14'hf86 	:	o_val <= 16'b0111111111011100;
                14'hf87 	:	o_val <= 16'b0111111111011101;
                14'hf88 	:	o_val <= 16'b0111111111011101;
                14'hf89 	:	o_val <= 16'b0111111111011110;
                14'hf8a 	:	o_val <= 16'b0111111111011110;
                14'hf8b 	:	o_val <= 16'b0111111111011111;
                14'hf8c 	:	o_val <= 16'b0111111111011111;
                14'hf8d 	:	o_val <= 16'b0111111111100000;
                14'hf8e 	:	o_val <= 16'b0111111111100000;
                14'hf8f 	:	o_val <= 16'b0111111111100001;
                14'hf90 	:	o_val <= 16'b0111111111100010;
                14'hf91 	:	o_val <= 16'b0111111111100010;
                14'hf92 	:	o_val <= 16'b0111111111100011;
                14'hf93 	:	o_val <= 16'b0111111111100011;
                14'hf94 	:	o_val <= 16'b0111111111100100;
                14'hf95 	:	o_val <= 16'b0111111111100100;
                14'hf96 	:	o_val <= 16'b0111111111100101;
                14'hf97 	:	o_val <= 16'b0111111111100101;
                14'hf98 	:	o_val <= 16'b0111111111100110;
                14'hf99 	:	o_val <= 16'b0111111111100110;
                14'hf9a 	:	o_val <= 16'b0111111111100111;
                14'hf9b 	:	o_val <= 16'b0111111111100111;
                14'hf9c 	:	o_val <= 16'b0111111111101000;
                14'hf9d 	:	o_val <= 16'b0111111111101000;
                14'hf9e 	:	o_val <= 16'b0111111111101001;
                14'hf9f 	:	o_val <= 16'b0111111111101001;
                14'hfa0 	:	o_val <= 16'b0111111111101010;
                14'hfa1 	:	o_val <= 16'b0111111111101010;
                14'hfa2 	:	o_val <= 16'b0111111111101010;
                14'hfa3 	:	o_val <= 16'b0111111111101011;
                14'hfa4 	:	o_val <= 16'b0111111111101011;
                14'hfa5 	:	o_val <= 16'b0111111111101100;
                14'hfa6 	:	o_val <= 16'b0111111111101100;
                14'hfa7 	:	o_val <= 16'b0111111111101101;
                14'hfa8 	:	o_val <= 16'b0111111111101101;
                14'hfa9 	:	o_val <= 16'b0111111111101101;
                14'hfaa 	:	o_val <= 16'b0111111111101110;
                14'hfab 	:	o_val <= 16'b0111111111101110;
                14'hfac 	:	o_val <= 16'b0111111111101111;
                14'hfad 	:	o_val <= 16'b0111111111101111;
                14'hfae 	:	o_val <= 16'b0111111111101111;
                14'hfaf 	:	o_val <= 16'b0111111111110000;
                14'hfb0 	:	o_val <= 16'b0111111111110000;
                14'hfb1 	:	o_val <= 16'b0111111111110001;
                14'hfb2 	:	o_val <= 16'b0111111111110001;
                14'hfb3 	:	o_val <= 16'b0111111111110001;
                14'hfb4 	:	o_val <= 16'b0111111111110010;
                14'hfb5 	:	o_val <= 16'b0111111111110010;
                14'hfb6 	:	o_val <= 16'b0111111111110010;
                14'hfb7 	:	o_val <= 16'b0111111111110011;
                14'hfb8 	:	o_val <= 16'b0111111111110011;
                14'hfb9 	:	o_val <= 16'b0111111111110100;
                14'hfba 	:	o_val <= 16'b0111111111110100;
                14'hfbb 	:	o_val <= 16'b0111111111110100;
                14'hfbc 	:	o_val <= 16'b0111111111110101;
                14'hfbd 	:	o_val <= 16'b0111111111110101;
                14'hfbe 	:	o_val <= 16'b0111111111110101;
                14'hfbf 	:	o_val <= 16'b0111111111110101;
                14'hfc0 	:	o_val <= 16'b0111111111110110;
                14'hfc1 	:	o_val <= 16'b0111111111110110;
                14'hfc2 	:	o_val <= 16'b0111111111110110;
                14'hfc3 	:	o_val <= 16'b0111111111110111;
                14'hfc4 	:	o_val <= 16'b0111111111110111;
                14'hfc5 	:	o_val <= 16'b0111111111110111;
                14'hfc6 	:	o_val <= 16'b0111111111111000;
                14'hfc7 	:	o_val <= 16'b0111111111111000;
                14'hfc8 	:	o_val <= 16'b0111111111111000;
                14'hfc9 	:	o_val <= 16'b0111111111111000;
                14'hfca 	:	o_val <= 16'b0111111111111001;
                14'hfcb 	:	o_val <= 16'b0111111111111001;
                14'hfcc 	:	o_val <= 16'b0111111111111001;
                14'hfcd 	:	o_val <= 16'b0111111111111001;
                14'hfce 	:	o_val <= 16'b0111111111111010;
                14'hfcf 	:	o_val <= 16'b0111111111111010;
                14'hfd0 	:	o_val <= 16'b0111111111111010;
                14'hfd1 	:	o_val <= 16'b0111111111111010;
                14'hfd2 	:	o_val <= 16'b0111111111111011;
                14'hfd3 	:	o_val <= 16'b0111111111111011;
                14'hfd4 	:	o_val <= 16'b0111111111111011;
                14'hfd5 	:	o_val <= 16'b0111111111111011;
                14'hfd6 	:	o_val <= 16'b0111111111111011;
                14'hfd7 	:	o_val <= 16'b0111111111111100;
                14'hfd8 	:	o_val <= 16'b0111111111111100;
                14'hfd9 	:	o_val <= 16'b0111111111111100;
                14'hfda 	:	o_val <= 16'b0111111111111100;
                14'hfdb 	:	o_val <= 16'b0111111111111100;
                14'hfdc 	:	o_val <= 16'b0111111111111100;
                14'hfdd 	:	o_val <= 16'b0111111111111101;
                14'hfde 	:	o_val <= 16'b0111111111111101;
                14'hfdf 	:	o_val <= 16'b0111111111111101;
                14'hfe0 	:	o_val <= 16'b0111111111111101;
                14'hfe1 	:	o_val <= 16'b0111111111111101;
                14'hfe2 	:	o_val <= 16'b0111111111111101;
                14'hfe3 	:	o_val <= 16'b0111111111111110;
                14'hfe4 	:	o_val <= 16'b0111111111111110;
                14'hfe5 	:	o_val <= 16'b0111111111111110;
                14'hfe6 	:	o_val <= 16'b0111111111111110;
                14'hfe7 	:	o_val <= 16'b0111111111111110;
                14'hfe8 	:	o_val <= 16'b0111111111111110;
                14'hfe9 	:	o_val <= 16'b0111111111111110;
                14'hfea 	:	o_val <= 16'b0111111111111110;
                14'hfeb 	:	o_val <= 16'b0111111111111110;
                14'hfec 	:	o_val <= 16'b0111111111111111;
                14'hfed 	:	o_val <= 16'b0111111111111111;
                14'hfee 	:	o_val <= 16'b0111111111111111;
                14'hfef 	:	o_val <= 16'b0111111111111111;
                14'hff0 	:	o_val <= 16'b0111111111111111;
                14'hff1 	:	o_val <= 16'b0111111111111111;
                14'hff2 	:	o_val <= 16'b0111111111111111;
                14'hff3 	:	o_val <= 16'b0111111111111111;
                14'hff4 	:	o_val <= 16'b0111111111111111;
                14'hff5 	:	o_val <= 16'b0111111111111111;
                14'hff6 	:	o_val <= 16'b0111111111111111;
                14'hff7 	:	o_val <= 16'b0111111111111111;
                14'hff8 	:	o_val <= 16'b0111111111111111;
                14'hff9 	:	o_val <= 16'b0111111111111111;
                14'hffa 	:	o_val <= 16'b0111111111111111;
                14'hffb 	:	o_val <= 16'b0111111111111111;
                14'hffc 	:	o_val <= 16'b0111111111111111;
                14'hffd 	:	o_val <= 16'b0111111111111111;
                14'hffe 	:	o_val <= 16'b0111111111111111;
                14'hfff 	:	o_val <= 16'b0111111111111111;
				 default		:	o_val <= 16'b0;
			endcase
		end
endmodule
                                        
