module sawtooth_lut(input[9:0] i_phase,
								output reg signed[15:0] o_val);
        initial o_val = 16'b0;

		always @(i_phase) begin
			case(i_phase)
            10'h000 	:	o_val <= 16'b0000000000000000;
            10'h001 	:	o_val <= 16'b0000000000100000;
            10'h002 	:	o_val <= 16'b0000000001000000;
            10'h003 	:	o_val <= 16'b0000000001100000;
            10'h004 	:	o_val <= 16'b0000000010000000;
            10'h005 	:	o_val <= 16'b0000000010100000;
            10'h006 	:	o_val <= 16'b0000000011000000;
            10'h007 	:	o_val <= 16'b0000000011100000;
            10'h008 	:	o_val <= 16'b0000000100000000;
            10'h009 	:	o_val <= 16'b0000000100100000;
            10'h00a 	:	o_val <= 16'b0000000101000000;
            10'h00b 	:	o_val <= 16'b0000000101100000;
            10'h00c 	:	o_val <= 16'b0000000110000000;
            10'h00d 	:	o_val <= 16'b0000000110100000;
            10'h00e 	:	o_val <= 16'b0000000111000000;
            10'h00f 	:	o_val <= 16'b0000000111100000;
            10'h010 	:	o_val <= 16'b0000001000000000;
            10'h011 	:	o_val <= 16'b0000001000100000;
            10'h012 	:	o_val <= 16'b0000001001000000;
            10'h013 	:	o_val <= 16'b0000001001100000;
            10'h014 	:	o_val <= 16'b0000001010000000;
            10'h015 	:	o_val <= 16'b0000001010100000;
            10'h016 	:	o_val <= 16'b0000001011000000;
            10'h017 	:	o_val <= 16'b0000001011100000;
            10'h018 	:	o_val <= 16'b0000001100000000;
            10'h019 	:	o_val <= 16'b0000001100100000;
            10'h01a 	:	o_val <= 16'b0000001101000000;
            10'h01b 	:	o_val <= 16'b0000001101100000;
            10'h01c 	:	o_val <= 16'b0000001110000000;
            10'h01d 	:	o_val <= 16'b0000001110100000;
            10'h01e 	:	o_val <= 16'b0000001111000000;
            10'h01f 	:	o_val <= 16'b0000001111100000;
            10'h020 	:	o_val <= 16'b0000010000000000;
            10'h021 	:	o_val <= 16'b0000010000100000;
            10'h022 	:	o_val <= 16'b0000010001000000;
            10'h023 	:	o_val <= 16'b0000010001100000;
            10'h024 	:	o_val <= 16'b0000010010000000;
            10'h025 	:	o_val <= 16'b0000010010100000;
            10'h026 	:	o_val <= 16'b0000010011000000;
            10'h027 	:	o_val <= 16'b0000010011100000;
            10'h028 	:	o_val <= 16'b0000010100000000;
            10'h029 	:	o_val <= 16'b0000010100100000;
            10'h02a 	:	o_val <= 16'b0000010101000000;
            10'h02b 	:	o_val <= 16'b0000010101100000;
            10'h02c 	:	o_val <= 16'b0000010110000000;
            10'h02d 	:	o_val <= 16'b0000010110100000;
            10'h02e 	:	o_val <= 16'b0000010111000000;
            10'h02f 	:	o_val <= 16'b0000010111100000;
            10'h030 	:	o_val <= 16'b0000011000000000;
            10'h031 	:	o_val <= 16'b0000011000100000;
            10'h032 	:	o_val <= 16'b0000011001000000;
            10'h033 	:	o_val <= 16'b0000011001100000;
            10'h034 	:	o_val <= 16'b0000011010000000;
            10'h035 	:	o_val <= 16'b0000011010100000;
            10'h036 	:	o_val <= 16'b0000011011000000;
            10'h037 	:	o_val <= 16'b0000011011100000;
            10'h038 	:	o_val <= 16'b0000011100000000;
            10'h039 	:	o_val <= 16'b0000011100100000;
            10'h03a 	:	o_val <= 16'b0000011101000000;
            10'h03b 	:	o_val <= 16'b0000011101100000;
            10'h03c 	:	o_val <= 16'b0000011110000000;
            10'h03d 	:	o_val <= 16'b0000011110100000;
            10'h03e 	:	o_val <= 16'b0000011111000000;
            10'h03f 	:	o_val <= 16'b0000011111100000;
            10'h040 	:	o_val <= 16'b0000100000000000;
            10'h041 	:	o_val <= 16'b0000100000100000;
            10'h042 	:	o_val <= 16'b0000100001000000;
            10'h043 	:	o_val <= 16'b0000100001100000;
            10'h044 	:	o_val <= 16'b0000100010000000;
            10'h045 	:	o_val <= 16'b0000100010100000;
            10'h046 	:	o_val <= 16'b0000100011000000;
            10'h047 	:	o_val <= 16'b0000100011100000;
            10'h048 	:	o_val <= 16'b0000100100000000;
            10'h049 	:	o_val <= 16'b0000100100100000;
            10'h04a 	:	o_val <= 16'b0000100101000000;
            10'h04b 	:	o_val <= 16'b0000100101100000;
            10'h04c 	:	o_val <= 16'b0000100110000000;
            10'h04d 	:	o_val <= 16'b0000100110100000;
            10'h04e 	:	o_val <= 16'b0000100111000000;
            10'h04f 	:	o_val <= 16'b0000100111100000;
            10'h050 	:	o_val <= 16'b0000101000000000;
            10'h051 	:	o_val <= 16'b0000101000100000;
            10'h052 	:	o_val <= 16'b0000101001000000;
            10'h053 	:	o_val <= 16'b0000101001100000;
            10'h054 	:	o_val <= 16'b0000101010000000;
            10'h055 	:	o_val <= 16'b0000101010100000;
            10'h056 	:	o_val <= 16'b0000101011000000;
            10'h057 	:	o_val <= 16'b0000101011100000;
            10'h058 	:	o_val <= 16'b0000101100000000;
            10'h059 	:	o_val <= 16'b0000101100100000;
            10'h05a 	:	o_val <= 16'b0000101101000000;
            10'h05b 	:	o_val <= 16'b0000101101100000;
            10'h05c 	:	o_val <= 16'b0000101110000000;
            10'h05d 	:	o_val <= 16'b0000101110100000;
            10'h05e 	:	o_val <= 16'b0000101111000000;
            10'h05f 	:	o_val <= 16'b0000101111100000;
            10'h060 	:	o_val <= 16'b0000110000000000;
            10'h061 	:	o_val <= 16'b0000110000100000;
            10'h062 	:	o_val <= 16'b0000110001000000;
            10'h063 	:	o_val <= 16'b0000110001100000;
            10'h064 	:	o_val <= 16'b0000110010000000;
            10'h065 	:	o_val <= 16'b0000110010100000;
            10'h066 	:	o_val <= 16'b0000110011000000;
            10'h067 	:	o_val <= 16'b0000110011100000;
            10'h068 	:	o_val <= 16'b0000110100000000;
            10'h069 	:	o_val <= 16'b0000110100100000;
            10'h06a 	:	o_val <= 16'b0000110101000000;
            10'h06b 	:	o_val <= 16'b0000110101100000;
            10'h06c 	:	o_val <= 16'b0000110110000000;
            10'h06d 	:	o_val <= 16'b0000110110100000;
            10'h06e 	:	o_val <= 16'b0000110111000000;
            10'h06f 	:	o_val <= 16'b0000110111100000;
            10'h070 	:	o_val <= 16'b0000111000000000;
            10'h071 	:	o_val <= 16'b0000111000100000;
            10'h072 	:	o_val <= 16'b0000111001000000;
            10'h073 	:	o_val <= 16'b0000111001100000;
            10'h074 	:	o_val <= 16'b0000111010000000;
            10'h075 	:	o_val <= 16'b0000111010100000;
            10'h076 	:	o_val <= 16'b0000111011000000;
            10'h077 	:	o_val <= 16'b0000111011100000;
            10'h078 	:	o_val <= 16'b0000111100000000;
            10'h079 	:	o_val <= 16'b0000111100100000;
            10'h07a 	:	o_val <= 16'b0000111101000000;
            10'h07b 	:	o_val <= 16'b0000111101100000;
            10'h07c 	:	o_val <= 16'b0000111110000000;
            10'h07d 	:	o_val <= 16'b0000111110100000;
            10'h07e 	:	o_val <= 16'b0000111111000000;
            10'h07f 	:	o_val <= 16'b0000111111100000;
            10'h080 	:	o_val <= 16'b0001000000000000;
            10'h081 	:	o_val <= 16'b0001000000100000;
            10'h082 	:	o_val <= 16'b0001000001000000;
            10'h083 	:	o_val <= 16'b0001000001100000;
            10'h084 	:	o_val <= 16'b0001000010000000;
            10'h085 	:	o_val <= 16'b0001000010100000;
            10'h086 	:	o_val <= 16'b0001000011000000;
            10'h087 	:	o_val <= 16'b0001000011100000;
            10'h088 	:	o_val <= 16'b0001000100000000;
            10'h089 	:	o_val <= 16'b0001000100100000;
            10'h08a 	:	o_val <= 16'b0001000101000000;
            10'h08b 	:	o_val <= 16'b0001000101100000;
            10'h08c 	:	o_val <= 16'b0001000110000000;
            10'h08d 	:	o_val <= 16'b0001000110100000;
            10'h08e 	:	o_val <= 16'b0001000111000000;
            10'h08f 	:	o_val <= 16'b0001000111100000;
            10'h090 	:	o_val <= 16'b0001001000000000;
            10'h091 	:	o_val <= 16'b0001001000100000;
            10'h092 	:	o_val <= 16'b0001001001000000;
            10'h093 	:	o_val <= 16'b0001001001100000;
            10'h094 	:	o_val <= 16'b0001001010000000;
            10'h095 	:	o_val <= 16'b0001001010100000;
            10'h096 	:	o_val <= 16'b0001001011000000;
            10'h097 	:	o_val <= 16'b0001001011100000;
            10'h098 	:	o_val <= 16'b0001001100000000;
            10'h099 	:	o_val <= 16'b0001001100100000;
            10'h09a 	:	o_val <= 16'b0001001101000000;
            10'h09b 	:	o_val <= 16'b0001001101100000;
            10'h09c 	:	o_val <= 16'b0001001110000000;
            10'h09d 	:	o_val <= 16'b0001001110100000;
            10'h09e 	:	o_val <= 16'b0001001111000000;
            10'h09f 	:	o_val <= 16'b0001001111100000;
            10'h0a0 	:	o_val <= 16'b0001010000000000;
            10'h0a1 	:	o_val <= 16'b0001010000100000;
            10'h0a2 	:	o_val <= 16'b0001010001000000;
            10'h0a3 	:	o_val <= 16'b0001010001100000;
            10'h0a4 	:	o_val <= 16'b0001010010000000;
            10'h0a5 	:	o_val <= 16'b0001010010100000;
            10'h0a6 	:	o_val <= 16'b0001010011000000;
            10'h0a7 	:	o_val <= 16'b0001010011100000;
            10'h0a8 	:	o_val <= 16'b0001010100000000;
            10'h0a9 	:	o_val <= 16'b0001010100100000;
            10'h0aa 	:	o_val <= 16'b0001010101000000;
            10'h0ab 	:	o_val <= 16'b0001010101100000;
            10'h0ac 	:	o_val <= 16'b0001010110000000;
            10'h0ad 	:	o_val <= 16'b0001010110100000;
            10'h0ae 	:	o_val <= 16'b0001010111000000;
            10'h0af 	:	o_val <= 16'b0001010111100000;
            10'h0b0 	:	o_val <= 16'b0001011000000000;
            10'h0b1 	:	o_val <= 16'b0001011000100000;
            10'h0b2 	:	o_val <= 16'b0001011001000000;
            10'h0b3 	:	o_val <= 16'b0001011001100000;
            10'h0b4 	:	o_val <= 16'b0001011010000000;
            10'h0b5 	:	o_val <= 16'b0001011010100000;
            10'h0b6 	:	o_val <= 16'b0001011011000000;
            10'h0b7 	:	o_val <= 16'b0001011011100000;
            10'h0b8 	:	o_val <= 16'b0001011100000000;
            10'h0b9 	:	o_val <= 16'b0001011100100000;
            10'h0ba 	:	o_val <= 16'b0001011101000000;
            10'h0bb 	:	o_val <= 16'b0001011101100000;
            10'h0bc 	:	o_val <= 16'b0001011110000000;
            10'h0bd 	:	o_val <= 16'b0001011110100000;
            10'h0be 	:	o_val <= 16'b0001011111000000;
            10'h0bf 	:	o_val <= 16'b0001011111100000;
            10'h0c0 	:	o_val <= 16'b0001100000000000;
            10'h0c1 	:	o_val <= 16'b0001100000100000;
            10'h0c2 	:	o_val <= 16'b0001100001000000;
            10'h0c3 	:	o_val <= 16'b0001100001100000;
            10'h0c4 	:	o_val <= 16'b0001100010000000;
            10'h0c5 	:	o_val <= 16'b0001100010100000;
            10'h0c6 	:	o_val <= 16'b0001100011000000;
            10'h0c7 	:	o_val <= 16'b0001100011100000;
            10'h0c8 	:	o_val <= 16'b0001100100000000;
            10'h0c9 	:	o_val <= 16'b0001100100100000;
            10'h0ca 	:	o_val <= 16'b0001100101000000;
            10'h0cb 	:	o_val <= 16'b0001100101100000;
            10'h0cc 	:	o_val <= 16'b0001100110000000;
            10'h0cd 	:	o_val <= 16'b0001100110100000;
            10'h0ce 	:	o_val <= 16'b0001100111000000;
            10'h0cf 	:	o_val <= 16'b0001100111100000;
            10'h0d0 	:	o_val <= 16'b0001101000000000;
            10'h0d1 	:	o_val <= 16'b0001101000100000;
            10'h0d2 	:	o_val <= 16'b0001101001000000;
            10'h0d3 	:	o_val <= 16'b0001101001100000;
            10'h0d4 	:	o_val <= 16'b0001101010000000;
            10'h0d5 	:	o_val <= 16'b0001101010100000;
            10'h0d6 	:	o_val <= 16'b0001101011000000;
            10'h0d7 	:	o_val <= 16'b0001101011100000;
            10'h0d8 	:	o_val <= 16'b0001101100000000;
            10'h0d9 	:	o_val <= 16'b0001101100100000;
            10'h0da 	:	o_val <= 16'b0001101101000000;
            10'h0db 	:	o_val <= 16'b0001101101100000;
            10'h0dc 	:	o_val <= 16'b0001101110000000;
            10'h0dd 	:	o_val <= 16'b0001101110100000;
            10'h0de 	:	o_val <= 16'b0001101111000000;
            10'h0df 	:	o_val <= 16'b0001101111100000;
            10'h0e0 	:	o_val <= 16'b0001110000000000;
            10'h0e1 	:	o_val <= 16'b0001110000100000;
            10'h0e2 	:	o_val <= 16'b0001110001000000;
            10'h0e3 	:	o_val <= 16'b0001110001100000;
            10'h0e4 	:	o_val <= 16'b0001110010000000;
            10'h0e5 	:	o_val <= 16'b0001110010100000;
            10'h0e6 	:	o_val <= 16'b0001110011000000;
            10'h0e7 	:	o_val <= 16'b0001110011100000;
            10'h0e8 	:	o_val <= 16'b0001110100000000;
            10'h0e9 	:	o_val <= 16'b0001110100100000;
            10'h0ea 	:	o_val <= 16'b0001110101000000;
            10'h0eb 	:	o_val <= 16'b0001110101100000;
            10'h0ec 	:	o_val <= 16'b0001110110000000;
            10'h0ed 	:	o_val <= 16'b0001110110100000;
            10'h0ee 	:	o_val <= 16'b0001110111000000;
            10'h0ef 	:	o_val <= 16'b0001110111100000;
            10'h0f0 	:	o_val <= 16'b0001111000000000;
            10'h0f1 	:	o_val <= 16'b0001111000100000;
            10'h0f2 	:	o_val <= 16'b0001111001000000;
            10'h0f3 	:	o_val <= 16'b0001111001100000;
            10'h0f4 	:	o_val <= 16'b0001111010000000;
            10'h0f5 	:	o_val <= 16'b0001111010100000;
            10'h0f6 	:	o_val <= 16'b0001111011000000;
            10'h0f7 	:	o_val <= 16'b0001111011100000;
            10'h0f8 	:	o_val <= 16'b0001111100000000;
            10'h0f9 	:	o_val <= 16'b0001111100100000;
            10'h0fa 	:	o_val <= 16'b0001111101000000;
            10'h0fb 	:	o_val <= 16'b0001111101100000;
            10'h0fc 	:	o_val <= 16'b0001111110000000;
            10'h0fd 	:	o_val <= 16'b0001111110100000;
            10'h0fe 	:	o_val <= 16'b0001111111000000;
            10'h0ff 	:	o_val <= 16'b0001111111100000;
            10'h100 	:	o_val <= 16'b0010000000000000;
            10'h101 	:	o_val <= 16'b0010000000100000;
            10'h102 	:	o_val <= 16'b0010000001000000;
            10'h103 	:	o_val <= 16'b0010000001100000;
            10'h104 	:	o_val <= 16'b0010000010000000;
            10'h105 	:	o_val <= 16'b0010000010100000;
            10'h106 	:	o_val <= 16'b0010000011000000;
            10'h107 	:	o_val <= 16'b0010000011100000;
            10'h108 	:	o_val <= 16'b0010000100000000;
            10'h109 	:	o_val <= 16'b0010000100100000;
            10'h10a 	:	o_val <= 16'b0010000101000000;
            10'h10b 	:	o_val <= 16'b0010000101100000;
            10'h10c 	:	o_val <= 16'b0010000110000000;
            10'h10d 	:	o_val <= 16'b0010000110100000;
            10'h10e 	:	o_val <= 16'b0010000111000000;
            10'h10f 	:	o_val <= 16'b0010000111100000;
            10'h110 	:	o_val <= 16'b0010001000000000;
            10'h111 	:	o_val <= 16'b0010001000100000;
            10'h112 	:	o_val <= 16'b0010001001000000;
            10'h113 	:	o_val <= 16'b0010001001100000;
            10'h114 	:	o_val <= 16'b0010001010000000;
            10'h115 	:	o_val <= 16'b0010001010100000;
            10'h116 	:	o_val <= 16'b0010001011000000;
            10'h117 	:	o_val <= 16'b0010001011100000;
            10'h118 	:	o_val <= 16'b0010001100000000;
            10'h119 	:	o_val <= 16'b0010001100100000;
            10'h11a 	:	o_val <= 16'b0010001101000000;
            10'h11b 	:	o_val <= 16'b0010001101100000;
            10'h11c 	:	o_val <= 16'b0010001110000000;
            10'h11d 	:	o_val <= 16'b0010001110100000;
            10'h11e 	:	o_val <= 16'b0010001111000000;
            10'h11f 	:	o_val <= 16'b0010001111100000;
            10'h120 	:	o_val <= 16'b0010010000000000;
            10'h121 	:	o_val <= 16'b0010010000100000;
            10'h122 	:	o_val <= 16'b0010010001000000;
            10'h123 	:	o_val <= 16'b0010010001100000;
            10'h124 	:	o_val <= 16'b0010010010000000;
            10'h125 	:	o_val <= 16'b0010010010100000;
            10'h126 	:	o_val <= 16'b0010010011000000;
            10'h127 	:	o_val <= 16'b0010010011100000;
            10'h128 	:	o_val <= 16'b0010010100000000;
            10'h129 	:	o_val <= 16'b0010010100100000;
            10'h12a 	:	o_val <= 16'b0010010101000000;
            10'h12b 	:	o_val <= 16'b0010010101100000;
            10'h12c 	:	o_val <= 16'b0010010110000000;
            10'h12d 	:	o_val <= 16'b0010010110100000;
            10'h12e 	:	o_val <= 16'b0010010111000000;
            10'h12f 	:	o_val <= 16'b0010010111100000;
            10'h130 	:	o_val <= 16'b0010011000000000;
            10'h131 	:	o_val <= 16'b0010011000100000;
            10'h132 	:	o_val <= 16'b0010011001000000;
            10'h133 	:	o_val <= 16'b0010011001100000;
            10'h134 	:	o_val <= 16'b0010011010000000;
            10'h135 	:	o_val <= 16'b0010011010100000;
            10'h136 	:	o_val <= 16'b0010011011000000;
            10'h137 	:	o_val <= 16'b0010011011100000;
            10'h138 	:	o_val <= 16'b0010011100000000;
            10'h139 	:	o_val <= 16'b0010011100100000;
            10'h13a 	:	o_val <= 16'b0010011101000000;
            10'h13b 	:	o_val <= 16'b0010011101100000;
            10'h13c 	:	o_val <= 16'b0010011110000000;
            10'h13d 	:	o_val <= 16'b0010011110100000;
            10'h13e 	:	o_val <= 16'b0010011111000000;
            10'h13f 	:	o_val <= 16'b0010011111100000;
            10'h140 	:	o_val <= 16'b0010100000000000;
            10'h141 	:	o_val <= 16'b0010100000100000;
            10'h142 	:	o_val <= 16'b0010100001000000;
            10'h143 	:	o_val <= 16'b0010100001100000;
            10'h144 	:	o_val <= 16'b0010100010000000;
            10'h145 	:	o_val <= 16'b0010100010100000;
            10'h146 	:	o_val <= 16'b0010100011000000;
            10'h147 	:	o_val <= 16'b0010100011100000;
            10'h148 	:	o_val <= 16'b0010100100000000;
            10'h149 	:	o_val <= 16'b0010100100100000;
            10'h14a 	:	o_val <= 16'b0010100101000000;
            10'h14b 	:	o_val <= 16'b0010100101100000;
            10'h14c 	:	o_val <= 16'b0010100110000000;
            10'h14d 	:	o_val <= 16'b0010100110100000;
            10'h14e 	:	o_val <= 16'b0010100111000000;
            10'h14f 	:	o_val <= 16'b0010100111100000;
            10'h150 	:	o_val <= 16'b0010101000000000;
            10'h151 	:	o_val <= 16'b0010101000100000;
            10'h152 	:	o_val <= 16'b0010101001000000;
            10'h153 	:	o_val <= 16'b0010101001100000;
            10'h154 	:	o_val <= 16'b0010101010000000;
            10'h155 	:	o_val <= 16'b0010101010100000;
            10'h156 	:	o_val <= 16'b0010101011000000;
            10'h157 	:	o_val <= 16'b0010101011100000;
            10'h158 	:	o_val <= 16'b0010101100000000;
            10'h159 	:	o_val <= 16'b0010101100100000;
            10'h15a 	:	o_val <= 16'b0010101101000000;
            10'h15b 	:	o_val <= 16'b0010101101100000;
            10'h15c 	:	o_val <= 16'b0010101110000000;
            10'h15d 	:	o_val <= 16'b0010101110100000;
            10'h15e 	:	o_val <= 16'b0010101111000000;
            10'h15f 	:	o_val <= 16'b0010101111100000;
            10'h160 	:	o_val <= 16'b0010110000000000;
            10'h161 	:	o_val <= 16'b0010110000100000;
            10'h162 	:	o_val <= 16'b0010110001000000;
            10'h163 	:	o_val <= 16'b0010110001100000;
            10'h164 	:	o_val <= 16'b0010110010000000;
            10'h165 	:	o_val <= 16'b0010110010100000;
            10'h166 	:	o_val <= 16'b0010110011000000;
            10'h167 	:	o_val <= 16'b0010110011100000;
            10'h168 	:	o_val <= 16'b0010110100000000;
            10'h169 	:	o_val <= 16'b0010110100100000;
            10'h16a 	:	o_val <= 16'b0010110101000000;
            10'h16b 	:	o_val <= 16'b0010110101100000;
            10'h16c 	:	o_val <= 16'b0010110110000000;
            10'h16d 	:	o_val <= 16'b0010110110100000;
            10'h16e 	:	o_val <= 16'b0010110111000000;
            10'h16f 	:	o_val <= 16'b0010110111100000;
            10'h170 	:	o_val <= 16'b0010111000000000;
            10'h171 	:	o_val <= 16'b0010111000100000;
            10'h172 	:	o_val <= 16'b0010111001000000;
            10'h173 	:	o_val <= 16'b0010111001100000;
            10'h174 	:	o_val <= 16'b0010111010000000;
            10'h175 	:	o_val <= 16'b0010111010100000;
            10'h176 	:	o_val <= 16'b0010111011000000;
            10'h177 	:	o_val <= 16'b0010111011100000;
            10'h178 	:	o_val <= 16'b0010111100000000;
            10'h179 	:	o_val <= 16'b0010111100100000;
            10'h17a 	:	o_val <= 16'b0010111101000000;
            10'h17b 	:	o_val <= 16'b0010111101100000;
            10'h17c 	:	o_val <= 16'b0010111110000000;
            10'h17d 	:	o_val <= 16'b0010111110100000;
            10'h17e 	:	o_val <= 16'b0010111111000000;
            10'h17f 	:	o_val <= 16'b0010111111100000;
            10'h180 	:	o_val <= 16'b0011000000000000;
            10'h181 	:	o_val <= 16'b0011000000100000;
            10'h182 	:	o_val <= 16'b0011000001000000;
            10'h183 	:	o_val <= 16'b0011000001100000;
            10'h184 	:	o_val <= 16'b0011000010000000;
            10'h185 	:	o_val <= 16'b0011000010100000;
            10'h186 	:	o_val <= 16'b0011000011000000;
            10'h187 	:	o_val <= 16'b0011000011100000;
            10'h188 	:	o_val <= 16'b0011000100000000;
            10'h189 	:	o_val <= 16'b0011000100100000;
            10'h18a 	:	o_val <= 16'b0011000101000000;
            10'h18b 	:	o_val <= 16'b0011000101100000;
            10'h18c 	:	o_val <= 16'b0011000110000000;
            10'h18d 	:	o_val <= 16'b0011000110100000;
            10'h18e 	:	o_val <= 16'b0011000111000000;
            10'h18f 	:	o_val <= 16'b0011000111100000;
            10'h190 	:	o_val <= 16'b0011001000000000;
            10'h191 	:	o_val <= 16'b0011001000100000;
            10'h192 	:	o_val <= 16'b0011001001000000;
            10'h193 	:	o_val <= 16'b0011001001100000;
            10'h194 	:	o_val <= 16'b0011001010000000;
            10'h195 	:	o_val <= 16'b0011001010100000;
            10'h196 	:	o_val <= 16'b0011001011000000;
            10'h197 	:	o_val <= 16'b0011001011100000;
            10'h198 	:	o_val <= 16'b0011001100000000;
            10'h199 	:	o_val <= 16'b0011001100100000;
            10'h19a 	:	o_val <= 16'b0011001101000000;
            10'h19b 	:	o_val <= 16'b0011001101100000;
            10'h19c 	:	o_val <= 16'b0011001110000000;
            10'h19d 	:	o_val <= 16'b0011001110100000;
            10'h19e 	:	o_val <= 16'b0011001111000000;
            10'h19f 	:	o_val <= 16'b0011001111100000;
            10'h1a0 	:	o_val <= 16'b0011010000000000;
            10'h1a1 	:	o_val <= 16'b0011010000100000;
            10'h1a2 	:	o_val <= 16'b0011010001000000;
            10'h1a3 	:	o_val <= 16'b0011010001100000;
            10'h1a4 	:	o_val <= 16'b0011010010000000;
            10'h1a5 	:	o_val <= 16'b0011010010100000;
            10'h1a6 	:	o_val <= 16'b0011010011000000;
            10'h1a7 	:	o_val <= 16'b0011010011100000;
            10'h1a8 	:	o_val <= 16'b0011010100000000;
            10'h1a9 	:	o_val <= 16'b0011010100100000;
            10'h1aa 	:	o_val <= 16'b0011010101000000;
            10'h1ab 	:	o_val <= 16'b0011010101100000;
            10'h1ac 	:	o_val <= 16'b0011010110000000;
            10'h1ad 	:	o_val <= 16'b0011010110100000;
            10'h1ae 	:	o_val <= 16'b0011010111000000;
            10'h1af 	:	o_val <= 16'b0011010111100000;
            10'h1b0 	:	o_val <= 16'b0011011000000000;
            10'h1b1 	:	o_val <= 16'b0011011000100000;
            10'h1b2 	:	o_val <= 16'b0011011001000000;
            10'h1b3 	:	o_val <= 16'b0011011001100000;
            10'h1b4 	:	o_val <= 16'b0011011010000000;
            10'h1b5 	:	o_val <= 16'b0011011010100000;
            10'h1b6 	:	o_val <= 16'b0011011011000000;
            10'h1b7 	:	o_val <= 16'b0011011011100000;
            10'h1b8 	:	o_val <= 16'b0011011100000000;
            10'h1b9 	:	o_val <= 16'b0011011100100000;
            10'h1ba 	:	o_val <= 16'b0011011101000000;
            10'h1bb 	:	o_val <= 16'b0011011101100000;
            10'h1bc 	:	o_val <= 16'b0011011110000000;
            10'h1bd 	:	o_val <= 16'b0011011110100000;
            10'h1be 	:	o_val <= 16'b0011011111000000;
            10'h1bf 	:	o_val <= 16'b0011011111100000;
            10'h1c0 	:	o_val <= 16'b0011100000000000;
            10'h1c1 	:	o_val <= 16'b0011100000100000;
            10'h1c2 	:	o_val <= 16'b0011100001000000;
            10'h1c3 	:	o_val <= 16'b0011100001100000;
            10'h1c4 	:	o_val <= 16'b0011100010000000;
            10'h1c5 	:	o_val <= 16'b0011100010100000;
            10'h1c6 	:	o_val <= 16'b0011100011000000;
            10'h1c7 	:	o_val <= 16'b0011100011100000;
            10'h1c8 	:	o_val <= 16'b0011100100000000;
            10'h1c9 	:	o_val <= 16'b0011100100100000;
            10'h1ca 	:	o_val <= 16'b0011100101000000;
            10'h1cb 	:	o_val <= 16'b0011100101100000;
            10'h1cc 	:	o_val <= 16'b0011100110000000;
            10'h1cd 	:	o_val <= 16'b0011100110100000;
            10'h1ce 	:	o_val <= 16'b0011100111000000;
            10'h1cf 	:	o_val <= 16'b0011100111100000;
            10'h1d0 	:	o_val <= 16'b0011101000000000;
            10'h1d1 	:	o_val <= 16'b0011101000100000;
            10'h1d2 	:	o_val <= 16'b0011101001000000;
            10'h1d3 	:	o_val <= 16'b0011101001100000;
            10'h1d4 	:	o_val <= 16'b0011101010000000;
            10'h1d5 	:	o_val <= 16'b0011101010100000;
            10'h1d6 	:	o_val <= 16'b0011101011000000;
            10'h1d7 	:	o_val <= 16'b0011101011100000;
            10'h1d8 	:	o_val <= 16'b0011101100000000;
            10'h1d9 	:	o_val <= 16'b0011101100100000;
            10'h1da 	:	o_val <= 16'b0011101101000000;
            10'h1db 	:	o_val <= 16'b0011101101100000;
            10'h1dc 	:	o_val <= 16'b0011101110000000;
            10'h1dd 	:	o_val <= 16'b0011101110100000;
            10'h1de 	:	o_val <= 16'b0011101111000000;
            10'h1df 	:	o_val <= 16'b0011101111100000;
            10'h1e0 	:	o_val <= 16'b0011110000000000;
            10'h1e1 	:	o_val <= 16'b0011110000100000;
            10'h1e2 	:	o_val <= 16'b0011110001000000;
            10'h1e3 	:	o_val <= 16'b0011110001100000;
            10'h1e4 	:	o_val <= 16'b0011110010000000;
            10'h1e5 	:	o_val <= 16'b0011110010100000;
            10'h1e6 	:	o_val <= 16'b0011110011000000;
            10'h1e7 	:	o_val <= 16'b0011110011100000;
            10'h1e8 	:	o_val <= 16'b0011110100000000;
            10'h1e9 	:	o_val <= 16'b0011110100100000;
            10'h1ea 	:	o_val <= 16'b0011110101000000;
            10'h1eb 	:	o_val <= 16'b0011110101100000;
            10'h1ec 	:	o_val <= 16'b0011110110000000;
            10'h1ed 	:	o_val <= 16'b0011110110100000;
            10'h1ee 	:	o_val <= 16'b0011110111000000;
            10'h1ef 	:	o_val <= 16'b0011110111100000;
            10'h1f0 	:	o_val <= 16'b0011111000000000;
            10'h1f1 	:	o_val <= 16'b0011111000100000;
            10'h1f2 	:	o_val <= 16'b0011111001000000;
            10'h1f3 	:	o_val <= 16'b0011111001100000;
            10'h1f4 	:	o_val <= 16'b0011111010000000;
            10'h1f5 	:	o_val <= 16'b0011111010100000;
            10'h1f6 	:	o_val <= 16'b0011111011000000;
            10'h1f7 	:	o_val <= 16'b0011111011100000;
            10'h1f8 	:	o_val <= 16'b0011111100000000;
            10'h1f9 	:	o_val <= 16'b0011111100100000;
            10'h1fa 	:	o_val <= 16'b0011111101000000;
            10'h1fb 	:	o_val <= 16'b0011111101100000;
            10'h1fc 	:	o_val <= 16'b0011111110000000;
            10'h1fd 	:	o_val <= 16'b0011111110100000;
            10'h1fe 	:	o_val <= 16'b0011111111000000;
            10'h1ff 	:	o_val <= 16'b0011111111100000;
            10'h200 	:	o_val <= 16'b0100000000000000;
            10'h201 	:	o_val <= 16'b0100000000100000;
            10'h202 	:	o_val <= 16'b0100000001000000;
            10'h203 	:	o_val <= 16'b0100000001100000;
            10'h204 	:	o_val <= 16'b0100000010000000;
            10'h205 	:	o_val <= 16'b0100000010100000;
            10'h206 	:	o_val <= 16'b0100000011000000;
            10'h207 	:	o_val <= 16'b0100000011100000;
            10'h208 	:	o_val <= 16'b0100000100000000;
            10'h209 	:	o_val <= 16'b0100000100100000;
            10'h20a 	:	o_val <= 16'b0100000101000000;
            10'h20b 	:	o_val <= 16'b0100000101100000;
            10'h20c 	:	o_val <= 16'b0100000110000000;
            10'h20d 	:	o_val <= 16'b0100000110100000;
            10'h20e 	:	o_val <= 16'b0100000111000000;
            10'h20f 	:	o_val <= 16'b0100000111100000;
            10'h210 	:	o_val <= 16'b0100001000000000;
            10'h211 	:	o_val <= 16'b0100001000100000;
            10'h212 	:	o_val <= 16'b0100001001000000;
            10'h213 	:	o_val <= 16'b0100001001100000;
            10'h214 	:	o_val <= 16'b0100001010000000;
            10'h215 	:	o_val <= 16'b0100001010100000;
            10'h216 	:	o_val <= 16'b0100001011000000;
            10'h217 	:	o_val <= 16'b0100001011100000;
            10'h218 	:	o_val <= 16'b0100001100000000;
            10'h219 	:	o_val <= 16'b0100001100100000;
            10'h21a 	:	o_val <= 16'b0100001101000000;
            10'h21b 	:	o_val <= 16'b0100001101100000;
            10'h21c 	:	o_val <= 16'b0100001110000000;
            10'h21d 	:	o_val <= 16'b0100001110100000;
            10'h21e 	:	o_val <= 16'b0100001111000000;
            10'h21f 	:	o_val <= 16'b0100001111100000;
            10'h220 	:	o_val <= 16'b0100010000000000;
            10'h221 	:	o_val <= 16'b0100010000100000;
            10'h222 	:	o_val <= 16'b0100010001000000;
            10'h223 	:	o_val <= 16'b0100010001100000;
            10'h224 	:	o_val <= 16'b0100010010000000;
            10'h225 	:	o_val <= 16'b0100010010100000;
            10'h226 	:	o_val <= 16'b0100010011000000;
            10'h227 	:	o_val <= 16'b0100010011100000;
            10'h228 	:	o_val <= 16'b0100010100000000;
            10'h229 	:	o_val <= 16'b0100010100100000;
            10'h22a 	:	o_val <= 16'b0100010101000000;
            10'h22b 	:	o_val <= 16'b0100010101100000;
            10'h22c 	:	o_val <= 16'b0100010110000000;
            10'h22d 	:	o_val <= 16'b0100010110100000;
            10'h22e 	:	o_val <= 16'b0100010111000000;
            10'h22f 	:	o_val <= 16'b0100010111100000;
            10'h230 	:	o_val <= 16'b0100011000000000;
            10'h231 	:	o_val <= 16'b0100011000100000;
            10'h232 	:	o_val <= 16'b0100011001000000;
            10'h233 	:	o_val <= 16'b0100011001100000;
            10'h234 	:	o_val <= 16'b0100011010000000;
            10'h235 	:	o_val <= 16'b0100011010100000;
            10'h236 	:	o_val <= 16'b0100011011000000;
            10'h237 	:	o_val <= 16'b0100011011100000;
            10'h238 	:	o_val <= 16'b0100011100000000;
            10'h239 	:	o_val <= 16'b0100011100100000;
            10'h23a 	:	o_val <= 16'b0100011101000000;
            10'h23b 	:	o_val <= 16'b0100011101100000;
            10'h23c 	:	o_val <= 16'b0100011110000000;
            10'h23d 	:	o_val <= 16'b0100011110100000;
            10'h23e 	:	o_val <= 16'b0100011111000000;
            10'h23f 	:	o_val <= 16'b0100011111100000;
            10'h240 	:	o_val <= 16'b0100100000000000;
            10'h241 	:	o_val <= 16'b0100100000100000;
            10'h242 	:	o_val <= 16'b0100100001000000;
            10'h243 	:	o_val <= 16'b0100100001100000;
            10'h244 	:	o_val <= 16'b0100100010000000;
            10'h245 	:	o_val <= 16'b0100100010100000;
            10'h246 	:	o_val <= 16'b0100100011000000;
            10'h247 	:	o_val <= 16'b0100100011100000;
            10'h248 	:	o_val <= 16'b0100100100000000;
            10'h249 	:	o_val <= 16'b0100100100100000;
            10'h24a 	:	o_val <= 16'b0100100101000000;
            10'h24b 	:	o_val <= 16'b0100100101100000;
            10'h24c 	:	o_val <= 16'b0100100110000000;
            10'h24d 	:	o_val <= 16'b0100100110100000;
            10'h24e 	:	o_val <= 16'b0100100111000000;
            10'h24f 	:	o_val <= 16'b0100100111100000;
            10'h250 	:	o_val <= 16'b0100101000000000;
            10'h251 	:	o_val <= 16'b0100101000100000;
            10'h252 	:	o_val <= 16'b0100101001000000;
            10'h253 	:	o_val <= 16'b0100101001100000;
            10'h254 	:	o_val <= 16'b0100101010000000;
            10'h255 	:	o_val <= 16'b0100101010100000;
            10'h256 	:	o_val <= 16'b0100101011000000;
            10'h257 	:	o_val <= 16'b0100101011100000;
            10'h258 	:	o_val <= 16'b0100101100000000;
            10'h259 	:	o_val <= 16'b0100101100100000;
            10'h25a 	:	o_val <= 16'b0100101101000000;
            10'h25b 	:	o_val <= 16'b0100101101100000;
            10'h25c 	:	o_val <= 16'b0100101110000000;
            10'h25d 	:	o_val <= 16'b0100101110100000;
            10'h25e 	:	o_val <= 16'b0100101111000000;
            10'h25f 	:	o_val <= 16'b0100101111100000;
            10'h260 	:	o_val <= 16'b0100110000000000;
            10'h261 	:	o_val <= 16'b0100110000100000;
            10'h262 	:	o_val <= 16'b0100110001000000;
            10'h263 	:	o_val <= 16'b0100110001100000;
            10'h264 	:	o_val <= 16'b0100110010000000;
            10'h265 	:	o_val <= 16'b0100110010100000;
            10'h266 	:	o_val <= 16'b0100110011000000;
            10'h267 	:	o_val <= 16'b0100110011100000;
            10'h268 	:	o_val <= 16'b0100110100000000;
            10'h269 	:	o_val <= 16'b0100110100100000;
            10'h26a 	:	o_val <= 16'b0100110101000000;
            10'h26b 	:	o_val <= 16'b0100110101100000;
            10'h26c 	:	o_val <= 16'b0100110110000000;
            10'h26d 	:	o_val <= 16'b0100110110100000;
            10'h26e 	:	o_val <= 16'b0100110111000000;
            10'h26f 	:	o_val <= 16'b0100110111100000;
            10'h270 	:	o_val <= 16'b0100111000000000;
            10'h271 	:	o_val <= 16'b0100111000100000;
            10'h272 	:	o_val <= 16'b0100111001000000;
            10'h273 	:	o_val <= 16'b0100111001100000;
            10'h274 	:	o_val <= 16'b0100111010000000;
            10'h275 	:	o_val <= 16'b0100111010100000;
            10'h276 	:	o_val <= 16'b0100111011000000;
            10'h277 	:	o_val <= 16'b0100111011100000;
            10'h278 	:	o_val <= 16'b0100111100000000;
            10'h279 	:	o_val <= 16'b0100111100100000;
            10'h27a 	:	o_val <= 16'b0100111101000000;
            10'h27b 	:	o_val <= 16'b0100111101100000;
            10'h27c 	:	o_val <= 16'b0100111110000000;
            10'h27d 	:	o_val <= 16'b0100111110100000;
            10'h27e 	:	o_val <= 16'b0100111111000000;
            10'h27f 	:	o_val <= 16'b0100111111100000;
            10'h280 	:	o_val <= 16'b0101000000000000;
            10'h281 	:	o_val <= 16'b0101000000100000;
            10'h282 	:	o_val <= 16'b0101000001000000;
            10'h283 	:	o_val <= 16'b0101000001100000;
            10'h284 	:	o_val <= 16'b0101000010000000;
            10'h285 	:	o_val <= 16'b0101000010100000;
            10'h286 	:	o_val <= 16'b0101000011000000;
            10'h287 	:	o_val <= 16'b0101000011100000;
            10'h288 	:	o_val <= 16'b0101000100000000;
            10'h289 	:	o_val <= 16'b0101000100100000;
            10'h28a 	:	o_val <= 16'b0101000101000000;
            10'h28b 	:	o_val <= 16'b0101000101100000;
            10'h28c 	:	o_val <= 16'b0101000110000000;
            10'h28d 	:	o_val <= 16'b0101000110100000;
            10'h28e 	:	o_val <= 16'b0101000111000000;
            10'h28f 	:	o_val <= 16'b0101000111100000;
            10'h290 	:	o_val <= 16'b0101001000000000;
            10'h291 	:	o_val <= 16'b0101001000100000;
            10'h292 	:	o_val <= 16'b0101001001000000;
            10'h293 	:	o_val <= 16'b0101001001100000;
            10'h294 	:	o_val <= 16'b0101001010000000;
            10'h295 	:	o_val <= 16'b0101001010100000;
            10'h296 	:	o_val <= 16'b0101001011000000;
            10'h297 	:	o_val <= 16'b0101001011100000;
            10'h298 	:	o_val <= 16'b0101001100000000;
            10'h299 	:	o_val <= 16'b0101001100100000;
            10'h29a 	:	o_val <= 16'b0101001101000000;
            10'h29b 	:	o_val <= 16'b0101001101100000;
            10'h29c 	:	o_val <= 16'b0101001110000000;
            10'h29d 	:	o_val <= 16'b0101001110100000;
            10'h29e 	:	o_val <= 16'b0101001111000000;
            10'h29f 	:	o_val <= 16'b0101001111100000;
            10'h2a0 	:	o_val <= 16'b0101010000000000;
            10'h2a1 	:	o_val <= 16'b0101010000100000;
            10'h2a2 	:	o_val <= 16'b0101010001000000;
            10'h2a3 	:	o_val <= 16'b0101010001100000;
            10'h2a4 	:	o_val <= 16'b0101010010000000;
            10'h2a5 	:	o_val <= 16'b0101010010100000;
            10'h2a6 	:	o_val <= 16'b0101010011000000;
            10'h2a7 	:	o_val <= 16'b0101010011100000;
            10'h2a8 	:	o_val <= 16'b0101010100000000;
            10'h2a9 	:	o_val <= 16'b0101010100100000;
            10'h2aa 	:	o_val <= 16'b0101010101000000;
            10'h2ab 	:	o_val <= 16'b0101010101100000;
            10'h2ac 	:	o_val <= 16'b0101010110000000;
            10'h2ad 	:	o_val <= 16'b0101010110100000;
            10'h2ae 	:	o_val <= 16'b0101010111000000;
            10'h2af 	:	o_val <= 16'b0101010111100000;
            10'h2b0 	:	o_val <= 16'b0101011000000000;
            10'h2b1 	:	o_val <= 16'b0101011000100000;
            10'h2b2 	:	o_val <= 16'b0101011001000000;
            10'h2b3 	:	o_val <= 16'b0101011001100000;
            10'h2b4 	:	o_val <= 16'b0101011010000000;
            10'h2b5 	:	o_val <= 16'b0101011010100000;
            10'h2b6 	:	o_val <= 16'b0101011011000000;
            10'h2b7 	:	o_val <= 16'b0101011011100000;
            10'h2b8 	:	o_val <= 16'b0101011100000000;
            10'h2b9 	:	o_val <= 16'b0101011100100000;
            10'h2ba 	:	o_val <= 16'b0101011101000000;
            10'h2bb 	:	o_val <= 16'b0101011101100000;
            10'h2bc 	:	o_val <= 16'b0101011110000000;
            10'h2bd 	:	o_val <= 16'b0101011110100000;
            10'h2be 	:	o_val <= 16'b0101011111000000;
            10'h2bf 	:	o_val <= 16'b0101011111100000;
            10'h2c0 	:	o_val <= 16'b0101100000000000;
            10'h2c1 	:	o_val <= 16'b0101100000100000;
            10'h2c2 	:	o_val <= 16'b0101100001000000;
            10'h2c3 	:	o_val <= 16'b0101100001100000;
            10'h2c4 	:	o_val <= 16'b0101100010000000;
            10'h2c5 	:	o_val <= 16'b0101100010100000;
            10'h2c6 	:	o_val <= 16'b0101100011000000;
            10'h2c7 	:	o_val <= 16'b0101100011100000;
            10'h2c8 	:	o_val <= 16'b0101100100000000;
            10'h2c9 	:	o_val <= 16'b0101100100100000;
            10'h2ca 	:	o_val <= 16'b0101100101000000;
            10'h2cb 	:	o_val <= 16'b0101100101100000;
            10'h2cc 	:	o_val <= 16'b0101100110000000;
            10'h2cd 	:	o_val <= 16'b0101100110100000;
            10'h2ce 	:	o_val <= 16'b0101100111000000;
            10'h2cf 	:	o_val <= 16'b0101100111100000;
            10'h2d0 	:	o_val <= 16'b0101101000000000;
            10'h2d1 	:	o_val <= 16'b0101101000100000;
            10'h2d2 	:	o_val <= 16'b0101101001000000;
            10'h2d3 	:	o_val <= 16'b0101101001100000;
            10'h2d4 	:	o_val <= 16'b0101101010000000;
            10'h2d5 	:	o_val <= 16'b0101101010100000;
            10'h2d6 	:	o_val <= 16'b0101101011000000;
            10'h2d7 	:	o_val <= 16'b0101101011100000;
            10'h2d8 	:	o_val <= 16'b0101101100000000;
            10'h2d9 	:	o_val <= 16'b0101101100100000;
            10'h2da 	:	o_val <= 16'b0101101101000000;
            10'h2db 	:	o_val <= 16'b0101101101100000;
            10'h2dc 	:	o_val <= 16'b0101101110000000;
            10'h2dd 	:	o_val <= 16'b0101101110100000;
            10'h2de 	:	o_val <= 16'b0101101111000000;
            10'h2df 	:	o_val <= 16'b0101101111100000;
            10'h2e0 	:	o_val <= 16'b0101110000000000;
            10'h2e1 	:	o_val <= 16'b0101110000100000;
            10'h2e2 	:	o_val <= 16'b0101110001000000;
            10'h2e3 	:	o_val <= 16'b0101110001100000;
            10'h2e4 	:	o_val <= 16'b0101110010000000;
            10'h2e5 	:	o_val <= 16'b0101110010100000;
            10'h2e6 	:	o_val <= 16'b0101110011000000;
            10'h2e7 	:	o_val <= 16'b0101110011100000;
            10'h2e8 	:	o_val <= 16'b0101110100000000;
            10'h2e9 	:	o_val <= 16'b0101110100100000;
            10'h2ea 	:	o_val <= 16'b0101110101000000;
            10'h2eb 	:	o_val <= 16'b0101110101100000;
            10'h2ec 	:	o_val <= 16'b0101110110000000;
            10'h2ed 	:	o_val <= 16'b0101110110100000;
            10'h2ee 	:	o_val <= 16'b0101110111000000;
            10'h2ef 	:	o_val <= 16'b0101110111100000;
            10'h2f0 	:	o_val <= 16'b0101111000000000;
            10'h2f1 	:	o_val <= 16'b0101111000100000;
            10'h2f2 	:	o_val <= 16'b0101111001000000;
            10'h2f3 	:	o_val <= 16'b0101111001100000;
            10'h2f4 	:	o_val <= 16'b0101111010000000;
            10'h2f5 	:	o_val <= 16'b0101111010100000;
            10'h2f6 	:	o_val <= 16'b0101111011000000;
            10'h2f7 	:	o_val <= 16'b0101111011100000;
            10'h2f8 	:	o_val <= 16'b0101111100000000;
            10'h2f9 	:	o_val <= 16'b0101111100100000;
            10'h2fa 	:	o_val <= 16'b0101111101000000;
            10'h2fb 	:	o_val <= 16'b0101111101100000;
            10'h2fc 	:	o_val <= 16'b0101111110000000;
            10'h2fd 	:	o_val <= 16'b0101111110100000;
            10'h2fe 	:	o_val <= 16'b0101111111000000;
            10'h2ff 	:	o_val <= 16'b0101111111100000;
            10'h300 	:	o_val <= 16'b0110000000000000;
            10'h301 	:	o_val <= 16'b0110000000100000;
            10'h302 	:	o_val <= 16'b0110000001000000;
            10'h303 	:	o_val <= 16'b0110000001100000;
            10'h304 	:	o_val <= 16'b0110000010000000;
            10'h305 	:	o_val <= 16'b0110000010100000;
            10'h306 	:	o_val <= 16'b0110000011000000;
            10'h307 	:	o_val <= 16'b0110000011100000;
            10'h308 	:	o_val <= 16'b0110000100000000;
            10'h309 	:	o_val <= 16'b0110000100100000;
            10'h30a 	:	o_val <= 16'b0110000101000000;
            10'h30b 	:	o_val <= 16'b0110000101100000;
            10'h30c 	:	o_val <= 16'b0110000110000000;
            10'h30d 	:	o_val <= 16'b0110000110100000;
            10'h30e 	:	o_val <= 16'b0110000111000000;
            10'h30f 	:	o_val <= 16'b0110000111100000;
            10'h310 	:	o_val <= 16'b0110001000000000;
            10'h311 	:	o_val <= 16'b0110001000100000;
            10'h312 	:	o_val <= 16'b0110001001000000;
            10'h313 	:	o_val <= 16'b0110001001100000;
            10'h314 	:	o_val <= 16'b0110001010000000;
            10'h315 	:	o_val <= 16'b0110001010100000;
            10'h316 	:	o_val <= 16'b0110001011000000;
            10'h317 	:	o_val <= 16'b0110001011100000;
            10'h318 	:	o_val <= 16'b0110001100000000;
            10'h319 	:	o_val <= 16'b0110001100100000;
            10'h31a 	:	o_val <= 16'b0110001101000000;
            10'h31b 	:	o_val <= 16'b0110001101100000;
            10'h31c 	:	o_val <= 16'b0110001110000000;
            10'h31d 	:	o_val <= 16'b0110001110100000;
            10'h31e 	:	o_val <= 16'b0110001111000000;
            10'h31f 	:	o_val <= 16'b0110001111100000;
            10'h320 	:	o_val <= 16'b0110010000000000;
            10'h321 	:	o_val <= 16'b0110010000100000;
            10'h322 	:	o_val <= 16'b0110010001000000;
            10'h323 	:	o_val <= 16'b0110010001100000;
            10'h324 	:	o_val <= 16'b0110010010000000;
            10'h325 	:	o_val <= 16'b0110010010100000;
            10'h326 	:	o_val <= 16'b0110010011000000;
            10'h327 	:	o_val <= 16'b0110010011100000;
            10'h328 	:	o_val <= 16'b0110010100000000;
            10'h329 	:	o_val <= 16'b0110010100100000;
            10'h32a 	:	o_val <= 16'b0110010101000000;
            10'h32b 	:	o_val <= 16'b0110010101100000;
            10'h32c 	:	o_val <= 16'b0110010110000000;
            10'h32d 	:	o_val <= 16'b0110010110100000;
            10'h32e 	:	o_val <= 16'b0110010111000000;
            10'h32f 	:	o_val <= 16'b0110010111100000;
            10'h330 	:	o_val <= 16'b0110011000000000;
            10'h331 	:	o_val <= 16'b0110011000100000;
            10'h332 	:	o_val <= 16'b0110011001000000;
            10'h333 	:	o_val <= 16'b0110011001100000;
            10'h334 	:	o_val <= 16'b0110011010000000;
            10'h335 	:	o_val <= 16'b0110011010100000;
            10'h336 	:	o_val <= 16'b0110011011000000;
            10'h337 	:	o_val <= 16'b0110011011100000;
            10'h338 	:	o_val <= 16'b0110011100000000;
            10'h339 	:	o_val <= 16'b0110011100100000;
            10'h33a 	:	o_val <= 16'b0110011101000000;
            10'h33b 	:	o_val <= 16'b0110011101100000;
            10'h33c 	:	o_val <= 16'b0110011110000000;
            10'h33d 	:	o_val <= 16'b0110011110100000;
            10'h33e 	:	o_val <= 16'b0110011111000000;
            10'h33f 	:	o_val <= 16'b0110011111100000;
            10'h340 	:	o_val <= 16'b0110100000000000;
            10'h341 	:	o_val <= 16'b0110100000100000;
            10'h342 	:	o_val <= 16'b0110100001000000;
            10'h343 	:	o_val <= 16'b0110100001100000;
            10'h344 	:	o_val <= 16'b0110100010000000;
            10'h345 	:	o_val <= 16'b0110100010100000;
            10'h346 	:	o_val <= 16'b0110100011000000;
            10'h347 	:	o_val <= 16'b0110100011100000;
            10'h348 	:	o_val <= 16'b0110100100000000;
            10'h349 	:	o_val <= 16'b0110100100100000;
            10'h34a 	:	o_val <= 16'b0110100101000000;
            10'h34b 	:	o_val <= 16'b0110100101100000;
            10'h34c 	:	o_val <= 16'b0110100110000000;
            10'h34d 	:	o_val <= 16'b0110100110100000;
            10'h34e 	:	o_val <= 16'b0110100111000000;
            10'h34f 	:	o_val <= 16'b0110100111100000;
            10'h350 	:	o_val <= 16'b0110101000000000;
            10'h351 	:	o_val <= 16'b0110101000100000;
            10'h352 	:	o_val <= 16'b0110101001000000;
            10'h353 	:	o_val <= 16'b0110101001100000;
            10'h354 	:	o_val <= 16'b0110101010000000;
            10'h355 	:	o_val <= 16'b0110101010100000;
            10'h356 	:	o_val <= 16'b0110101011000000;
            10'h357 	:	o_val <= 16'b0110101011100000;
            10'h358 	:	o_val <= 16'b0110101100000000;
            10'h359 	:	o_val <= 16'b0110101100100000;
            10'h35a 	:	o_val <= 16'b0110101101000000;
            10'h35b 	:	o_val <= 16'b0110101101100000;
            10'h35c 	:	o_val <= 16'b0110101110000000;
            10'h35d 	:	o_val <= 16'b0110101110100000;
            10'h35e 	:	o_val <= 16'b0110101111000000;
            10'h35f 	:	o_val <= 16'b0110101111100000;
            10'h360 	:	o_val <= 16'b0110110000000000;
            10'h361 	:	o_val <= 16'b0110110000100000;
            10'h362 	:	o_val <= 16'b0110110001000000;
            10'h363 	:	o_val <= 16'b0110110001100000;
            10'h364 	:	o_val <= 16'b0110110010000000;
            10'h365 	:	o_val <= 16'b0110110010100000;
            10'h366 	:	o_val <= 16'b0110110011000000;
            10'h367 	:	o_val <= 16'b0110110011100000;
            10'h368 	:	o_val <= 16'b0110110100000000;
            10'h369 	:	o_val <= 16'b0110110100100000;
            10'h36a 	:	o_val <= 16'b0110110101000000;
            10'h36b 	:	o_val <= 16'b0110110101100000;
            10'h36c 	:	o_val <= 16'b0110110110000000;
            10'h36d 	:	o_val <= 16'b0110110110100000;
            10'h36e 	:	o_val <= 16'b0110110111000000;
            10'h36f 	:	o_val <= 16'b0110110111100000;
            10'h370 	:	o_val <= 16'b0110111000000000;
            10'h371 	:	o_val <= 16'b0110111000100000;
            10'h372 	:	o_val <= 16'b0110111001000000;
            10'h373 	:	o_val <= 16'b0110111001100000;
            10'h374 	:	o_val <= 16'b0110111010000000;
            10'h375 	:	o_val <= 16'b0110111010100000;
            10'h376 	:	o_val <= 16'b0110111011000000;
            10'h377 	:	o_val <= 16'b0110111011100000;
            10'h378 	:	o_val <= 16'b0110111100000000;
            10'h379 	:	o_val <= 16'b0110111100100000;
            10'h37a 	:	o_val <= 16'b0110111101000000;
            10'h37b 	:	o_val <= 16'b0110111101100000;
            10'h37c 	:	o_val <= 16'b0110111110000000;
            10'h37d 	:	o_val <= 16'b0110111110100000;
            10'h37e 	:	o_val <= 16'b0110111111000000;
            10'h37f 	:	o_val <= 16'b0110111111100000;
            10'h380 	:	o_val <= 16'b0111000000000000;
            10'h381 	:	o_val <= 16'b0111000000100000;
            10'h382 	:	o_val <= 16'b0111000001000000;
            10'h383 	:	o_val <= 16'b0111000001100000;
            10'h384 	:	o_val <= 16'b0111000010000000;
            10'h385 	:	o_val <= 16'b0111000010100000;
            10'h386 	:	o_val <= 16'b0111000011000000;
            10'h387 	:	o_val <= 16'b0111000011100000;
            10'h388 	:	o_val <= 16'b0111000100000000;
            10'h389 	:	o_val <= 16'b0111000100100000;
            10'h38a 	:	o_val <= 16'b0111000101000000;
            10'h38b 	:	o_val <= 16'b0111000101100000;
            10'h38c 	:	o_val <= 16'b0111000110000000;
            10'h38d 	:	o_val <= 16'b0111000110100000;
            10'h38e 	:	o_val <= 16'b0111000111000000;
            10'h38f 	:	o_val <= 16'b0111000111100000;
            10'h390 	:	o_val <= 16'b0111001000000000;
            10'h391 	:	o_val <= 16'b0111001000100000;
            10'h392 	:	o_val <= 16'b0111001001000000;
            10'h393 	:	o_val <= 16'b0111001001100000;
            10'h394 	:	o_val <= 16'b0111001010000000;
            10'h395 	:	o_val <= 16'b0111001010100000;
            10'h396 	:	o_val <= 16'b0111001011000000;
            10'h397 	:	o_val <= 16'b0111001011100000;
            10'h398 	:	o_val <= 16'b0111001100000000;
            10'h399 	:	o_val <= 16'b0111001100100000;
            10'h39a 	:	o_val <= 16'b0111001101000000;
            10'h39b 	:	o_val <= 16'b0111001101100000;
            10'h39c 	:	o_val <= 16'b0111001110000000;
            10'h39d 	:	o_val <= 16'b0111001110100000;
            10'h39e 	:	o_val <= 16'b0111001111000000;
            10'h39f 	:	o_val <= 16'b0111001111100000;
            10'h3a0 	:	o_val <= 16'b0111010000000000;
            10'h3a1 	:	o_val <= 16'b0111010000100000;
            10'h3a2 	:	o_val <= 16'b0111010001000000;
            10'h3a3 	:	o_val <= 16'b0111010001100000;
            10'h3a4 	:	o_val <= 16'b0111010010000000;
            10'h3a5 	:	o_val <= 16'b0111010010100000;
            10'h3a6 	:	o_val <= 16'b0111010011000000;
            10'h3a7 	:	o_val <= 16'b0111010011100000;
            10'h3a8 	:	o_val <= 16'b0111010100000000;
            10'h3a9 	:	o_val <= 16'b0111010100100000;
            10'h3aa 	:	o_val <= 16'b0111010101000000;
            10'h3ab 	:	o_val <= 16'b0111010101100000;
            10'h3ac 	:	o_val <= 16'b0111010110000000;
            10'h3ad 	:	o_val <= 16'b0111010110100000;
            10'h3ae 	:	o_val <= 16'b0111010111000000;
            10'h3af 	:	o_val <= 16'b0111010111100000;
            10'h3b0 	:	o_val <= 16'b0111011000000000;
            10'h3b1 	:	o_val <= 16'b0111011000100000;
            10'h3b2 	:	o_val <= 16'b0111011001000000;
            10'h3b3 	:	o_val <= 16'b0111011001100000;
            10'h3b4 	:	o_val <= 16'b0111011010000000;
            10'h3b5 	:	o_val <= 16'b0111011010100000;
            10'h3b6 	:	o_val <= 16'b0111011011000000;
            10'h3b7 	:	o_val <= 16'b0111011011100000;
            10'h3b8 	:	o_val <= 16'b0111011100000000;
            10'h3b9 	:	o_val <= 16'b0111011100100000;
            10'h3ba 	:	o_val <= 16'b0111011101000000;
            10'h3bb 	:	o_val <= 16'b0111011101100000;
            10'h3bc 	:	o_val <= 16'b0111011110000000;
            10'h3bd 	:	o_val <= 16'b0111011110100000;
            10'h3be 	:	o_val <= 16'b0111011111000000;
            10'h3bf 	:	o_val <= 16'b0111011111100000;
            10'h3c0 	:	o_val <= 16'b0111100000000000;
            10'h3c1 	:	o_val <= 16'b0111100000100000;
            10'h3c2 	:	o_val <= 16'b0111100001000000;
            10'h3c3 	:	o_val <= 16'b0111100001100000;
            10'h3c4 	:	o_val <= 16'b0111100010000000;
            10'h3c5 	:	o_val <= 16'b0111100010100000;
            10'h3c6 	:	o_val <= 16'b0111100011000000;
            10'h3c7 	:	o_val <= 16'b0111100011100000;
            10'h3c8 	:	o_val <= 16'b0111100100000000;
            10'h3c9 	:	o_val <= 16'b0111100100100000;
            10'h3ca 	:	o_val <= 16'b0111100101000000;
            10'h3cb 	:	o_val <= 16'b0111100101100000;
            10'h3cc 	:	o_val <= 16'b0111100110000000;
            10'h3cd 	:	o_val <= 16'b0111100110100000;
            10'h3ce 	:	o_val <= 16'b0111100111000000;
            10'h3cf 	:	o_val <= 16'b0111100111100000;
            10'h3d0 	:	o_val <= 16'b0111101000000000;
            10'h3d1 	:	o_val <= 16'b0111101000100000;
            10'h3d2 	:	o_val <= 16'b0111101001000000;
            10'h3d3 	:	o_val <= 16'b0111101001100000;
            10'h3d4 	:	o_val <= 16'b0111101010000000;
            10'h3d5 	:	o_val <= 16'b0111101010100000;
            10'h3d6 	:	o_val <= 16'b0111101011000000;
            10'h3d7 	:	o_val <= 16'b0111101011100000;
            10'h3d8 	:	o_val <= 16'b0111101100000000;
            10'h3d9 	:	o_val <= 16'b0111101100100000;
            10'h3da 	:	o_val <= 16'b0111101101000000;
            10'h3db 	:	o_val <= 16'b0111101101100000;
            10'h3dc 	:	o_val <= 16'b0111101110000000;
            10'h3dd 	:	o_val <= 16'b0111101110100000;
            10'h3de 	:	o_val <= 16'b0111101111000000;
            10'h3df 	:	o_val <= 16'b0111101111100000;
            10'h3e0 	:	o_val <= 16'b0111110000000000;
            10'h3e1 	:	o_val <= 16'b0111110000100000;
            10'h3e2 	:	o_val <= 16'b0111110001000000;
            10'h3e3 	:	o_val <= 16'b0111110001100000;
            10'h3e4 	:	o_val <= 16'b0111110010000000;
            10'h3e5 	:	o_val <= 16'b0111110010100000;
            10'h3e6 	:	o_val <= 16'b0111110011000000;
            10'h3e7 	:	o_val <= 16'b0111110011100000;
            10'h3e8 	:	o_val <= 16'b0111110100000000;
            10'h3e9 	:	o_val <= 16'b0111110100100000;
            10'h3ea 	:	o_val <= 16'b0111110101000000;
            10'h3eb 	:	o_val <= 16'b0111110101100000;
            10'h3ec 	:	o_val <= 16'b0111110110000000;
            10'h3ed 	:	o_val <= 16'b0111110110100000;
            10'h3ee 	:	o_val <= 16'b0111110111000000;
            10'h3ef 	:	o_val <= 16'b0111110111100000;
            10'h3f0 	:	o_val <= 16'b0111111000000000;
            10'h3f1 	:	o_val <= 16'b0111111000100000;
            10'h3f2 	:	o_val <= 16'b0111111001000000;
            10'h3f3 	:	o_val <= 16'b0111111001100000;
            10'h3f4 	:	o_val <= 16'b0111111010000000;
            10'h3f5 	:	o_val <= 16'b0111111010100000;
            10'h3f6 	:	o_val <= 16'b0111111011000000;
            10'h3f7 	:	o_val <= 16'b0111111011100000;
            10'h3f8 	:	o_val <= 16'b0111111100000000;
            10'h3f9 	:	o_val <= 16'b0111111100100000;
            10'h3fa 	:	o_val <= 16'b0111111101000000;
            10'h3fb 	:	o_val <= 16'b0111111101100000;
            10'h3fc 	:	o_val <= 16'b0111111110000000;
            10'h3fd 	:	o_val <= 16'b0111111110100000;
            10'h3fe 	:	o_val <= 16'b0111111111000000;
            10'h3ff 	:	o_val <= 16'b0111111111100000;
				default		:	o_val <= 16'b0;
			endcase
		end
endmodule
              
