// modules for LUT's for multiple sinewaves for SIMPLE synthesis


//TODO: clock enable has to be given because it cannot be always enabled
// for now just A4 (440kHz) generating module (for phase calculation) 
module dummyA4(clk, phase_out); // maybe different style of coding, everything in module declaration?
	input clk;
	output reg [31:0] phase_out = 32'b0; // does it need to be initialized?
	// Phase increment can be precalculated = 188978561.024 (ignoring the truncated part) -> 2^32 * fd /fs
	
	always @(posedge clk) begin
		phase_out <= phase_out + 32'h0b43_9581;
	end
	
endmodule

// for now let's assume 8192 samples = 2^13, generate four quarters of one cycle for now (simplify later, but requires more logic)
module sineLUT(phase, val_out);
	input [15:0] phase;
	output reg [15:0] val_out;
	
	always @(phase) begin
		case (phase)         
			16'h0000, 16'h0001, 16'h0002, 16'h0003, 16'h0004, 16'h0005, 16'h0006, 16'h0007 	:	val_out <= 16'h8000;
         16'h0008, 16'h0009, 16'h000a, 16'h000b, 16'h000c, 16'h000d, 16'h000e, 16'h000f 	:	val_out <= 16'h8019;
         16'h0010, 16'h0011, 16'h0012, 16'h0013, 16'h0014, 16'h0015, 16'h0016, 16'h0017 	:	val_out <= 16'h8032;
         16'h0018, 16'h0019, 16'h001a, 16'h001b, 16'h001c, 16'h001d, 16'h001e, 16'h001f 	:	val_out <= 16'h804b;
         16'h0020, 16'h0021, 16'h0022, 16'h0023, 16'h0024, 16'h0025, 16'h0026, 16'h0027 	:	val_out <= 16'h8064;
         16'h0028, 16'h0029, 16'h002a, 16'h002b, 16'h002c, 16'h002d, 16'h002e, 16'h002f 	:	val_out <= 16'h807d;
         16'h0030, 16'h0031, 16'h0032, 16'h0033, 16'h0034, 16'h0035, 16'h0036, 16'h0037 	:	val_out <= 16'h8096;
         16'h0038, 16'h0039, 16'h003a, 16'h003b, 16'h003c, 16'h003d, 16'h003e, 16'h003f 	:	val_out <= 16'h80af;
         16'h0040, 16'h0041, 16'h0042, 16'h0043, 16'h0044, 16'h0045, 16'h0046, 16'h0047 	:	val_out <= 16'h80c9;
         16'h0048, 16'h0049, 16'h004a, 16'h004b, 16'h004c, 16'h004d, 16'h004e, 16'h004f 	:	val_out <= 16'h80e2;
         16'h0050, 16'h0051, 16'h0052, 16'h0053, 16'h0054, 16'h0055, 16'h0056, 16'h0057 	:	val_out <= 16'h80fb;
         16'h0058, 16'h0059, 16'h005a, 16'h005b, 16'h005c, 16'h005d, 16'h005e, 16'h005f 	:	val_out <= 16'h8114;
         16'h0060, 16'h0061, 16'h0062, 16'h0063, 16'h0064, 16'h0065, 16'h0066, 16'h0067 	:	val_out <= 16'h812d;
         16'h0068, 16'h0069, 16'h006a, 16'h006b, 16'h006c, 16'h006d, 16'h006e, 16'h006f 	:	val_out <= 16'h8146;
         16'h0070, 16'h0071, 16'h0072, 16'h0073, 16'h0074, 16'h0075, 16'h0076, 16'h0077 	:	val_out <= 16'h815f;
         16'h0078, 16'h0079, 16'h007a, 16'h007b, 16'h007c, 16'h007d, 16'h007e, 16'h007f 	:	val_out <= 16'h8178;
         16'h0080, 16'h0081, 16'h0082, 16'h0083, 16'h0084, 16'h0085, 16'h0086, 16'h0087 	:	val_out <= 16'h8192;
         16'h0088, 16'h0089, 16'h008a, 16'h008b, 16'h008c, 16'h008d, 16'h008e, 16'h008f 	:	val_out <= 16'h81ab;
         16'h0090, 16'h0091, 16'h0092, 16'h0093, 16'h0094, 16'h0095, 16'h0096, 16'h0097 	:	val_out <= 16'h81c4;
         16'h0098, 16'h0099, 16'h009a, 16'h009b, 16'h009c, 16'h009d, 16'h009e, 16'h009f 	:	val_out <= 16'h81dd;
         16'h00a0, 16'h00a1, 16'h00a2, 16'h00a3, 16'h00a4, 16'h00a5, 16'h00a6, 16'h00a7 	:	val_out <= 16'h81f6;
         16'h00a8, 16'h00a9, 16'h00aa, 16'h00ab, 16'h00ac, 16'h00ad, 16'h00ae, 16'h00af 	:	val_out <= 16'h820f;
         16'h00b0, 16'h00b1, 16'h00b2, 16'h00b3, 16'h00b4, 16'h00b5, 16'h00b6, 16'h00b7 	:	val_out <= 16'h8228;
         16'h00b8, 16'h00b9, 16'h00ba, 16'h00bb, 16'h00bc, 16'h00bd, 16'h00be, 16'h00bf 	:	val_out <= 16'h8242;
         16'h00c0, 16'h00c1, 16'h00c2, 16'h00c3, 16'h00c4, 16'h00c5, 16'h00c6, 16'h00c7 	:	val_out <= 16'h825b;
         16'h00c8, 16'h00c9, 16'h00ca, 16'h00cb, 16'h00cc, 16'h00cd, 16'h00ce, 16'h00cf 	:	val_out <= 16'h8274;
         16'h00d0, 16'h00d1, 16'h00d2, 16'h00d3, 16'h00d4, 16'h00d5, 16'h00d6, 16'h00d7 	:	val_out <= 16'h828d;
         16'h00d8, 16'h00d9, 16'h00da, 16'h00db, 16'h00dc, 16'h00dd, 16'h00de, 16'h00df 	:	val_out <= 16'h82a6;
         16'h00e0, 16'h00e1, 16'h00e2, 16'h00e3, 16'h00e4, 16'h00e5, 16'h00e6, 16'h00e7 	:	val_out <= 16'h82bf;
         16'h00e8, 16'h00e9, 16'h00ea, 16'h00eb, 16'h00ec, 16'h00ed, 16'h00ee, 16'h00ef 	:	val_out <= 16'h82d8;
         16'h00f0, 16'h00f1, 16'h00f2, 16'h00f3, 16'h00f4, 16'h00f5, 16'h00f6, 16'h00f7 	:	val_out <= 16'h82f1;
         16'h00f8, 16'h00f9, 16'h00fa, 16'h00fb, 16'h00fc, 16'h00fd, 16'h00fe, 16'h00ff 	:	val_out <= 16'h830b;
         16'h0100, 16'h0101, 16'h0102, 16'h0103, 16'h0104, 16'h0105, 16'h0106, 16'h0107 	:	val_out <= 16'h8324;
         16'h0108, 16'h0109, 16'h010a, 16'h010b, 16'h010c, 16'h010d, 16'h010e, 16'h010f 	:	val_out <= 16'h833d;
         16'h0110, 16'h0111, 16'h0112, 16'h0113, 16'h0114, 16'h0115, 16'h0116, 16'h0117 	:	val_out <= 16'h8356;
         16'h0118, 16'h0119, 16'h011a, 16'h011b, 16'h011c, 16'h011d, 16'h011e, 16'h011f 	:	val_out <= 16'h836f;
         16'h0120, 16'h0121, 16'h0122, 16'h0123, 16'h0124, 16'h0125, 16'h0126, 16'h0127 	:	val_out <= 16'h8388;
         16'h0128, 16'h0129, 16'h012a, 16'h012b, 16'h012c, 16'h012d, 16'h012e, 16'h012f 	:	val_out <= 16'h83a1;
         16'h0130, 16'h0131, 16'h0132, 16'h0133, 16'h0134, 16'h0135, 16'h0136, 16'h0137 	:	val_out <= 16'h83ba;
         16'h0138, 16'h0139, 16'h013a, 16'h013b, 16'h013c, 16'h013d, 16'h013e, 16'h013f 	:	val_out <= 16'h83d4;
         16'h0140, 16'h0141, 16'h0142, 16'h0143, 16'h0144, 16'h0145, 16'h0146, 16'h0147 	:	val_out <= 16'h83ed;
         16'h0148, 16'h0149, 16'h014a, 16'h014b, 16'h014c, 16'h014d, 16'h014e, 16'h014f 	:	val_out <= 16'h8406;
         16'h0150, 16'h0151, 16'h0152, 16'h0153, 16'h0154, 16'h0155, 16'h0156, 16'h0157 	:	val_out <= 16'h841f;
         16'h0158, 16'h0159, 16'h015a, 16'h015b, 16'h015c, 16'h015d, 16'h015e, 16'h015f 	:	val_out <= 16'h8438;
         16'h0160, 16'h0161, 16'h0162, 16'h0163, 16'h0164, 16'h0165, 16'h0166, 16'h0167 	:	val_out <= 16'h8451;
         16'h0168, 16'h0169, 16'h016a, 16'h016b, 16'h016c, 16'h016d, 16'h016e, 16'h016f 	:	val_out <= 16'h846a;
         16'h0170, 16'h0171, 16'h0172, 16'h0173, 16'h0174, 16'h0175, 16'h0176, 16'h0177 	:	val_out <= 16'h8483;
         16'h0178, 16'h0179, 16'h017a, 16'h017b, 16'h017c, 16'h017d, 16'h017e, 16'h017f 	:	val_out <= 16'h849c;
         16'h0180, 16'h0181, 16'h0182, 16'h0183, 16'h0184, 16'h0185, 16'h0186, 16'h0187 	:	val_out <= 16'h84b6;
         16'h0188, 16'h0189, 16'h018a, 16'h018b, 16'h018c, 16'h018d, 16'h018e, 16'h018f 	:	val_out <= 16'h84cf;
         16'h0190, 16'h0191, 16'h0192, 16'h0193, 16'h0194, 16'h0195, 16'h0196, 16'h0197 	:	val_out <= 16'h84e8;
         16'h0198, 16'h0199, 16'h019a, 16'h019b, 16'h019c, 16'h019d, 16'h019e, 16'h019f 	:	val_out <= 16'h8501;
         16'h01a0, 16'h01a1, 16'h01a2, 16'h01a3, 16'h01a4, 16'h01a5, 16'h01a6, 16'h01a7 	:	val_out <= 16'h851a;
         16'h01a8, 16'h01a9, 16'h01aa, 16'h01ab, 16'h01ac, 16'h01ad, 16'h01ae, 16'h01af 	:	val_out <= 16'h8533;
         16'h01b0, 16'h01b1, 16'h01b2, 16'h01b3, 16'h01b4, 16'h01b5, 16'h01b6, 16'h01b7 	:	val_out <= 16'h854c;
         16'h01b8, 16'h01b9, 16'h01ba, 16'h01bb, 16'h01bc, 16'h01bd, 16'h01be, 16'h01bf 	:	val_out <= 16'h8565;
         16'h01c0, 16'h01c1, 16'h01c2, 16'h01c3, 16'h01c4, 16'h01c5, 16'h01c6, 16'h01c7 	:	val_out <= 16'h857f;
         16'h01c8, 16'h01c9, 16'h01ca, 16'h01cb, 16'h01cc, 16'h01cd, 16'h01ce, 16'h01cf 	:	val_out <= 16'h8598;
         16'h01d0, 16'h01d1, 16'h01d2, 16'h01d3, 16'h01d4, 16'h01d5, 16'h01d6, 16'h01d7 	:	val_out <= 16'h85b1;
         16'h01d8, 16'h01d9, 16'h01da, 16'h01db, 16'h01dc, 16'h01dd, 16'h01de, 16'h01df 	:	val_out <= 16'h85ca;
         16'h01e0, 16'h01e1, 16'h01e2, 16'h01e3, 16'h01e4, 16'h01e5, 16'h01e6, 16'h01e7 	:	val_out <= 16'h85e3;
         16'h01e8, 16'h01e9, 16'h01ea, 16'h01eb, 16'h01ec, 16'h01ed, 16'h01ee, 16'h01ef 	:	val_out <= 16'h85fc;
         16'h01f0, 16'h01f1, 16'h01f2, 16'h01f3, 16'h01f4, 16'h01f5, 16'h01f6, 16'h01f7 	:	val_out <= 16'h8615;
         16'h01f8, 16'h01f9, 16'h01fa, 16'h01fb, 16'h01fc, 16'h01fd, 16'h01fe, 16'h01ff 	:	val_out <= 16'h862e;
         16'h0200, 16'h0201, 16'h0202, 16'h0203, 16'h0204, 16'h0205, 16'h0206, 16'h0207 	:	val_out <= 16'h8647;
         16'h0208, 16'h0209, 16'h020a, 16'h020b, 16'h020c, 16'h020d, 16'h020e, 16'h020f 	:	val_out <= 16'h8660;
         16'h0210, 16'h0211, 16'h0212, 16'h0213, 16'h0214, 16'h0215, 16'h0216, 16'h0217 	:	val_out <= 16'h867a;
         16'h0218, 16'h0219, 16'h021a, 16'h021b, 16'h021c, 16'h021d, 16'h021e, 16'h021f 	:	val_out <= 16'h8693;
         16'h0220, 16'h0221, 16'h0222, 16'h0223, 16'h0224, 16'h0225, 16'h0226, 16'h0227 	:	val_out <= 16'h86ac;
         16'h0228, 16'h0229, 16'h022a, 16'h022b, 16'h022c, 16'h022d, 16'h022e, 16'h022f 	:	val_out <= 16'h86c5;
         16'h0230, 16'h0231, 16'h0232, 16'h0233, 16'h0234, 16'h0235, 16'h0236, 16'h0237 	:	val_out <= 16'h86de;
         16'h0238, 16'h0239, 16'h023a, 16'h023b, 16'h023c, 16'h023d, 16'h023e, 16'h023f 	:	val_out <= 16'h86f7;
         16'h0240, 16'h0241, 16'h0242, 16'h0243, 16'h0244, 16'h0245, 16'h0246, 16'h0247 	:	val_out <= 16'h8710;
         16'h0248, 16'h0249, 16'h024a, 16'h024b, 16'h024c, 16'h024d, 16'h024e, 16'h024f 	:	val_out <= 16'h8729;
         16'h0250, 16'h0251, 16'h0252, 16'h0253, 16'h0254, 16'h0255, 16'h0256, 16'h0257 	:	val_out <= 16'h8742;
         16'h0258, 16'h0259, 16'h025a, 16'h025b, 16'h025c, 16'h025d, 16'h025e, 16'h025f 	:	val_out <= 16'h875b;
         16'h0260, 16'h0261, 16'h0262, 16'h0263, 16'h0264, 16'h0265, 16'h0266, 16'h0267 	:	val_out <= 16'h8775;
         16'h0268, 16'h0269, 16'h026a, 16'h026b, 16'h026c, 16'h026d, 16'h026e, 16'h026f 	:	val_out <= 16'h878e;
         16'h0270, 16'h0271, 16'h0272, 16'h0273, 16'h0274, 16'h0275, 16'h0276, 16'h0277 	:	val_out <= 16'h87a7;
         16'h0278, 16'h0279, 16'h027a, 16'h027b, 16'h027c, 16'h027d, 16'h027e, 16'h027f 	:	val_out <= 16'h87c0;
         16'h0280, 16'h0281, 16'h0282, 16'h0283, 16'h0284, 16'h0285, 16'h0286, 16'h0287 	:	val_out <= 16'h87d9;
         16'h0288, 16'h0289, 16'h028a, 16'h028b, 16'h028c, 16'h028d, 16'h028e, 16'h028f 	:	val_out <= 16'h87f2;
         16'h0290, 16'h0291, 16'h0292, 16'h0293, 16'h0294, 16'h0295, 16'h0296, 16'h0297 	:	val_out <= 16'h880b;
         16'h0298, 16'h0299, 16'h029a, 16'h029b, 16'h029c, 16'h029d, 16'h029e, 16'h029f 	:	val_out <= 16'h8824;
         16'h02a0, 16'h02a1, 16'h02a2, 16'h02a3, 16'h02a4, 16'h02a5, 16'h02a6, 16'h02a7 	:	val_out <= 16'h883d;
         16'h02a8, 16'h02a9, 16'h02aa, 16'h02ab, 16'h02ac, 16'h02ad, 16'h02ae, 16'h02af 	:	val_out <= 16'h8856;
         16'h02b0, 16'h02b1, 16'h02b2, 16'h02b3, 16'h02b4, 16'h02b5, 16'h02b6, 16'h02b7 	:	val_out <= 16'h886f;
         16'h02b8, 16'h02b9, 16'h02ba, 16'h02bb, 16'h02bc, 16'h02bd, 16'h02be, 16'h02bf 	:	val_out <= 16'h8888;
         16'h02c0, 16'h02c1, 16'h02c2, 16'h02c3, 16'h02c4, 16'h02c5, 16'h02c6, 16'h02c7 	:	val_out <= 16'h88a2;
         16'h02c8, 16'h02c9, 16'h02ca, 16'h02cb, 16'h02cc, 16'h02cd, 16'h02ce, 16'h02cf 	:	val_out <= 16'h88bb;
         16'h02d0, 16'h02d1, 16'h02d2, 16'h02d3, 16'h02d4, 16'h02d5, 16'h02d6, 16'h02d7 	:	val_out <= 16'h88d4;
         16'h02d8, 16'h02d9, 16'h02da, 16'h02db, 16'h02dc, 16'h02dd, 16'h02de, 16'h02df 	:	val_out <= 16'h88ed;
         16'h02e0, 16'h02e1, 16'h02e2, 16'h02e3, 16'h02e4, 16'h02e5, 16'h02e6, 16'h02e7 	:	val_out <= 16'h8906;
         16'h02e8, 16'h02e9, 16'h02ea, 16'h02eb, 16'h02ec, 16'h02ed, 16'h02ee, 16'h02ef 	:	val_out <= 16'h891f;
         16'h02f0, 16'h02f1, 16'h02f2, 16'h02f3, 16'h02f4, 16'h02f5, 16'h02f6, 16'h02f7 	:	val_out <= 16'h8938;
         16'h02f8, 16'h02f9, 16'h02fa, 16'h02fb, 16'h02fc, 16'h02fd, 16'h02fe, 16'h02ff 	:	val_out <= 16'h8951;
         16'h0300, 16'h0301, 16'h0302, 16'h0303, 16'h0304, 16'h0305, 16'h0306, 16'h0307 	:	val_out <= 16'h896a;
         16'h0308, 16'h0309, 16'h030a, 16'h030b, 16'h030c, 16'h030d, 16'h030e, 16'h030f 	:	val_out <= 16'h8983;
         16'h0310, 16'h0311, 16'h0312, 16'h0313, 16'h0314, 16'h0315, 16'h0316, 16'h0317 	:	val_out <= 16'h899c;
         16'h0318, 16'h0319, 16'h031a, 16'h031b, 16'h031c, 16'h031d, 16'h031e, 16'h031f 	:	val_out <= 16'h89b5;
         16'h0320, 16'h0321, 16'h0322, 16'h0323, 16'h0324, 16'h0325, 16'h0326, 16'h0327 	:	val_out <= 16'h89ce;
         16'h0328, 16'h0329, 16'h032a, 16'h032b, 16'h032c, 16'h032d, 16'h032e, 16'h032f 	:	val_out <= 16'h89e7;
         16'h0330, 16'h0331, 16'h0332, 16'h0333, 16'h0334, 16'h0335, 16'h0336, 16'h0337 	:	val_out <= 16'h8a00;
         16'h0338, 16'h0339, 16'h033a, 16'h033b, 16'h033c, 16'h033d, 16'h033e, 16'h033f 	:	val_out <= 16'h8a19;
         16'h0340, 16'h0341, 16'h0342, 16'h0343, 16'h0344, 16'h0345, 16'h0346, 16'h0347 	:	val_out <= 16'h8a33;
         16'h0348, 16'h0349, 16'h034a, 16'h034b, 16'h034c, 16'h034d, 16'h034e, 16'h034f 	:	val_out <= 16'h8a4c;
         16'h0350, 16'h0351, 16'h0352, 16'h0353, 16'h0354, 16'h0355, 16'h0356, 16'h0357 	:	val_out <= 16'h8a65;
         16'h0358, 16'h0359, 16'h035a, 16'h035b, 16'h035c, 16'h035d, 16'h035e, 16'h035f 	:	val_out <= 16'h8a7e;
         16'h0360, 16'h0361, 16'h0362, 16'h0363, 16'h0364, 16'h0365, 16'h0366, 16'h0367 	:	val_out <= 16'h8a97;
         16'h0368, 16'h0369, 16'h036a, 16'h036b, 16'h036c, 16'h036d, 16'h036e, 16'h036f 	:	val_out <= 16'h8ab0;
         16'h0370, 16'h0371, 16'h0372, 16'h0373, 16'h0374, 16'h0375, 16'h0376, 16'h0377 	:	val_out <= 16'h8ac9;
         16'h0378, 16'h0379, 16'h037a, 16'h037b, 16'h037c, 16'h037d, 16'h037e, 16'h037f 	:	val_out <= 16'h8ae2;
         16'h0380, 16'h0381, 16'h0382, 16'h0383, 16'h0384, 16'h0385, 16'h0386, 16'h0387 	:	val_out <= 16'h8afb;
         16'h0388, 16'h0389, 16'h038a, 16'h038b, 16'h038c, 16'h038d, 16'h038e, 16'h038f 	:	val_out <= 16'h8b14;
         16'h0390, 16'h0391, 16'h0392, 16'h0393, 16'h0394, 16'h0395, 16'h0396, 16'h0397 	:	val_out <= 16'h8b2d;
         16'h0398, 16'h0399, 16'h039a, 16'h039b, 16'h039c, 16'h039d, 16'h039e, 16'h039f 	:	val_out <= 16'h8b46;
         16'h03a0, 16'h03a1, 16'h03a2, 16'h03a3, 16'h03a4, 16'h03a5, 16'h03a6, 16'h03a7 	:	val_out <= 16'h8b5f;
         16'h03a8, 16'h03a9, 16'h03aa, 16'h03ab, 16'h03ac, 16'h03ad, 16'h03ae, 16'h03af 	:	val_out <= 16'h8b78;
         16'h03b0, 16'h03b1, 16'h03b2, 16'h03b3, 16'h03b4, 16'h03b5, 16'h03b6, 16'h03b7 	:	val_out <= 16'h8b91;
         16'h03b8, 16'h03b9, 16'h03ba, 16'h03bb, 16'h03bc, 16'h03bd, 16'h03be, 16'h03bf 	:	val_out <= 16'h8baa;
         16'h03c0, 16'h03c1, 16'h03c2, 16'h03c3, 16'h03c4, 16'h03c5, 16'h03c6, 16'h03c7 	:	val_out <= 16'h8bc3;
         16'h03c8, 16'h03c9, 16'h03ca, 16'h03cb, 16'h03cc, 16'h03cd, 16'h03ce, 16'h03cf 	:	val_out <= 16'h8bdc;
         16'h03d0, 16'h03d1, 16'h03d2, 16'h03d3, 16'h03d4, 16'h03d5, 16'h03d6, 16'h03d7 	:	val_out <= 16'h8bf5;
         16'h03d8, 16'h03d9, 16'h03da, 16'h03db, 16'h03dc, 16'h03dd, 16'h03de, 16'h03df 	:	val_out <= 16'h8c0e;
         16'h03e0, 16'h03e1, 16'h03e2, 16'h03e3, 16'h03e4, 16'h03e5, 16'h03e6, 16'h03e7 	:	val_out <= 16'h8c27;
         16'h03e8, 16'h03e9, 16'h03ea, 16'h03eb, 16'h03ec, 16'h03ed, 16'h03ee, 16'h03ef 	:	val_out <= 16'h8c40;
         16'h03f0, 16'h03f1, 16'h03f2, 16'h03f3, 16'h03f4, 16'h03f5, 16'h03f6, 16'h03f7 	:	val_out <= 16'h8c59;
         16'h03f8, 16'h03f9, 16'h03fa, 16'h03fb, 16'h03fc, 16'h03fd, 16'h03fe, 16'h03ff 	:	val_out <= 16'h8c72;
         16'h0400, 16'h0401, 16'h0402, 16'h0403, 16'h0404, 16'h0405, 16'h0406, 16'h0407 	:	val_out <= 16'h8c8b;
         16'h0408, 16'h0409, 16'h040a, 16'h040b, 16'h040c, 16'h040d, 16'h040e, 16'h040f 	:	val_out <= 16'h8ca4;
         16'h0410, 16'h0411, 16'h0412, 16'h0413, 16'h0414, 16'h0415, 16'h0416, 16'h0417 	:	val_out <= 16'h8cbd;
         16'h0418, 16'h0419, 16'h041a, 16'h041b, 16'h041c, 16'h041d, 16'h041e, 16'h041f 	:	val_out <= 16'h8cd6;
         16'h0420, 16'h0421, 16'h0422, 16'h0423, 16'h0424, 16'h0425, 16'h0426, 16'h0427 	:	val_out <= 16'h8cef;
         16'h0428, 16'h0429, 16'h042a, 16'h042b, 16'h042c, 16'h042d, 16'h042e, 16'h042f 	:	val_out <= 16'h8d08;
         16'h0430, 16'h0431, 16'h0432, 16'h0433, 16'h0434, 16'h0435, 16'h0436, 16'h0437 	:	val_out <= 16'h8d21;
         16'h0438, 16'h0439, 16'h043a, 16'h043b, 16'h043c, 16'h043d, 16'h043e, 16'h043f 	:	val_out <= 16'h8d3a;
         16'h0440, 16'h0441, 16'h0442, 16'h0443, 16'h0444, 16'h0445, 16'h0446, 16'h0447 	:	val_out <= 16'h8d53;
         16'h0448, 16'h0449, 16'h044a, 16'h044b, 16'h044c, 16'h044d, 16'h044e, 16'h044f 	:	val_out <= 16'h8d6c;
         16'h0450, 16'h0451, 16'h0452, 16'h0453, 16'h0454, 16'h0455, 16'h0456, 16'h0457 	:	val_out <= 16'h8d85;
         16'h0458, 16'h0459, 16'h045a, 16'h045b, 16'h045c, 16'h045d, 16'h045e, 16'h045f 	:	val_out <= 16'h8d9e;
         16'h0460, 16'h0461, 16'h0462, 16'h0463, 16'h0464, 16'h0465, 16'h0466, 16'h0467 	:	val_out <= 16'h8db7;
         16'h0468, 16'h0469, 16'h046a, 16'h046b, 16'h046c, 16'h046d, 16'h046e, 16'h046f 	:	val_out <= 16'h8dd0;
         16'h0470, 16'h0471, 16'h0472, 16'h0473, 16'h0474, 16'h0475, 16'h0476, 16'h0477 	:	val_out <= 16'h8de9;
         16'h0478, 16'h0479, 16'h047a, 16'h047b, 16'h047c, 16'h047d, 16'h047e, 16'h047f 	:	val_out <= 16'h8e02;
         16'h0480, 16'h0481, 16'h0482, 16'h0483, 16'h0484, 16'h0485, 16'h0486, 16'h0487 	:	val_out <= 16'h8e1b;
         16'h0488, 16'h0489, 16'h048a, 16'h048b, 16'h048c, 16'h048d, 16'h048e, 16'h048f 	:	val_out <= 16'h8e34;
         16'h0490, 16'h0491, 16'h0492, 16'h0493, 16'h0494, 16'h0495, 16'h0496, 16'h0497 	:	val_out <= 16'h8e4d;
         16'h0498, 16'h0499, 16'h049a, 16'h049b, 16'h049c, 16'h049d, 16'h049e, 16'h049f 	:	val_out <= 16'h8e66;
         16'h04a0, 16'h04a1, 16'h04a2, 16'h04a3, 16'h04a4, 16'h04a5, 16'h04a6, 16'h04a7 	:	val_out <= 16'h8e7f;
         16'h04a8, 16'h04a9, 16'h04aa, 16'h04ab, 16'h04ac, 16'h04ad, 16'h04ae, 16'h04af 	:	val_out <= 16'h8e98;
         16'h04b0, 16'h04b1, 16'h04b2, 16'h04b3, 16'h04b4, 16'h04b5, 16'h04b6, 16'h04b7 	:	val_out <= 16'h8eb1;
         16'h04b8, 16'h04b9, 16'h04ba, 16'h04bb, 16'h04bc, 16'h04bd, 16'h04be, 16'h04bf 	:	val_out <= 16'h8eca;
         16'h04c0, 16'h04c1, 16'h04c2, 16'h04c3, 16'h04c4, 16'h04c5, 16'h04c6, 16'h04c7 	:	val_out <= 16'h8ee3;
         16'h04c8, 16'h04c9, 16'h04ca, 16'h04cb, 16'h04cc, 16'h04cd, 16'h04ce, 16'h04cf 	:	val_out <= 16'h8efc;
         16'h04d0, 16'h04d1, 16'h04d2, 16'h04d3, 16'h04d4, 16'h04d5, 16'h04d6, 16'h04d7 	:	val_out <= 16'h8f15;
         16'h04d8, 16'h04d9, 16'h04da, 16'h04db, 16'h04dc, 16'h04dd, 16'h04de, 16'h04df 	:	val_out <= 16'h8f2e;
         16'h04e0, 16'h04e1, 16'h04e2, 16'h04e3, 16'h04e4, 16'h04e5, 16'h04e6, 16'h04e7 	:	val_out <= 16'h8f47;
         16'h04e8, 16'h04e9, 16'h04ea, 16'h04eb, 16'h04ec, 16'h04ed, 16'h04ee, 16'h04ef 	:	val_out <= 16'h8f60;
         16'h04f0, 16'h04f1, 16'h04f2, 16'h04f3, 16'h04f4, 16'h04f5, 16'h04f6, 16'h04f7 	:	val_out <= 16'h8f79;
         16'h04f8, 16'h04f9, 16'h04fa, 16'h04fb, 16'h04fc, 16'h04fd, 16'h04fe, 16'h04ff 	:	val_out <= 16'h8f92;
         16'h0500, 16'h0501, 16'h0502, 16'h0503, 16'h0504, 16'h0505, 16'h0506, 16'h0507 	:	val_out <= 16'h8fab;
         16'h0508, 16'h0509, 16'h050a, 16'h050b, 16'h050c, 16'h050d, 16'h050e, 16'h050f 	:	val_out <= 16'h8fc4;
         16'h0510, 16'h0511, 16'h0512, 16'h0513, 16'h0514, 16'h0515, 16'h0516, 16'h0517 	:	val_out <= 16'h8fdd;
         16'h0518, 16'h0519, 16'h051a, 16'h051b, 16'h051c, 16'h051d, 16'h051e, 16'h051f 	:	val_out <= 16'h8ff5;
         16'h0520, 16'h0521, 16'h0522, 16'h0523, 16'h0524, 16'h0525, 16'h0526, 16'h0527 	:	val_out <= 16'h900e;
         16'h0528, 16'h0529, 16'h052a, 16'h052b, 16'h052c, 16'h052d, 16'h052e, 16'h052f 	:	val_out <= 16'h9027;
         16'h0530, 16'h0531, 16'h0532, 16'h0533, 16'h0534, 16'h0535, 16'h0536, 16'h0537 	:	val_out <= 16'h9040;
         16'h0538, 16'h0539, 16'h053a, 16'h053b, 16'h053c, 16'h053d, 16'h053e, 16'h053f 	:	val_out <= 16'h9059;
         16'h0540, 16'h0541, 16'h0542, 16'h0543, 16'h0544, 16'h0545, 16'h0546, 16'h0547 	:	val_out <= 16'h9072;
         16'h0548, 16'h0549, 16'h054a, 16'h054b, 16'h054c, 16'h054d, 16'h054e, 16'h054f 	:	val_out <= 16'h908b;
         16'h0550, 16'h0551, 16'h0552, 16'h0553, 16'h0554, 16'h0555, 16'h0556, 16'h0557 	:	val_out <= 16'h90a4;
         16'h0558, 16'h0559, 16'h055a, 16'h055b, 16'h055c, 16'h055d, 16'h055e, 16'h055f 	:	val_out <= 16'h90bd;
         16'h0560, 16'h0561, 16'h0562, 16'h0563, 16'h0564, 16'h0565, 16'h0566, 16'h0567 	:	val_out <= 16'h90d6;
         16'h0568, 16'h0569, 16'h056a, 16'h056b, 16'h056c, 16'h056d, 16'h056e, 16'h056f 	:	val_out <= 16'h90ef;
         16'h0570, 16'h0571, 16'h0572, 16'h0573, 16'h0574, 16'h0575, 16'h0576, 16'h0577 	:	val_out <= 16'h9108;
         16'h0578, 16'h0579, 16'h057a, 16'h057b, 16'h057c, 16'h057d, 16'h057e, 16'h057f 	:	val_out <= 16'h9121;
         16'h0580, 16'h0581, 16'h0582, 16'h0583, 16'h0584, 16'h0585, 16'h0586, 16'h0587 	:	val_out <= 16'h9139;
         16'h0588, 16'h0589, 16'h058a, 16'h058b, 16'h058c, 16'h058d, 16'h058e, 16'h058f 	:	val_out <= 16'h9152;
         16'h0590, 16'h0591, 16'h0592, 16'h0593, 16'h0594, 16'h0595, 16'h0596, 16'h0597 	:	val_out <= 16'h916b;
         16'h0598, 16'h0599, 16'h059a, 16'h059b, 16'h059c, 16'h059d, 16'h059e, 16'h059f 	:	val_out <= 16'h9184;
         16'h05a0, 16'h05a1, 16'h05a2, 16'h05a3, 16'h05a4, 16'h05a5, 16'h05a6, 16'h05a7 	:	val_out <= 16'h919d;
         16'h05a8, 16'h05a9, 16'h05aa, 16'h05ab, 16'h05ac, 16'h05ad, 16'h05ae, 16'h05af 	:	val_out <= 16'h91b6;
         16'h05b0, 16'h05b1, 16'h05b2, 16'h05b3, 16'h05b4, 16'h05b5, 16'h05b6, 16'h05b7 	:	val_out <= 16'h91cf;
         16'h05b8, 16'h05b9, 16'h05ba, 16'h05bb, 16'h05bc, 16'h05bd, 16'h05be, 16'h05bf 	:	val_out <= 16'h91e8;
         16'h05c0, 16'h05c1, 16'h05c2, 16'h05c3, 16'h05c4, 16'h05c5, 16'h05c6, 16'h05c7 	:	val_out <= 16'h9201;
         16'h05c8, 16'h05c9, 16'h05ca, 16'h05cb, 16'h05cc, 16'h05cd, 16'h05ce, 16'h05cf 	:	val_out <= 16'h9219;
         16'h05d0, 16'h05d1, 16'h05d2, 16'h05d3, 16'h05d4, 16'h05d5, 16'h05d6, 16'h05d7 	:	val_out <= 16'h9232;
         16'h05d8, 16'h05d9, 16'h05da, 16'h05db, 16'h05dc, 16'h05dd, 16'h05de, 16'h05df 	:	val_out <= 16'h924b;
         16'h05e0, 16'h05e1, 16'h05e2, 16'h05e3, 16'h05e4, 16'h05e5, 16'h05e6, 16'h05e7 	:	val_out <= 16'h9264;
         16'h05e8, 16'h05e9, 16'h05ea, 16'h05eb, 16'h05ec, 16'h05ed, 16'h05ee, 16'h05ef 	:	val_out <= 16'h927d;
         16'h05f0, 16'h05f1, 16'h05f2, 16'h05f3, 16'h05f4, 16'h05f5, 16'h05f6, 16'h05f7 	:	val_out <= 16'h9296;
         16'h05f8, 16'h05f9, 16'h05fa, 16'h05fb, 16'h05fc, 16'h05fd, 16'h05fe, 16'h05ff 	:	val_out <= 16'h92af;
         16'h0600, 16'h0601, 16'h0602, 16'h0603, 16'h0604, 16'h0605, 16'h0606, 16'h0607 	:	val_out <= 16'h92c8;
         16'h0608, 16'h0609, 16'h060a, 16'h060b, 16'h060c, 16'h060d, 16'h060e, 16'h060f 	:	val_out <= 16'h92e0;
         16'h0610, 16'h0611, 16'h0612, 16'h0613, 16'h0614, 16'h0615, 16'h0616, 16'h0617 	:	val_out <= 16'h92f9;
         16'h0618, 16'h0619, 16'h061a, 16'h061b, 16'h061c, 16'h061d, 16'h061e, 16'h061f 	:	val_out <= 16'h9312;
         16'h0620, 16'h0621, 16'h0622, 16'h0623, 16'h0624, 16'h0625, 16'h0626, 16'h0627 	:	val_out <= 16'h932b;
         16'h0628, 16'h0629, 16'h062a, 16'h062b, 16'h062c, 16'h062d, 16'h062e, 16'h062f 	:	val_out <= 16'h9344;
         16'h0630, 16'h0631, 16'h0632, 16'h0633, 16'h0634, 16'h0635, 16'h0636, 16'h0637 	:	val_out <= 16'h935d;
         16'h0638, 16'h0639, 16'h063a, 16'h063b, 16'h063c, 16'h063d, 16'h063e, 16'h063f 	:	val_out <= 16'h9376;
         16'h0640, 16'h0641, 16'h0642, 16'h0643, 16'h0644, 16'h0645, 16'h0646, 16'h0647 	:	val_out <= 16'h938e;
         16'h0648, 16'h0649, 16'h064a, 16'h064b, 16'h064c, 16'h064d, 16'h064e, 16'h064f 	:	val_out <= 16'h93a7;
         16'h0650, 16'h0651, 16'h0652, 16'h0653, 16'h0654, 16'h0655, 16'h0656, 16'h0657 	:	val_out <= 16'h93c0;
         16'h0658, 16'h0659, 16'h065a, 16'h065b, 16'h065c, 16'h065d, 16'h065e, 16'h065f 	:	val_out <= 16'h93d9;
         16'h0660, 16'h0661, 16'h0662, 16'h0663, 16'h0664, 16'h0665, 16'h0666, 16'h0667 	:	val_out <= 16'h93f2;
         16'h0668, 16'h0669, 16'h066a, 16'h066b, 16'h066c, 16'h066d, 16'h066e, 16'h066f 	:	val_out <= 16'h940b;
         16'h0670, 16'h0671, 16'h0672, 16'h0673, 16'h0674, 16'h0675, 16'h0676, 16'h0677 	:	val_out <= 16'h9423;
         16'h0678, 16'h0679, 16'h067a, 16'h067b, 16'h067c, 16'h067d, 16'h067e, 16'h067f 	:	val_out <= 16'h943c;
         16'h0680, 16'h0681, 16'h0682, 16'h0683, 16'h0684, 16'h0685, 16'h0686, 16'h0687 	:	val_out <= 16'h9455;
         16'h0688, 16'h0689, 16'h068a, 16'h068b, 16'h068c, 16'h068d, 16'h068e, 16'h068f 	:	val_out <= 16'h946e;
         16'h0690, 16'h0691, 16'h0692, 16'h0693, 16'h0694, 16'h0695, 16'h0696, 16'h0697 	:	val_out <= 16'h9487;
         16'h0698, 16'h0699, 16'h069a, 16'h069b, 16'h069c, 16'h069d, 16'h069e, 16'h069f 	:	val_out <= 16'h949f;
         16'h06a0, 16'h06a1, 16'h06a2, 16'h06a3, 16'h06a4, 16'h06a5, 16'h06a6, 16'h06a7 	:	val_out <= 16'h94b8;
         16'h06a8, 16'h06a9, 16'h06aa, 16'h06ab, 16'h06ac, 16'h06ad, 16'h06ae, 16'h06af 	:	val_out <= 16'h94d1;
         16'h06b0, 16'h06b1, 16'h06b2, 16'h06b3, 16'h06b4, 16'h06b5, 16'h06b6, 16'h06b7 	:	val_out <= 16'h94ea;
         16'h06b8, 16'h06b9, 16'h06ba, 16'h06bb, 16'h06bc, 16'h06bd, 16'h06be, 16'h06bf 	:	val_out <= 16'h9503;
         16'h06c0, 16'h06c1, 16'h06c2, 16'h06c3, 16'h06c4, 16'h06c5, 16'h06c6, 16'h06c7 	:	val_out <= 16'h951b;
         16'h06c8, 16'h06c9, 16'h06ca, 16'h06cb, 16'h06cc, 16'h06cd, 16'h06ce, 16'h06cf 	:	val_out <= 16'h9534;
         16'h06d0, 16'h06d1, 16'h06d2, 16'h06d3, 16'h06d4, 16'h06d5, 16'h06d6, 16'h06d7 	:	val_out <= 16'h954d;
         16'h06d8, 16'h06d9, 16'h06da, 16'h06db, 16'h06dc, 16'h06dd, 16'h06de, 16'h06df 	:	val_out <= 16'h9566;
         16'h06e0, 16'h06e1, 16'h06e2, 16'h06e3, 16'h06e4, 16'h06e5, 16'h06e6, 16'h06e7 	:	val_out <= 16'h957f;
         16'h06e8, 16'h06e9, 16'h06ea, 16'h06eb, 16'h06ec, 16'h06ed, 16'h06ee, 16'h06ef 	:	val_out <= 16'h9597;
         16'h06f0, 16'h06f1, 16'h06f2, 16'h06f3, 16'h06f4, 16'h06f5, 16'h06f6, 16'h06f7 	:	val_out <= 16'h95b0;
         16'h06f8, 16'h06f9, 16'h06fa, 16'h06fb, 16'h06fc, 16'h06fd, 16'h06fe, 16'h06ff 	:	val_out <= 16'h95c9;
         16'h0700, 16'h0701, 16'h0702, 16'h0703, 16'h0704, 16'h0705, 16'h0706, 16'h0707 	:	val_out <= 16'h95e2;
         16'h0708, 16'h0709, 16'h070a, 16'h070b, 16'h070c, 16'h070d, 16'h070e, 16'h070f 	:	val_out <= 16'h95fa;
         16'h0710, 16'h0711, 16'h0712, 16'h0713, 16'h0714, 16'h0715, 16'h0716, 16'h0717 	:	val_out <= 16'h9613;
         16'h0718, 16'h0719, 16'h071a, 16'h071b, 16'h071c, 16'h071d, 16'h071e, 16'h071f 	:	val_out <= 16'h962c;
         16'h0720, 16'h0721, 16'h0722, 16'h0723, 16'h0724, 16'h0725, 16'h0726, 16'h0727 	:	val_out <= 16'h9645;
         16'h0728, 16'h0729, 16'h072a, 16'h072b, 16'h072c, 16'h072d, 16'h072e, 16'h072f 	:	val_out <= 16'h965d;
         16'h0730, 16'h0731, 16'h0732, 16'h0733, 16'h0734, 16'h0735, 16'h0736, 16'h0737 	:	val_out <= 16'h9676;
         16'h0738, 16'h0739, 16'h073a, 16'h073b, 16'h073c, 16'h073d, 16'h073e, 16'h073f 	:	val_out <= 16'h968f;
         16'h0740, 16'h0741, 16'h0742, 16'h0743, 16'h0744, 16'h0745, 16'h0746, 16'h0747 	:	val_out <= 16'h96a8;
         16'h0748, 16'h0749, 16'h074a, 16'h074b, 16'h074c, 16'h074d, 16'h074e, 16'h074f 	:	val_out <= 16'h96c0;
         16'h0750, 16'h0751, 16'h0752, 16'h0753, 16'h0754, 16'h0755, 16'h0756, 16'h0757 	:	val_out <= 16'h96d9;
         16'h0758, 16'h0759, 16'h075a, 16'h075b, 16'h075c, 16'h075d, 16'h075e, 16'h075f 	:	val_out <= 16'h96f2;
         16'h0760, 16'h0761, 16'h0762, 16'h0763, 16'h0764, 16'h0765, 16'h0766, 16'h0767 	:	val_out <= 16'h970a;
         16'h0768, 16'h0769, 16'h076a, 16'h076b, 16'h076c, 16'h076d, 16'h076e, 16'h076f 	:	val_out <= 16'h9723;
         16'h0770, 16'h0771, 16'h0772, 16'h0773, 16'h0774, 16'h0775, 16'h0776, 16'h0777 	:	val_out <= 16'h973c;
         16'h0778, 16'h0779, 16'h077a, 16'h077b, 16'h077c, 16'h077d, 16'h077e, 16'h077f 	:	val_out <= 16'h9755;
         16'h0780, 16'h0781, 16'h0782, 16'h0783, 16'h0784, 16'h0785, 16'h0786, 16'h0787 	:	val_out <= 16'h976d;
         16'h0788, 16'h0789, 16'h078a, 16'h078b, 16'h078c, 16'h078d, 16'h078e, 16'h078f 	:	val_out <= 16'h9786;
         16'h0790, 16'h0791, 16'h0792, 16'h0793, 16'h0794, 16'h0795, 16'h0796, 16'h0797 	:	val_out <= 16'h979f;
         16'h0798, 16'h0799, 16'h079a, 16'h079b, 16'h079c, 16'h079d, 16'h079e, 16'h079f 	:	val_out <= 16'h97b7;
         16'h07a0, 16'h07a1, 16'h07a2, 16'h07a3, 16'h07a4, 16'h07a5, 16'h07a6, 16'h07a7 	:	val_out <= 16'h97d0;
         16'h07a8, 16'h07a9, 16'h07aa, 16'h07ab, 16'h07ac, 16'h07ad, 16'h07ae, 16'h07af 	:	val_out <= 16'h97e9;
         16'h07b0, 16'h07b1, 16'h07b2, 16'h07b3, 16'h07b4, 16'h07b5, 16'h07b6, 16'h07b7 	:	val_out <= 16'h9802;
         16'h07b8, 16'h07b9, 16'h07ba, 16'h07bb, 16'h07bc, 16'h07bd, 16'h07be, 16'h07bf 	:	val_out <= 16'h981a;
         16'h07c0, 16'h07c1, 16'h07c2, 16'h07c3, 16'h07c4, 16'h07c5, 16'h07c6, 16'h07c7 	:	val_out <= 16'h9833;
         16'h07c8, 16'h07c9, 16'h07ca, 16'h07cb, 16'h07cc, 16'h07cd, 16'h07ce, 16'h07cf 	:	val_out <= 16'h984c;
         16'h07d0, 16'h07d1, 16'h07d2, 16'h07d3, 16'h07d4, 16'h07d5, 16'h07d6, 16'h07d7 	:	val_out <= 16'h9864;
         16'h07d8, 16'h07d9, 16'h07da, 16'h07db, 16'h07dc, 16'h07dd, 16'h07de, 16'h07df 	:	val_out <= 16'h987d;
         16'h07e0, 16'h07e1, 16'h07e2, 16'h07e3, 16'h07e4, 16'h07e5, 16'h07e6, 16'h07e7 	:	val_out <= 16'h9896;
         16'h07e8, 16'h07e9, 16'h07ea, 16'h07eb, 16'h07ec, 16'h07ed, 16'h07ee, 16'h07ef 	:	val_out <= 16'h98ae;
         16'h07f0, 16'h07f1, 16'h07f2, 16'h07f3, 16'h07f4, 16'h07f5, 16'h07f6, 16'h07f7 	:	val_out <= 16'h98c7;
         16'h07f8, 16'h07f9, 16'h07fa, 16'h07fb, 16'h07fc, 16'h07fd, 16'h07fe, 16'h07ff 	:	val_out <= 16'h98e0;
         16'h0800, 16'h0801, 16'h0802, 16'h0803, 16'h0804, 16'h0805, 16'h0806, 16'h0807 	:	val_out <= 16'h98f8;
         16'h0808, 16'h0809, 16'h080a, 16'h080b, 16'h080c, 16'h080d, 16'h080e, 16'h080f 	:	val_out <= 16'h9911;
         16'h0810, 16'h0811, 16'h0812, 16'h0813, 16'h0814, 16'h0815, 16'h0816, 16'h0817 	:	val_out <= 16'h992a;
         16'h0818, 16'h0819, 16'h081a, 16'h081b, 16'h081c, 16'h081d, 16'h081e, 16'h081f 	:	val_out <= 16'h9942;
         16'h0820, 16'h0821, 16'h0822, 16'h0823, 16'h0824, 16'h0825, 16'h0826, 16'h0827 	:	val_out <= 16'h995b;
         16'h0828, 16'h0829, 16'h082a, 16'h082b, 16'h082c, 16'h082d, 16'h082e, 16'h082f 	:	val_out <= 16'h9973;
         16'h0830, 16'h0831, 16'h0832, 16'h0833, 16'h0834, 16'h0835, 16'h0836, 16'h0837 	:	val_out <= 16'h998c;
         16'h0838, 16'h0839, 16'h083a, 16'h083b, 16'h083c, 16'h083d, 16'h083e, 16'h083f 	:	val_out <= 16'h99a5;
         16'h0840, 16'h0841, 16'h0842, 16'h0843, 16'h0844, 16'h0845, 16'h0846, 16'h0847 	:	val_out <= 16'h99bd;
         16'h0848, 16'h0849, 16'h084a, 16'h084b, 16'h084c, 16'h084d, 16'h084e, 16'h084f 	:	val_out <= 16'h99d6;
         16'h0850, 16'h0851, 16'h0852, 16'h0853, 16'h0854, 16'h0855, 16'h0856, 16'h0857 	:	val_out <= 16'h99ef;
         16'h0858, 16'h0859, 16'h085a, 16'h085b, 16'h085c, 16'h085d, 16'h085e, 16'h085f 	:	val_out <= 16'h9a07;
         16'h0860, 16'h0861, 16'h0862, 16'h0863, 16'h0864, 16'h0865, 16'h0866, 16'h0867 	:	val_out <= 16'h9a20;
         16'h0868, 16'h0869, 16'h086a, 16'h086b, 16'h086c, 16'h086d, 16'h086e, 16'h086f 	:	val_out <= 16'h9a38;
         16'h0870, 16'h0871, 16'h0872, 16'h0873, 16'h0874, 16'h0875, 16'h0876, 16'h0877 	:	val_out <= 16'h9a51;
         16'h0878, 16'h0879, 16'h087a, 16'h087b, 16'h087c, 16'h087d, 16'h087e, 16'h087f 	:	val_out <= 16'h9a6a;
         16'h0880, 16'h0881, 16'h0882, 16'h0883, 16'h0884, 16'h0885, 16'h0886, 16'h0887 	:	val_out <= 16'h9a82;
         16'h0888, 16'h0889, 16'h088a, 16'h088b, 16'h088c, 16'h088d, 16'h088e, 16'h088f 	:	val_out <= 16'h9a9b;
         16'h0890, 16'h0891, 16'h0892, 16'h0893, 16'h0894, 16'h0895, 16'h0896, 16'h0897 	:	val_out <= 16'h9ab3;
         16'h0898, 16'h0899, 16'h089a, 16'h089b, 16'h089c, 16'h089d, 16'h089e, 16'h089f 	:	val_out <= 16'h9acc;
         16'h08a0, 16'h08a1, 16'h08a2, 16'h08a3, 16'h08a4, 16'h08a5, 16'h08a6, 16'h08a7 	:	val_out <= 16'h9ae4;
         16'h08a8, 16'h08a9, 16'h08aa, 16'h08ab, 16'h08ac, 16'h08ad, 16'h08ae, 16'h08af 	:	val_out <= 16'h9afd;
         16'h08b0, 16'h08b1, 16'h08b2, 16'h08b3, 16'h08b4, 16'h08b5, 16'h08b6, 16'h08b7 	:	val_out <= 16'h9b16;
         16'h08b8, 16'h08b9, 16'h08ba, 16'h08bb, 16'h08bc, 16'h08bd, 16'h08be, 16'h08bf 	:	val_out <= 16'h9b2e;
         16'h08c0, 16'h08c1, 16'h08c2, 16'h08c3, 16'h08c4, 16'h08c5, 16'h08c6, 16'h08c7 	:	val_out <= 16'h9b47;
         16'h08c8, 16'h08c9, 16'h08ca, 16'h08cb, 16'h08cc, 16'h08cd, 16'h08ce, 16'h08cf 	:	val_out <= 16'h9b5f;
         16'h08d0, 16'h08d1, 16'h08d2, 16'h08d3, 16'h08d4, 16'h08d5, 16'h08d6, 16'h08d7 	:	val_out <= 16'h9b78;
         16'h08d8, 16'h08d9, 16'h08da, 16'h08db, 16'h08dc, 16'h08dd, 16'h08de, 16'h08df 	:	val_out <= 16'h9b90;
         16'h08e0, 16'h08e1, 16'h08e2, 16'h08e3, 16'h08e4, 16'h08e5, 16'h08e6, 16'h08e7 	:	val_out <= 16'h9ba9;
         16'h08e8, 16'h08e9, 16'h08ea, 16'h08eb, 16'h08ec, 16'h08ed, 16'h08ee, 16'h08ef 	:	val_out <= 16'h9bc1;
         16'h08f0, 16'h08f1, 16'h08f2, 16'h08f3, 16'h08f4, 16'h08f5, 16'h08f6, 16'h08f7 	:	val_out <= 16'h9bda;
         16'h08f8, 16'h08f9, 16'h08fa, 16'h08fb, 16'h08fc, 16'h08fd, 16'h08fe, 16'h08ff 	:	val_out <= 16'h9bf2;
         16'h0900, 16'h0901, 16'h0902, 16'h0903, 16'h0904, 16'h0905, 16'h0906, 16'h0907 	:	val_out <= 16'h9c0b;
         16'h0908, 16'h0909, 16'h090a, 16'h090b, 16'h090c, 16'h090d, 16'h090e, 16'h090f 	:	val_out <= 16'h9c24;
         16'h0910, 16'h0911, 16'h0912, 16'h0913, 16'h0914, 16'h0915, 16'h0916, 16'h0917 	:	val_out <= 16'h9c3c;
         16'h0918, 16'h0919, 16'h091a, 16'h091b, 16'h091c, 16'h091d, 16'h091e, 16'h091f 	:	val_out <= 16'h9c55;
         16'h0920, 16'h0921, 16'h0922, 16'h0923, 16'h0924, 16'h0925, 16'h0926, 16'h0927 	:	val_out <= 16'h9c6d;
         16'h0928, 16'h0929, 16'h092a, 16'h092b, 16'h092c, 16'h092d, 16'h092e, 16'h092f 	:	val_out <= 16'h9c86;
         16'h0930, 16'h0931, 16'h0932, 16'h0933, 16'h0934, 16'h0935, 16'h0936, 16'h0937 	:	val_out <= 16'h9c9e;
         16'h0938, 16'h0939, 16'h093a, 16'h093b, 16'h093c, 16'h093d, 16'h093e, 16'h093f 	:	val_out <= 16'h9cb7;
         16'h0940, 16'h0941, 16'h0942, 16'h0943, 16'h0944, 16'h0945, 16'h0946, 16'h0947 	:	val_out <= 16'h9ccf;
         16'h0948, 16'h0949, 16'h094a, 16'h094b, 16'h094c, 16'h094d, 16'h094e, 16'h094f 	:	val_out <= 16'h9ce8;
         16'h0950, 16'h0951, 16'h0952, 16'h0953, 16'h0954, 16'h0955, 16'h0956, 16'h0957 	:	val_out <= 16'h9d00;
         16'h0958, 16'h0959, 16'h095a, 16'h095b, 16'h095c, 16'h095d, 16'h095e, 16'h095f 	:	val_out <= 16'h9d18;
         16'h0960, 16'h0961, 16'h0962, 16'h0963, 16'h0964, 16'h0965, 16'h0966, 16'h0967 	:	val_out <= 16'h9d31;
         16'h0968, 16'h0969, 16'h096a, 16'h096b, 16'h096c, 16'h096d, 16'h096e, 16'h096f 	:	val_out <= 16'h9d49;
         16'h0970, 16'h0971, 16'h0972, 16'h0973, 16'h0974, 16'h0975, 16'h0976, 16'h0977 	:	val_out <= 16'h9d62;
         16'h0978, 16'h0979, 16'h097a, 16'h097b, 16'h097c, 16'h097d, 16'h097e, 16'h097f 	:	val_out <= 16'h9d7a;
         16'h0980, 16'h0981, 16'h0982, 16'h0983, 16'h0984, 16'h0985, 16'h0986, 16'h0987 	:	val_out <= 16'h9d93;
         16'h0988, 16'h0989, 16'h098a, 16'h098b, 16'h098c, 16'h098d, 16'h098e, 16'h098f 	:	val_out <= 16'h9dab;
         16'h0990, 16'h0991, 16'h0992, 16'h0993, 16'h0994, 16'h0995, 16'h0996, 16'h0997 	:	val_out <= 16'h9dc4;
         16'h0998, 16'h0999, 16'h099a, 16'h099b, 16'h099c, 16'h099d, 16'h099e, 16'h099f 	:	val_out <= 16'h9ddc;
         16'h09a0, 16'h09a1, 16'h09a2, 16'h09a3, 16'h09a4, 16'h09a5, 16'h09a6, 16'h09a7 	:	val_out <= 16'h9df5;
         16'h09a8, 16'h09a9, 16'h09aa, 16'h09ab, 16'h09ac, 16'h09ad, 16'h09ae, 16'h09af 	:	val_out <= 16'h9e0d;
         16'h09b0, 16'h09b1, 16'h09b2, 16'h09b3, 16'h09b4, 16'h09b5, 16'h09b6, 16'h09b7 	:	val_out <= 16'h9e25;
         16'h09b8, 16'h09b9, 16'h09ba, 16'h09bb, 16'h09bc, 16'h09bd, 16'h09be, 16'h09bf 	:	val_out <= 16'h9e3e;
         16'h09c0, 16'h09c1, 16'h09c2, 16'h09c3, 16'h09c4, 16'h09c5, 16'h09c6, 16'h09c7 	:	val_out <= 16'h9e56;
         16'h09c8, 16'h09c9, 16'h09ca, 16'h09cb, 16'h09cc, 16'h09cd, 16'h09ce, 16'h09cf 	:	val_out <= 16'h9e6f;
         16'h09d0, 16'h09d1, 16'h09d2, 16'h09d3, 16'h09d4, 16'h09d5, 16'h09d6, 16'h09d7 	:	val_out <= 16'h9e87;
         16'h09d8, 16'h09d9, 16'h09da, 16'h09db, 16'h09dc, 16'h09dd, 16'h09de, 16'h09df 	:	val_out <= 16'h9ea0;
         16'h09e0, 16'h09e1, 16'h09e2, 16'h09e3, 16'h09e4, 16'h09e5, 16'h09e6, 16'h09e7 	:	val_out <= 16'h9eb8;
         16'h09e8, 16'h09e9, 16'h09ea, 16'h09eb, 16'h09ec, 16'h09ed, 16'h09ee, 16'h09ef 	:	val_out <= 16'h9ed0;
         16'h09f0, 16'h09f1, 16'h09f2, 16'h09f3, 16'h09f4, 16'h09f5, 16'h09f6, 16'h09f7 	:	val_out <= 16'h9ee9;
         16'h09f8, 16'h09f9, 16'h09fa, 16'h09fb, 16'h09fc, 16'h09fd, 16'h09fe, 16'h09ff 	:	val_out <= 16'h9f01;
         16'h0a00, 16'h0a01, 16'h0a02, 16'h0a03, 16'h0a04, 16'h0a05, 16'h0a06, 16'h0a07 	:	val_out <= 16'h9f19;
         16'h0a08, 16'h0a09, 16'h0a0a, 16'h0a0b, 16'h0a0c, 16'h0a0d, 16'h0a0e, 16'h0a0f 	:	val_out <= 16'h9f32;
         16'h0a10, 16'h0a11, 16'h0a12, 16'h0a13, 16'h0a14, 16'h0a15, 16'h0a16, 16'h0a17 	:	val_out <= 16'h9f4a;
         16'h0a18, 16'h0a19, 16'h0a1a, 16'h0a1b, 16'h0a1c, 16'h0a1d, 16'h0a1e, 16'h0a1f 	:	val_out <= 16'h9f63;
         16'h0a20, 16'h0a21, 16'h0a22, 16'h0a23, 16'h0a24, 16'h0a25, 16'h0a26, 16'h0a27 	:	val_out <= 16'h9f7b;
         16'h0a28, 16'h0a29, 16'h0a2a, 16'h0a2b, 16'h0a2c, 16'h0a2d, 16'h0a2e, 16'h0a2f 	:	val_out <= 16'h9f93;
         16'h0a30, 16'h0a31, 16'h0a32, 16'h0a33, 16'h0a34, 16'h0a35, 16'h0a36, 16'h0a37 	:	val_out <= 16'h9fac;
         16'h0a38, 16'h0a39, 16'h0a3a, 16'h0a3b, 16'h0a3c, 16'h0a3d, 16'h0a3e, 16'h0a3f 	:	val_out <= 16'h9fc4;
         16'h0a40, 16'h0a41, 16'h0a42, 16'h0a43, 16'h0a44, 16'h0a45, 16'h0a46, 16'h0a47 	:	val_out <= 16'h9fdc;
         16'h0a48, 16'h0a49, 16'h0a4a, 16'h0a4b, 16'h0a4c, 16'h0a4d, 16'h0a4e, 16'h0a4f 	:	val_out <= 16'h9ff5;
         16'h0a50, 16'h0a51, 16'h0a52, 16'h0a53, 16'h0a54, 16'h0a55, 16'h0a56, 16'h0a57 	:	val_out <= 16'ha00d;
         16'h0a58, 16'h0a59, 16'h0a5a, 16'h0a5b, 16'h0a5c, 16'h0a5d, 16'h0a5e, 16'h0a5f 	:	val_out <= 16'ha025;
         16'h0a60, 16'h0a61, 16'h0a62, 16'h0a63, 16'h0a64, 16'h0a65, 16'h0a66, 16'h0a67 	:	val_out <= 16'ha03e;
         16'h0a68, 16'h0a69, 16'h0a6a, 16'h0a6b, 16'h0a6c, 16'h0a6d, 16'h0a6e, 16'h0a6f 	:	val_out <= 16'ha056;
         16'h0a70, 16'h0a71, 16'h0a72, 16'h0a73, 16'h0a74, 16'h0a75, 16'h0a76, 16'h0a77 	:	val_out <= 16'ha06e;
         16'h0a78, 16'h0a79, 16'h0a7a, 16'h0a7b, 16'h0a7c, 16'h0a7d, 16'h0a7e, 16'h0a7f 	:	val_out <= 16'ha087;
         16'h0a80, 16'h0a81, 16'h0a82, 16'h0a83, 16'h0a84, 16'h0a85, 16'h0a86, 16'h0a87 	:	val_out <= 16'ha09f;
         16'h0a88, 16'h0a89, 16'h0a8a, 16'h0a8b, 16'h0a8c, 16'h0a8d, 16'h0a8e, 16'h0a8f 	:	val_out <= 16'ha0b7;
         16'h0a90, 16'h0a91, 16'h0a92, 16'h0a93, 16'h0a94, 16'h0a95, 16'h0a96, 16'h0a97 	:	val_out <= 16'ha0d0;
         16'h0a98, 16'h0a99, 16'h0a9a, 16'h0a9b, 16'h0a9c, 16'h0a9d, 16'h0a9e, 16'h0a9f 	:	val_out <= 16'ha0e8;
         16'h0aa0, 16'h0aa1, 16'h0aa2, 16'h0aa3, 16'h0aa4, 16'h0aa5, 16'h0aa6, 16'h0aa7 	:	val_out <= 16'ha100;
         16'h0aa8, 16'h0aa9, 16'h0aaa, 16'h0aab, 16'h0aac, 16'h0aad, 16'h0aae, 16'h0aaf 	:	val_out <= 16'ha118;
         16'h0ab0, 16'h0ab1, 16'h0ab2, 16'h0ab3, 16'h0ab4, 16'h0ab5, 16'h0ab6, 16'h0ab7 	:	val_out <= 16'ha131;
         16'h0ab8, 16'h0ab9, 16'h0aba, 16'h0abb, 16'h0abc, 16'h0abd, 16'h0abe, 16'h0abf 	:	val_out <= 16'ha149;
         16'h0ac0, 16'h0ac1, 16'h0ac2, 16'h0ac3, 16'h0ac4, 16'h0ac5, 16'h0ac6, 16'h0ac7 	:	val_out <= 16'ha161;
         16'h0ac8, 16'h0ac9, 16'h0aca, 16'h0acb, 16'h0acc, 16'h0acd, 16'h0ace, 16'h0acf 	:	val_out <= 16'ha179;
         16'h0ad0, 16'h0ad1, 16'h0ad2, 16'h0ad3, 16'h0ad4, 16'h0ad5, 16'h0ad6, 16'h0ad7 	:	val_out <= 16'ha192;
         16'h0ad8, 16'h0ad9, 16'h0ada, 16'h0adb, 16'h0adc, 16'h0add, 16'h0ade, 16'h0adf 	:	val_out <= 16'ha1aa;
         16'h0ae0, 16'h0ae1, 16'h0ae2, 16'h0ae3, 16'h0ae4, 16'h0ae5, 16'h0ae6, 16'h0ae7 	:	val_out <= 16'ha1c2;
         16'h0ae8, 16'h0ae9, 16'h0aea, 16'h0aeb, 16'h0aec, 16'h0aed, 16'h0aee, 16'h0aef 	:	val_out <= 16'ha1da;
         16'h0af0, 16'h0af1, 16'h0af2, 16'h0af3, 16'h0af4, 16'h0af5, 16'h0af6, 16'h0af7 	:	val_out <= 16'ha1f3;
         16'h0af8, 16'h0af9, 16'h0afa, 16'h0afb, 16'h0afc, 16'h0afd, 16'h0afe, 16'h0aff 	:	val_out <= 16'ha20b;
         16'h0b00, 16'h0b01, 16'h0b02, 16'h0b03, 16'h0b04, 16'h0b05, 16'h0b06, 16'h0b07 	:	val_out <= 16'ha223;
         16'h0b08, 16'h0b09, 16'h0b0a, 16'h0b0b, 16'h0b0c, 16'h0b0d, 16'h0b0e, 16'h0b0f 	:	val_out <= 16'ha23b;
         16'h0b10, 16'h0b11, 16'h0b12, 16'h0b13, 16'h0b14, 16'h0b15, 16'h0b16, 16'h0b17 	:	val_out <= 16'ha254;
         16'h0b18, 16'h0b19, 16'h0b1a, 16'h0b1b, 16'h0b1c, 16'h0b1d, 16'h0b1e, 16'h0b1f 	:	val_out <= 16'ha26c;
         16'h0b20, 16'h0b21, 16'h0b22, 16'h0b23, 16'h0b24, 16'h0b25, 16'h0b26, 16'h0b27 	:	val_out <= 16'ha284;
         16'h0b28, 16'h0b29, 16'h0b2a, 16'h0b2b, 16'h0b2c, 16'h0b2d, 16'h0b2e, 16'h0b2f 	:	val_out <= 16'ha29c;
         16'h0b30, 16'h0b31, 16'h0b32, 16'h0b33, 16'h0b34, 16'h0b35, 16'h0b36, 16'h0b37 	:	val_out <= 16'ha2b4;
         16'h0b38, 16'h0b39, 16'h0b3a, 16'h0b3b, 16'h0b3c, 16'h0b3d, 16'h0b3e, 16'h0b3f 	:	val_out <= 16'ha2cd;
         16'h0b40, 16'h0b41, 16'h0b42, 16'h0b43, 16'h0b44, 16'h0b45, 16'h0b46, 16'h0b47 	:	val_out <= 16'ha2e5;
         16'h0b48, 16'h0b49, 16'h0b4a, 16'h0b4b, 16'h0b4c, 16'h0b4d, 16'h0b4e, 16'h0b4f 	:	val_out <= 16'ha2fd;
         16'h0b50, 16'h0b51, 16'h0b52, 16'h0b53, 16'h0b54, 16'h0b55, 16'h0b56, 16'h0b57 	:	val_out <= 16'ha315;
         16'h0b58, 16'h0b59, 16'h0b5a, 16'h0b5b, 16'h0b5c, 16'h0b5d, 16'h0b5e, 16'h0b5f 	:	val_out <= 16'ha32d;
         16'h0b60, 16'h0b61, 16'h0b62, 16'h0b63, 16'h0b64, 16'h0b65, 16'h0b66, 16'h0b67 	:	val_out <= 16'ha345;
         16'h0b68, 16'h0b69, 16'h0b6a, 16'h0b6b, 16'h0b6c, 16'h0b6d, 16'h0b6e, 16'h0b6f 	:	val_out <= 16'ha35e;
         16'h0b70, 16'h0b71, 16'h0b72, 16'h0b73, 16'h0b74, 16'h0b75, 16'h0b76, 16'h0b77 	:	val_out <= 16'ha376;
         16'h0b78, 16'h0b79, 16'h0b7a, 16'h0b7b, 16'h0b7c, 16'h0b7d, 16'h0b7e, 16'h0b7f 	:	val_out <= 16'ha38e;
         16'h0b80, 16'h0b81, 16'h0b82, 16'h0b83, 16'h0b84, 16'h0b85, 16'h0b86, 16'h0b87 	:	val_out <= 16'ha3a6;
         16'h0b88, 16'h0b89, 16'h0b8a, 16'h0b8b, 16'h0b8c, 16'h0b8d, 16'h0b8e, 16'h0b8f 	:	val_out <= 16'ha3be;
         16'h0b90, 16'h0b91, 16'h0b92, 16'h0b93, 16'h0b94, 16'h0b95, 16'h0b96, 16'h0b97 	:	val_out <= 16'ha3d6;
         16'h0b98, 16'h0b99, 16'h0b9a, 16'h0b9b, 16'h0b9c, 16'h0b9d, 16'h0b9e, 16'h0b9f 	:	val_out <= 16'ha3ee;
         16'h0ba0, 16'h0ba1, 16'h0ba2, 16'h0ba3, 16'h0ba4, 16'h0ba5, 16'h0ba6, 16'h0ba7 	:	val_out <= 16'ha407;
         16'h0ba8, 16'h0ba9, 16'h0baa, 16'h0bab, 16'h0bac, 16'h0bad, 16'h0bae, 16'h0baf 	:	val_out <= 16'ha41f;
         16'h0bb0, 16'h0bb1, 16'h0bb2, 16'h0bb3, 16'h0bb4, 16'h0bb5, 16'h0bb6, 16'h0bb7 	:	val_out <= 16'ha437;
         16'h0bb8, 16'h0bb9, 16'h0bba, 16'h0bbb, 16'h0bbc, 16'h0bbd, 16'h0bbe, 16'h0bbf 	:	val_out <= 16'ha44f;
         16'h0bc0, 16'h0bc1, 16'h0bc2, 16'h0bc3, 16'h0bc4, 16'h0bc5, 16'h0bc6, 16'h0bc7 	:	val_out <= 16'ha467;
         16'h0bc8, 16'h0bc9, 16'h0bca, 16'h0bcb, 16'h0bcc, 16'h0bcd, 16'h0bce, 16'h0bcf 	:	val_out <= 16'ha47f;
         16'h0bd0, 16'h0bd1, 16'h0bd2, 16'h0bd3, 16'h0bd4, 16'h0bd5, 16'h0bd6, 16'h0bd7 	:	val_out <= 16'ha497;
         16'h0bd8, 16'h0bd9, 16'h0bda, 16'h0bdb, 16'h0bdc, 16'h0bdd, 16'h0bde, 16'h0bdf 	:	val_out <= 16'ha4af;
         16'h0be0, 16'h0be1, 16'h0be2, 16'h0be3, 16'h0be4, 16'h0be5, 16'h0be6, 16'h0be7 	:	val_out <= 16'ha4c7;
         16'h0be8, 16'h0be9, 16'h0bea, 16'h0beb, 16'h0bec, 16'h0bed, 16'h0bee, 16'h0bef 	:	val_out <= 16'ha4df;
         16'h0bf0, 16'h0bf1, 16'h0bf2, 16'h0bf3, 16'h0bf4, 16'h0bf5, 16'h0bf6, 16'h0bf7 	:	val_out <= 16'ha4f7;
         16'h0bf8, 16'h0bf9, 16'h0bfa, 16'h0bfb, 16'h0bfc, 16'h0bfd, 16'h0bfe, 16'h0bff 	:	val_out <= 16'ha50f;
         16'h0c00, 16'h0c01, 16'h0c02, 16'h0c03, 16'h0c04, 16'h0c05, 16'h0c06, 16'h0c07 	:	val_out <= 16'ha528;
         16'h0c08, 16'h0c09, 16'h0c0a, 16'h0c0b, 16'h0c0c, 16'h0c0d, 16'h0c0e, 16'h0c0f 	:	val_out <= 16'ha540;
         16'h0c10, 16'h0c11, 16'h0c12, 16'h0c13, 16'h0c14, 16'h0c15, 16'h0c16, 16'h0c17 	:	val_out <= 16'ha558;
         16'h0c18, 16'h0c19, 16'h0c1a, 16'h0c1b, 16'h0c1c, 16'h0c1d, 16'h0c1e, 16'h0c1f 	:	val_out <= 16'ha570;
         16'h0c20, 16'h0c21, 16'h0c22, 16'h0c23, 16'h0c24, 16'h0c25, 16'h0c26, 16'h0c27 	:	val_out <= 16'ha588;
         16'h0c28, 16'h0c29, 16'h0c2a, 16'h0c2b, 16'h0c2c, 16'h0c2d, 16'h0c2e, 16'h0c2f 	:	val_out <= 16'ha5a0;
         16'h0c30, 16'h0c31, 16'h0c32, 16'h0c33, 16'h0c34, 16'h0c35, 16'h0c36, 16'h0c37 	:	val_out <= 16'ha5b8;
         16'h0c38, 16'h0c39, 16'h0c3a, 16'h0c3b, 16'h0c3c, 16'h0c3d, 16'h0c3e, 16'h0c3f 	:	val_out <= 16'ha5d0;
         16'h0c40, 16'h0c41, 16'h0c42, 16'h0c43, 16'h0c44, 16'h0c45, 16'h0c46, 16'h0c47 	:	val_out <= 16'ha5e8;
         16'h0c48, 16'h0c49, 16'h0c4a, 16'h0c4b, 16'h0c4c, 16'h0c4d, 16'h0c4e, 16'h0c4f 	:	val_out <= 16'ha600;
         16'h0c50, 16'h0c51, 16'h0c52, 16'h0c53, 16'h0c54, 16'h0c55, 16'h0c56, 16'h0c57 	:	val_out <= 16'ha618;
         16'h0c58, 16'h0c59, 16'h0c5a, 16'h0c5b, 16'h0c5c, 16'h0c5d, 16'h0c5e, 16'h0c5f 	:	val_out <= 16'ha630;
         16'h0c60, 16'h0c61, 16'h0c62, 16'h0c63, 16'h0c64, 16'h0c65, 16'h0c66, 16'h0c67 	:	val_out <= 16'ha648;
         16'h0c68, 16'h0c69, 16'h0c6a, 16'h0c6b, 16'h0c6c, 16'h0c6d, 16'h0c6e, 16'h0c6f 	:	val_out <= 16'ha660;
         16'h0c70, 16'h0c71, 16'h0c72, 16'h0c73, 16'h0c74, 16'h0c75, 16'h0c76, 16'h0c77 	:	val_out <= 16'ha678;
         16'h0c78, 16'h0c79, 16'h0c7a, 16'h0c7b, 16'h0c7c, 16'h0c7d, 16'h0c7e, 16'h0c7f 	:	val_out <= 16'ha690;
         16'h0c80, 16'h0c81, 16'h0c82, 16'h0c83, 16'h0c84, 16'h0c85, 16'h0c86, 16'h0c87 	:	val_out <= 16'ha6a8;
         16'h0c88, 16'h0c89, 16'h0c8a, 16'h0c8b, 16'h0c8c, 16'h0c8d, 16'h0c8e, 16'h0c8f 	:	val_out <= 16'ha6c0;
         16'h0c90, 16'h0c91, 16'h0c92, 16'h0c93, 16'h0c94, 16'h0c95, 16'h0c96, 16'h0c97 	:	val_out <= 16'ha6d8;
         16'h0c98, 16'h0c99, 16'h0c9a, 16'h0c9b, 16'h0c9c, 16'h0c9d, 16'h0c9e, 16'h0c9f 	:	val_out <= 16'ha6ef;
         16'h0ca0, 16'h0ca1, 16'h0ca2, 16'h0ca3, 16'h0ca4, 16'h0ca5, 16'h0ca6, 16'h0ca7 	:	val_out <= 16'ha707;
         16'h0ca8, 16'h0ca9, 16'h0caa, 16'h0cab, 16'h0cac, 16'h0cad, 16'h0cae, 16'h0caf 	:	val_out <= 16'ha71f;
         16'h0cb0, 16'h0cb1, 16'h0cb2, 16'h0cb3, 16'h0cb4, 16'h0cb5, 16'h0cb6, 16'h0cb7 	:	val_out <= 16'ha737;
         16'h0cb8, 16'h0cb9, 16'h0cba, 16'h0cbb, 16'h0cbc, 16'h0cbd, 16'h0cbe, 16'h0cbf 	:	val_out <= 16'ha74f;
         16'h0cc0, 16'h0cc1, 16'h0cc2, 16'h0cc3, 16'h0cc4, 16'h0cc5, 16'h0cc6, 16'h0cc7 	:	val_out <= 16'ha767;
         16'h0cc8, 16'h0cc9, 16'h0cca, 16'h0ccb, 16'h0ccc, 16'h0ccd, 16'h0cce, 16'h0ccf 	:	val_out <= 16'ha77f;
         16'h0cd0, 16'h0cd1, 16'h0cd2, 16'h0cd3, 16'h0cd4, 16'h0cd5, 16'h0cd6, 16'h0cd7 	:	val_out <= 16'ha797;
         16'h0cd8, 16'h0cd9, 16'h0cda, 16'h0cdb, 16'h0cdc, 16'h0cdd, 16'h0cde, 16'h0cdf 	:	val_out <= 16'ha7af;
         16'h0ce0, 16'h0ce1, 16'h0ce2, 16'h0ce3, 16'h0ce4, 16'h0ce5, 16'h0ce6, 16'h0ce7 	:	val_out <= 16'ha7c7;
         16'h0ce8, 16'h0ce9, 16'h0cea, 16'h0ceb, 16'h0cec, 16'h0ced, 16'h0cee, 16'h0cef 	:	val_out <= 16'ha7df;
         16'h0cf0, 16'h0cf1, 16'h0cf2, 16'h0cf3, 16'h0cf4, 16'h0cf5, 16'h0cf6, 16'h0cf7 	:	val_out <= 16'ha7f6;
         16'h0cf8, 16'h0cf9, 16'h0cfa, 16'h0cfb, 16'h0cfc, 16'h0cfd, 16'h0cfe, 16'h0cff 	:	val_out <= 16'ha80e;
         16'h0d00, 16'h0d01, 16'h0d02, 16'h0d03, 16'h0d04, 16'h0d05, 16'h0d06, 16'h0d07 	:	val_out <= 16'ha826;
         16'h0d08, 16'h0d09, 16'h0d0a, 16'h0d0b, 16'h0d0c, 16'h0d0d, 16'h0d0e, 16'h0d0f 	:	val_out <= 16'ha83e;
         16'h0d10, 16'h0d11, 16'h0d12, 16'h0d13, 16'h0d14, 16'h0d15, 16'h0d16, 16'h0d17 	:	val_out <= 16'ha856;
         16'h0d18, 16'h0d19, 16'h0d1a, 16'h0d1b, 16'h0d1c, 16'h0d1d, 16'h0d1e, 16'h0d1f 	:	val_out <= 16'ha86e;
         16'h0d20, 16'h0d21, 16'h0d22, 16'h0d23, 16'h0d24, 16'h0d25, 16'h0d26, 16'h0d27 	:	val_out <= 16'ha886;
         16'h0d28, 16'h0d29, 16'h0d2a, 16'h0d2b, 16'h0d2c, 16'h0d2d, 16'h0d2e, 16'h0d2f 	:	val_out <= 16'ha89d;
         16'h0d30, 16'h0d31, 16'h0d32, 16'h0d33, 16'h0d34, 16'h0d35, 16'h0d36, 16'h0d37 	:	val_out <= 16'ha8b5;
         16'h0d38, 16'h0d39, 16'h0d3a, 16'h0d3b, 16'h0d3c, 16'h0d3d, 16'h0d3e, 16'h0d3f 	:	val_out <= 16'ha8cd;
         16'h0d40, 16'h0d41, 16'h0d42, 16'h0d43, 16'h0d44, 16'h0d45, 16'h0d46, 16'h0d47 	:	val_out <= 16'ha8e5;
         16'h0d48, 16'h0d49, 16'h0d4a, 16'h0d4b, 16'h0d4c, 16'h0d4d, 16'h0d4e, 16'h0d4f 	:	val_out <= 16'ha8fd;
         16'h0d50, 16'h0d51, 16'h0d52, 16'h0d53, 16'h0d54, 16'h0d55, 16'h0d56, 16'h0d57 	:	val_out <= 16'ha915;
         16'h0d58, 16'h0d59, 16'h0d5a, 16'h0d5b, 16'h0d5c, 16'h0d5d, 16'h0d5e, 16'h0d5f 	:	val_out <= 16'ha92c;
         16'h0d60, 16'h0d61, 16'h0d62, 16'h0d63, 16'h0d64, 16'h0d65, 16'h0d66, 16'h0d67 	:	val_out <= 16'ha944;
         16'h0d68, 16'h0d69, 16'h0d6a, 16'h0d6b, 16'h0d6c, 16'h0d6d, 16'h0d6e, 16'h0d6f 	:	val_out <= 16'ha95c;
         16'h0d70, 16'h0d71, 16'h0d72, 16'h0d73, 16'h0d74, 16'h0d75, 16'h0d76, 16'h0d77 	:	val_out <= 16'ha974;
         16'h0d78, 16'h0d79, 16'h0d7a, 16'h0d7b, 16'h0d7c, 16'h0d7d, 16'h0d7e, 16'h0d7f 	:	val_out <= 16'ha98b;
         16'h0d80, 16'h0d81, 16'h0d82, 16'h0d83, 16'h0d84, 16'h0d85, 16'h0d86, 16'h0d87 	:	val_out <= 16'ha9a3;
         16'h0d88, 16'h0d89, 16'h0d8a, 16'h0d8b, 16'h0d8c, 16'h0d8d, 16'h0d8e, 16'h0d8f 	:	val_out <= 16'ha9bb;
         16'h0d90, 16'h0d91, 16'h0d92, 16'h0d93, 16'h0d94, 16'h0d95, 16'h0d96, 16'h0d97 	:	val_out <= 16'ha9d3;
         16'h0d98, 16'h0d99, 16'h0d9a, 16'h0d9b, 16'h0d9c, 16'h0d9d, 16'h0d9e, 16'h0d9f 	:	val_out <= 16'ha9eb;
         16'h0da0, 16'h0da1, 16'h0da2, 16'h0da3, 16'h0da4, 16'h0da5, 16'h0da6, 16'h0da7 	:	val_out <= 16'haa02;
         16'h0da8, 16'h0da9, 16'h0daa, 16'h0dab, 16'h0dac, 16'h0dad, 16'h0dae, 16'h0daf 	:	val_out <= 16'haa1a;
         16'h0db0, 16'h0db1, 16'h0db2, 16'h0db3, 16'h0db4, 16'h0db5, 16'h0db6, 16'h0db7 	:	val_out <= 16'haa32;
         16'h0db8, 16'h0db9, 16'h0dba, 16'h0dbb, 16'h0dbc, 16'h0dbd, 16'h0dbe, 16'h0dbf 	:	val_out <= 16'haa49;
         16'h0dc0, 16'h0dc1, 16'h0dc2, 16'h0dc3, 16'h0dc4, 16'h0dc5, 16'h0dc6, 16'h0dc7 	:	val_out <= 16'haa61;
         16'h0dc8, 16'h0dc9, 16'h0dca, 16'h0dcb, 16'h0dcc, 16'h0dcd, 16'h0dce, 16'h0dcf 	:	val_out <= 16'haa79;
         16'h0dd0, 16'h0dd1, 16'h0dd2, 16'h0dd3, 16'h0dd4, 16'h0dd5, 16'h0dd6, 16'h0dd7 	:	val_out <= 16'haa91;
         16'h0dd8, 16'h0dd9, 16'h0dda, 16'h0ddb, 16'h0ddc, 16'h0ddd, 16'h0dde, 16'h0ddf 	:	val_out <= 16'haaa8;
         16'h0de0, 16'h0de1, 16'h0de2, 16'h0de3, 16'h0de4, 16'h0de5, 16'h0de6, 16'h0de7 	:	val_out <= 16'haac0;
         16'h0de8, 16'h0de9, 16'h0dea, 16'h0deb, 16'h0dec, 16'h0ded, 16'h0dee, 16'h0def 	:	val_out <= 16'haad8;
         16'h0df0, 16'h0df1, 16'h0df2, 16'h0df3, 16'h0df4, 16'h0df5, 16'h0df6, 16'h0df7 	:	val_out <= 16'haaef;
         16'h0df8, 16'h0df9, 16'h0dfa, 16'h0dfb, 16'h0dfc, 16'h0dfd, 16'h0dfe, 16'h0dff 	:	val_out <= 16'hab07;
         16'h0e00, 16'h0e01, 16'h0e02, 16'h0e03, 16'h0e04, 16'h0e05, 16'h0e06, 16'h0e07 	:	val_out <= 16'hab1f;
         16'h0e08, 16'h0e09, 16'h0e0a, 16'h0e0b, 16'h0e0c, 16'h0e0d, 16'h0e0e, 16'h0e0f 	:	val_out <= 16'hab36;
         16'h0e10, 16'h0e11, 16'h0e12, 16'h0e13, 16'h0e14, 16'h0e15, 16'h0e16, 16'h0e17 	:	val_out <= 16'hab4e;
         16'h0e18, 16'h0e19, 16'h0e1a, 16'h0e1b, 16'h0e1c, 16'h0e1d, 16'h0e1e, 16'h0e1f 	:	val_out <= 16'hab66;
         16'h0e20, 16'h0e21, 16'h0e22, 16'h0e23, 16'h0e24, 16'h0e25, 16'h0e26, 16'h0e27 	:	val_out <= 16'hab7d;
         16'h0e28, 16'h0e29, 16'h0e2a, 16'h0e2b, 16'h0e2c, 16'h0e2d, 16'h0e2e, 16'h0e2f 	:	val_out <= 16'hab95;
         16'h0e30, 16'h0e31, 16'h0e32, 16'h0e33, 16'h0e34, 16'h0e35, 16'h0e36, 16'h0e37 	:	val_out <= 16'habad;
         16'h0e38, 16'h0e39, 16'h0e3a, 16'h0e3b, 16'h0e3c, 16'h0e3d, 16'h0e3e, 16'h0e3f 	:	val_out <= 16'habc4;
         16'h0e40, 16'h0e41, 16'h0e42, 16'h0e43, 16'h0e44, 16'h0e45, 16'h0e46, 16'h0e47 	:	val_out <= 16'habdc;
         16'h0e48, 16'h0e49, 16'h0e4a, 16'h0e4b, 16'h0e4c, 16'h0e4d, 16'h0e4e, 16'h0e4f 	:	val_out <= 16'habf3;
         16'h0e50, 16'h0e51, 16'h0e52, 16'h0e53, 16'h0e54, 16'h0e55, 16'h0e56, 16'h0e57 	:	val_out <= 16'hac0b;
         16'h0e58, 16'h0e59, 16'h0e5a, 16'h0e5b, 16'h0e5c, 16'h0e5d, 16'h0e5e, 16'h0e5f 	:	val_out <= 16'hac23;
         16'h0e60, 16'h0e61, 16'h0e62, 16'h0e63, 16'h0e64, 16'h0e65, 16'h0e66, 16'h0e67 	:	val_out <= 16'hac3a;
         16'h0e68, 16'h0e69, 16'h0e6a, 16'h0e6b, 16'h0e6c, 16'h0e6d, 16'h0e6e, 16'h0e6f 	:	val_out <= 16'hac52;
         16'h0e70, 16'h0e71, 16'h0e72, 16'h0e73, 16'h0e74, 16'h0e75, 16'h0e76, 16'h0e77 	:	val_out <= 16'hac69;
         16'h0e78, 16'h0e79, 16'h0e7a, 16'h0e7b, 16'h0e7c, 16'h0e7d, 16'h0e7e, 16'h0e7f 	:	val_out <= 16'hac81;
         16'h0e80, 16'h0e81, 16'h0e82, 16'h0e83, 16'h0e84, 16'h0e85, 16'h0e86, 16'h0e87 	:	val_out <= 16'hac98;
         16'h0e88, 16'h0e89, 16'h0e8a, 16'h0e8b, 16'h0e8c, 16'h0e8d, 16'h0e8e, 16'h0e8f 	:	val_out <= 16'hacb0;
         16'h0e90, 16'h0e91, 16'h0e92, 16'h0e93, 16'h0e94, 16'h0e95, 16'h0e96, 16'h0e97 	:	val_out <= 16'hacc8;
         16'h0e98, 16'h0e99, 16'h0e9a, 16'h0e9b, 16'h0e9c, 16'h0e9d, 16'h0e9e, 16'h0e9f 	:	val_out <= 16'hacdf;
         16'h0ea0, 16'h0ea1, 16'h0ea2, 16'h0ea3, 16'h0ea4, 16'h0ea5, 16'h0ea6, 16'h0ea7 	:	val_out <= 16'hacf7;
         16'h0ea8, 16'h0ea9, 16'h0eaa, 16'h0eab, 16'h0eac, 16'h0ead, 16'h0eae, 16'h0eaf 	:	val_out <= 16'had0e;
         16'h0eb0, 16'h0eb1, 16'h0eb2, 16'h0eb3, 16'h0eb4, 16'h0eb5, 16'h0eb6, 16'h0eb7 	:	val_out <= 16'had26;
         16'h0eb8, 16'h0eb9, 16'h0eba, 16'h0ebb, 16'h0ebc, 16'h0ebd, 16'h0ebe, 16'h0ebf 	:	val_out <= 16'had3d;
         16'h0ec0, 16'h0ec1, 16'h0ec2, 16'h0ec3, 16'h0ec4, 16'h0ec5, 16'h0ec6, 16'h0ec7 	:	val_out <= 16'had55;
         16'h0ec8, 16'h0ec9, 16'h0eca, 16'h0ecb, 16'h0ecc, 16'h0ecd, 16'h0ece, 16'h0ecf 	:	val_out <= 16'had6c;
         16'h0ed0, 16'h0ed1, 16'h0ed2, 16'h0ed3, 16'h0ed4, 16'h0ed5, 16'h0ed6, 16'h0ed7 	:	val_out <= 16'had84;
         16'h0ed8, 16'h0ed9, 16'h0eda, 16'h0edb, 16'h0edc, 16'h0edd, 16'h0ede, 16'h0edf 	:	val_out <= 16'had9b;
         16'h0ee0, 16'h0ee1, 16'h0ee2, 16'h0ee3, 16'h0ee4, 16'h0ee5, 16'h0ee6, 16'h0ee7 	:	val_out <= 16'hadb3;
         16'h0ee8, 16'h0ee9, 16'h0eea, 16'h0eeb, 16'h0eec, 16'h0eed, 16'h0eee, 16'h0eef 	:	val_out <= 16'hadca;
         16'h0ef0, 16'h0ef1, 16'h0ef2, 16'h0ef3, 16'h0ef4, 16'h0ef5, 16'h0ef6, 16'h0ef7 	:	val_out <= 16'hade2;
         16'h0ef8, 16'h0ef9, 16'h0efa, 16'h0efb, 16'h0efc, 16'h0efd, 16'h0efe, 16'h0eff 	:	val_out <= 16'hadf9;
         16'h0f00, 16'h0f01, 16'h0f02, 16'h0f03, 16'h0f04, 16'h0f05, 16'h0f06, 16'h0f07 	:	val_out <= 16'hae11;
         16'h0f08, 16'h0f09, 16'h0f0a, 16'h0f0b, 16'h0f0c, 16'h0f0d, 16'h0f0e, 16'h0f0f 	:	val_out <= 16'hae28;
         16'h0f10, 16'h0f11, 16'h0f12, 16'h0f13, 16'h0f14, 16'h0f15, 16'h0f16, 16'h0f17 	:	val_out <= 16'hae3f;
         16'h0f18, 16'h0f19, 16'h0f1a, 16'h0f1b, 16'h0f1c, 16'h0f1d, 16'h0f1e, 16'h0f1f 	:	val_out <= 16'hae57;
         16'h0f20, 16'h0f21, 16'h0f22, 16'h0f23, 16'h0f24, 16'h0f25, 16'h0f26, 16'h0f27 	:	val_out <= 16'hae6e;
         16'h0f28, 16'h0f29, 16'h0f2a, 16'h0f2b, 16'h0f2c, 16'h0f2d, 16'h0f2e, 16'h0f2f 	:	val_out <= 16'hae86;
         16'h0f30, 16'h0f31, 16'h0f32, 16'h0f33, 16'h0f34, 16'h0f35, 16'h0f36, 16'h0f37 	:	val_out <= 16'hae9d;
         16'h0f38, 16'h0f39, 16'h0f3a, 16'h0f3b, 16'h0f3c, 16'h0f3d, 16'h0f3e, 16'h0f3f 	:	val_out <= 16'haeb5;
         16'h0f40, 16'h0f41, 16'h0f42, 16'h0f43, 16'h0f44, 16'h0f45, 16'h0f46, 16'h0f47 	:	val_out <= 16'haecc;
         16'h0f48, 16'h0f49, 16'h0f4a, 16'h0f4b, 16'h0f4c, 16'h0f4d, 16'h0f4e, 16'h0f4f 	:	val_out <= 16'haee3;
         16'h0f50, 16'h0f51, 16'h0f52, 16'h0f53, 16'h0f54, 16'h0f55, 16'h0f56, 16'h0f57 	:	val_out <= 16'haefb;
         16'h0f58, 16'h0f59, 16'h0f5a, 16'h0f5b, 16'h0f5c, 16'h0f5d, 16'h0f5e, 16'h0f5f 	:	val_out <= 16'haf12;
         16'h0f60, 16'h0f61, 16'h0f62, 16'h0f63, 16'h0f64, 16'h0f65, 16'h0f66, 16'h0f67 	:	val_out <= 16'haf29;
         16'h0f68, 16'h0f69, 16'h0f6a, 16'h0f6b, 16'h0f6c, 16'h0f6d, 16'h0f6e, 16'h0f6f 	:	val_out <= 16'haf41;
         16'h0f70, 16'h0f71, 16'h0f72, 16'h0f73, 16'h0f74, 16'h0f75, 16'h0f76, 16'h0f77 	:	val_out <= 16'haf58;
         16'h0f78, 16'h0f79, 16'h0f7a, 16'h0f7b, 16'h0f7c, 16'h0f7d, 16'h0f7e, 16'h0f7f 	:	val_out <= 16'haf6f;
         16'h0f80, 16'h0f81, 16'h0f82, 16'h0f83, 16'h0f84, 16'h0f85, 16'h0f86, 16'h0f87 	:	val_out <= 16'haf87;
         16'h0f88, 16'h0f89, 16'h0f8a, 16'h0f8b, 16'h0f8c, 16'h0f8d, 16'h0f8e, 16'h0f8f 	:	val_out <= 16'haf9e;
         16'h0f90, 16'h0f91, 16'h0f92, 16'h0f93, 16'h0f94, 16'h0f95, 16'h0f96, 16'h0f97 	:	val_out <= 16'hafb5;
         16'h0f98, 16'h0f99, 16'h0f9a, 16'h0f9b, 16'h0f9c, 16'h0f9d, 16'h0f9e, 16'h0f9f 	:	val_out <= 16'hafcd;
         16'h0fa0, 16'h0fa1, 16'h0fa2, 16'h0fa3, 16'h0fa4, 16'h0fa5, 16'h0fa6, 16'h0fa7 	:	val_out <= 16'hafe4;
         16'h0fa8, 16'h0fa9, 16'h0faa, 16'h0fab, 16'h0fac, 16'h0fad, 16'h0fae, 16'h0faf 	:	val_out <= 16'haffb;
         16'h0fb0, 16'h0fb1, 16'h0fb2, 16'h0fb3, 16'h0fb4, 16'h0fb5, 16'h0fb6, 16'h0fb7 	:	val_out <= 16'hb013;
         16'h0fb8, 16'h0fb9, 16'h0fba, 16'h0fbb, 16'h0fbc, 16'h0fbd, 16'h0fbe, 16'h0fbf 	:	val_out <= 16'hb02a;
         16'h0fc0, 16'h0fc1, 16'h0fc2, 16'h0fc3, 16'h0fc4, 16'h0fc5, 16'h0fc6, 16'h0fc7 	:	val_out <= 16'hb041;
         16'h0fc8, 16'h0fc9, 16'h0fca, 16'h0fcb, 16'h0fcc, 16'h0fcd, 16'h0fce, 16'h0fcf 	:	val_out <= 16'hb059;
         16'h0fd0, 16'h0fd1, 16'h0fd2, 16'h0fd3, 16'h0fd4, 16'h0fd5, 16'h0fd6, 16'h0fd7 	:	val_out <= 16'hb070;
         16'h0fd8, 16'h0fd9, 16'h0fda, 16'h0fdb, 16'h0fdc, 16'h0fdd, 16'h0fde, 16'h0fdf 	:	val_out <= 16'hb087;
         16'h0fe0, 16'h0fe1, 16'h0fe2, 16'h0fe3, 16'h0fe4, 16'h0fe5, 16'h0fe6, 16'h0fe7 	:	val_out <= 16'hb09e;
         16'h0fe8, 16'h0fe9, 16'h0fea, 16'h0feb, 16'h0fec, 16'h0fed, 16'h0fee, 16'h0fef 	:	val_out <= 16'hb0b6;
         16'h0ff0, 16'h0ff1, 16'h0ff2, 16'h0ff3, 16'h0ff4, 16'h0ff5, 16'h0ff6, 16'h0ff7 	:	val_out <= 16'hb0cd;
         16'h0ff8, 16'h0ff9, 16'h0ffa, 16'h0ffb, 16'h0ffc, 16'h0ffd, 16'h0ffe, 16'h0fff 	:	val_out <= 16'hb0e4;
         16'h1000, 16'h1001, 16'h1002, 16'h1003, 16'h1004, 16'h1005, 16'h1006, 16'h1007 	:	val_out <= 16'hb0fb;
         16'h1008, 16'h1009, 16'h100a, 16'h100b, 16'h100c, 16'h100d, 16'h100e, 16'h100f 	:	val_out <= 16'hb112;
         16'h1010, 16'h1011, 16'h1012, 16'h1013, 16'h1014, 16'h1015, 16'h1016, 16'h1017 	:	val_out <= 16'hb12a;
         16'h1018, 16'h1019, 16'h101a, 16'h101b, 16'h101c, 16'h101d, 16'h101e, 16'h101f 	:	val_out <= 16'hb141;
         16'h1020, 16'h1021, 16'h1022, 16'h1023, 16'h1024, 16'h1025, 16'h1026, 16'h1027 	:	val_out <= 16'hb158;
         16'h1028, 16'h1029, 16'h102a, 16'h102b, 16'h102c, 16'h102d, 16'h102e, 16'h102f 	:	val_out <= 16'hb16f;
         16'h1030, 16'h1031, 16'h1032, 16'h1033, 16'h1034, 16'h1035, 16'h1036, 16'h1037 	:	val_out <= 16'hb186;
         16'h1038, 16'h1039, 16'h103a, 16'h103b, 16'h103c, 16'h103d, 16'h103e, 16'h103f 	:	val_out <= 16'hb19e;
         16'h1040, 16'h1041, 16'h1042, 16'h1043, 16'h1044, 16'h1045, 16'h1046, 16'h1047 	:	val_out <= 16'hb1b5;
         16'h1048, 16'h1049, 16'h104a, 16'h104b, 16'h104c, 16'h104d, 16'h104e, 16'h104f 	:	val_out <= 16'hb1cc;
         16'h1050, 16'h1051, 16'h1052, 16'h1053, 16'h1054, 16'h1055, 16'h1056, 16'h1057 	:	val_out <= 16'hb1e3;
         16'h1058, 16'h1059, 16'h105a, 16'h105b, 16'h105c, 16'h105d, 16'h105e, 16'h105f 	:	val_out <= 16'hb1fa;
         16'h1060, 16'h1061, 16'h1062, 16'h1063, 16'h1064, 16'h1065, 16'h1066, 16'h1067 	:	val_out <= 16'hb211;
         16'h1068, 16'h1069, 16'h106a, 16'h106b, 16'h106c, 16'h106d, 16'h106e, 16'h106f 	:	val_out <= 16'hb228;
         16'h1070, 16'h1071, 16'h1072, 16'h1073, 16'h1074, 16'h1075, 16'h1076, 16'h1077 	:	val_out <= 16'hb240;
         16'h1078, 16'h1079, 16'h107a, 16'h107b, 16'h107c, 16'h107d, 16'h107e, 16'h107f 	:	val_out <= 16'hb257;
         16'h1080, 16'h1081, 16'h1082, 16'h1083, 16'h1084, 16'h1085, 16'h1086, 16'h1087 	:	val_out <= 16'hb26e;
         16'h1088, 16'h1089, 16'h108a, 16'h108b, 16'h108c, 16'h108d, 16'h108e, 16'h108f 	:	val_out <= 16'hb285;
         16'h1090, 16'h1091, 16'h1092, 16'h1093, 16'h1094, 16'h1095, 16'h1096, 16'h1097 	:	val_out <= 16'hb29c;
         16'h1098, 16'h1099, 16'h109a, 16'h109b, 16'h109c, 16'h109d, 16'h109e, 16'h109f 	:	val_out <= 16'hb2b3;
         16'h10a0, 16'h10a1, 16'h10a2, 16'h10a3, 16'h10a4, 16'h10a5, 16'h10a6, 16'h10a7 	:	val_out <= 16'hb2ca;
         16'h10a8, 16'h10a9, 16'h10aa, 16'h10ab, 16'h10ac, 16'h10ad, 16'h10ae, 16'h10af 	:	val_out <= 16'hb2e1;
         16'h10b0, 16'h10b1, 16'h10b2, 16'h10b3, 16'h10b4, 16'h10b5, 16'h10b6, 16'h10b7 	:	val_out <= 16'hb2f8;
         16'h10b8, 16'h10b9, 16'h10ba, 16'h10bb, 16'h10bc, 16'h10bd, 16'h10be, 16'h10bf 	:	val_out <= 16'hb30f;
         16'h10c0, 16'h10c1, 16'h10c2, 16'h10c3, 16'h10c4, 16'h10c5, 16'h10c6, 16'h10c7 	:	val_out <= 16'hb326;
         16'h10c8, 16'h10c9, 16'h10ca, 16'h10cb, 16'h10cc, 16'h10cd, 16'h10ce, 16'h10cf 	:	val_out <= 16'hb33d;
         16'h10d0, 16'h10d1, 16'h10d2, 16'h10d3, 16'h10d4, 16'h10d5, 16'h10d6, 16'h10d7 	:	val_out <= 16'hb354;
         16'h10d8, 16'h10d9, 16'h10da, 16'h10db, 16'h10dc, 16'h10dd, 16'h10de, 16'h10df 	:	val_out <= 16'hb36b;
         16'h10e0, 16'h10e1, 16'h10e2, 16'h10e3, 16'h10e4, 16'h10e5, 16'h10e6, 16'h10e7 	:	val_out <= 16'hb382;
         16'h10e8, 16'h10e9, 16'h10ea, 16'h10eb, 16'h10ec, 16'h10ed, 16'h10ee, 16'h10ef 	:	val_out <= 16'hb399;
         16'h10f0, 16'h10f1, 16'h10f2, 16'h10f3, 16'h10f4, 16'h10f5, 16'h10f6, 16'h10f7 	:	val_out <= 16'hb3b0;
         16'h10f8, 16'h10f9, 16'h10fa, 16'h10fb, 16'h10fc, 16'h10fd, 16'h10fe, 16'h10ff 	:	val_out <= 16'hb3c7;
         16'h1100, 16'h1101, 16'h1102, 16'h1103, 16'h1104, 16'h1105, 16'h1106, 16'h1107 	:	val_out <= 16'hb3de;
         16'h1108, 16'h1109, 16'h110a, 16'h110b, 16'h110c, 16'h110d, 16'h110e, 16'h110f 	:	val_out <= 16'hb3f5;
         16'h1110, 16'h1111, 16'h1112, 16'h1113, 16'h1114, 16'h1115, 16'h1116, 16'h1117 	:	val_out <= 16'hb40c;
         16'h1118, 16'h1119, 16'h111a, 16'h111b, 16'h111c, 16'h111d, 16'h111e, 16'h111f 	:	val_out <= 16'hb423;
         16'h1120, 16'h1121, 16'h1122, 16'h1123, 16'h1124, 16'h1125, 16'h1126, 16'h1127 	:	val_out <= 16'hb43a;
         16'h1128, 16'h1129, 16'h112a, 16'h112b, 16'h112c, 16'h112d, 16'h112e, 16'h112f 	:	val_out <= 16'hb451;
         16'h1130, 16'h1131, 16'h1132, 16'h1133, 16'h1134, 16'h1135, 16'h1136, 16'h1137 	:	val_out <= 16'hb468;
         16'h1138, 16'h1139, 16'h113a, 16'h113b, 16'h113c, 16'h113d, 16'h113e, 16'h113f 	:	val_out <= 16'hb47f;
         16'h1140, 16'h1141, 16'h1142, 16'h1143, 16'h1144, 16'h1145, 16'h1146, 16'h1147 	:	val_out <= 16'hb496;
         16'h1148, 16'h1149, 16'h114a, 16'h114b, 16'h114c, 16'h114d, 16'h114e, 16'h114f 	:	val_out <= 16'hb4ad;
         16'h1150, 16'h1151, 16'h1152, 16'h1153, 16'h1154, 16'h1155, 16'h1156, 16'h1157 	:	val_out <= 16'hb4c4;
         16'h1158, 16'h1159, 16'h115a, 16'h115b, 16'h115c, 16'h115d, 16'h115e, 16'h115f 	:	val_out <= 16'hb4db;
         16'h1160, 16'h1161, 16'h1162, 16'h1163, 16'h1164, 16'h1165, 16'h1166, 16'h1167 	:	val_out <= 16'hb4f2;
         16'h1168, 16'h1169, 16'h116a, 16'h116b, 16'h116c, 16'h116d, 16'h116e, 16'h116f 	:	val_out <= 16'hb508;
         16'h1170, 16'h1171, 16'h1172, 16'h1173, 16'h1174, 16'h1175, 16'h1176, 16'h1177 	:	val_out <= 16'hb51f;
         16'h1178, 16'h1179, 16'h117a, 16'h117b, 16'h117c, 16'h117d, 16'h117e, 16'h117f 	:	val_out <= 16'hb536;
         16'h1180, 16'h1181, 16'h1182, 16'h1183, 16'h1184, 16'h1185, 16'h1186, 16'h1187 	:	val_out <= 16'hb54d;
         16'h1188, 16'h1189, 16'h118a, 16'h118b, 16'h118c, 16'h118d, 16'h118e, 16'h118f 	:	val_out <= 16'hb564;
         16'h1190, 16'h1191, 16'h1192, 16'h1193, 16'h1194, 16'h1195, 16'h1196, 16'h1197 	:	val_out <= 16'hb57b;
         16'h1198, 16'h1199, 16'h119a, 16'h119b, 16'h119c, 16'h119d, 16'h119e, 16'h119f 	:	val_out <= 16'hb592;
         16'h11a0, 16'h11a1, 16'h11a2, 16'h11a3, 16'h11a4, 16'h11a5, 16'h11a6, 16'h11a7 	:	val_out <= 16'hb5a8;
         16'h11a8, 16'h11a9, 16'h11aa, 16'h11ab, 16'h11ac, 16'h11ad, 16'h11ae, 16'h11af 	:	val_out <= 16'hb5bf;
         16'h11b0, 16'h11b1, 16'h11b2, 16'h11b3, 16'h11b4, 16'h11b5, 16'h11b6, 16'h11b7 	:	val_out <= 16'hb5d6;
         16'h11b8, 16'h11b9, 16'h11ba, 16'h11bb, 16'h11bc, 16'h11bd, 16'h11be, 16'h11bf 	:	val_out <= 16'hb5ed;
         16'h11c0, 16'h11c1, 16'h11c2, 16'h11c3, 16'h11c4, 16'h11c5, 16'h11c6, 16'h11c7 	:	val_out <= 16'hb604;
         16'h11c8, 16'h11c9, 16'h11ca, 16'h11cb, 16'h11cc, 16'h11cd, 16'h11ce, 16'h11cf 	:	val_out <= 16'hb61a;
         16'h11d0, 16'h11d1, 16'h11d2, 16'h11d3, 16'h11d4, 16'h11d5, 16'h11d6, 16'h11d7 	:	val_out <= 16'hb631;
         16'h11d8, 16'h11d9, 16'h11da, 16'h11db, 16'h11dc, 16'h11dd, 16'h11de, 16'h11df 	:	val_out <= 16'hb648;
         16'h11e0, 16'h11e1, 16'h11e2, 16'h11e3, 16'h11e4, 16'h11e5, 16'h11e6, 16'h11e7 	:	val_out <= 16'hb65f;
         16'h11e8, 16'h11e9, 16'h11ea, 16'h11eb, 16'h11ec, 16'h11ed, 16'h11ee, 16'h11ef 	:	val_out <= 16'hb675;
         16'h11f0, 16'h11f1, 16'h11f2, 16'h11f3, 16'h11f4, 16'h11f5, 16'h11f6, 16'h11f7 	:	val_out <= 16'hb68c;
         16'h11f8, 16'h11f9, 16'h11fa, 16'h11fb, 16'h11fc, 16'h11fd, 16'h11fe, 16'h11ff 	:	val_out <= 16'hb6a3;
         16'h1200, 16'h1201, 16'h1202, 16'h1203, 16'h1204, 16'h1205, 16'h1206, 16'h1207 	:	val_out <= 16'hb6ba;
         16'h1208, 16'h1209, 16'h120a, 16'h120b, 16'h120c, 16'h120d, 16'h120e, 16'h120f 	:	val_out <= 16'hb6d0;
         16'h1210, 16'h1211, 16'h1212, 16'h1213, 16'h1214, 16'h1215, 16'h1216, 16'h1217 	:	val_out <= 16'hb6e7;
         16'h1218, 16'h1219, 16'h121a, 16'h121b, 16'h121c, 16'h121d, 16'h121e, 16'h121f 	:	val_out <= 16'hb6fe;
         16'h1220, 16'h1221, 16'h1222, 16'h1223, 16'h1224, 16'h1225, 16'h1226, 16'h1227 	:	val_out <= 16'hb714;
         16'h1228, 16'h1229, 16'h122a, 16'h122b, 16'h122c, 16'h122d, 16'h122e, 16'h122f 	:	val_out <= 16'hb72b;
         16'h1230, 16'h1231, 16'h1232, 16'h1233, 16'h1234, 16'h1235, 16'h1236, 16'h1237 	:	val_out <= 16'hb742;
         16'h1238, 16'h1239, 16'h123a, 16'h123b, 16'h123c, 16'h123d, 16'h123e, 16'h123f 	:	val_out <= 16'hb758;
         16'h1240, 16'h1241, 16'h1242, 16'h1243, 16'h1244, 16'h1245, 16'h1246, 16'h1247 	:	val_out <= 16'hb76f;
         16'h1248, 16'h1249, 16'h124a, 16'h124b, 16'h124c, 16'h124d, 16'h124e, 16'h124f 	:	val_out <= 16'hb786;
         16'h1250, 16'h1251, 16'h1252, 16'h1253, 16'h1254, 16'h1255, 16'h1256, 16'h1257 	:	val_out <= 16'hb79c;
         16'h1258, 16'h1259, 16'h125a, 16'h125b, 16'h125c, 16'h125d, 16'h125e, 16'h125f 	:	val_out <= 16'hb7b3;
         16'h1260, 16'h1261, 16'h1262, 16'h1263, 16'h1264, 16'h1265, 16'h1266, 16'h1267 	:	val_out <= 16'hb7ca;
         16'h1268, 16'h1269, 16'h126a, 16'h126b, 16'h126c, 16'h126d, 16'h126e, 16'h126f 	:	val_out <= 16'hb7e0;
         16'h1270, 16'h1271, 16'h1272, 16'h1273, 16'h1274, 16'h1275, 16'h1276, 16'h1277 	:	val_out <= 16'hb7f7;
         16'h1278, 16'h1279, 16'h127a, 16'h127b, 16'h127c, 16'h127d, 16'h127e, 16'h127f 	:	val_out <= 16'hb80d;
         16'h1280, 16'h1281, 16'h1282, 16'h1283, 16'h1284, 16'h1285, 16'h1286, 16'h1287 	:	val_out <= 16'hb824;
         16'h1288, 16'h1289, 16'h128a, 16'h128b, 16'h128c, 16'h128d, 16'h128e, 16'h128f 	:	val_out <= 16'hb83b;
         16'h1290, 16'h1291, 16'h1292, 16'h1293, 16'h1294, 16'h1295, 16'h1296, 16'h1297 	:	val_out <= 16'hb851;
         16'h1298, 16'h1299, 16'h129a, 16'h129b, 16'h129c, 16'h129d, 16'h129e, 16'h129f 	:	val_out <= 16'hb868;
         16'h12a0, 16'h12a1, 16'h12a2, 16'h12a3, 16'h12a4, 16'h12a5, 16'h12a6, 16'h12a7 	:	val_out <= 16'hb87e;
         16'h12a8, 16'h12a9, 16'h12aa, 16'h12ab, 16'h12ac, 16'h12ad, 16'h12ae, 16'h12af 	:	val_out <= 16'hb895;
         16'h12b0, 16'h12b1, 16'h12b2, 16'h12b3, 16'h12b4, 16'h12b5, 16'h12b6, 16'h12b7 	:	val_out <= 16'hb8ab;
         16'h12b8, 16'h12b9, 16'h12ba, 16'h12bb, 16'h12bc, 16'h12bd, 16'h12be, 16'h12bf 	:	val_out <= 16'hb8c2;
         16'h12c0, 16'h12c1, 16'h12c2, 16'h12c3, 16'h12c4, 16'h12c5, 16'h12c6, 16'h12c7 	:	val_out <= 16'hb8d8;
         16'h12c8, 16'h12c9, 16'h12ca, 16'h12cb, 16'h12cc, 16'h12cd, 16'h12ce, 16'h12cf 	:	val_out <= 16'hb8ef;
         16'h12d0, 16'h12d1, 16'h12d2, 16'h12d3, 16'h12d4, 16'h12d5, 16'h12d6, 16'h12d7 	:	val_out <= 16'hb906;
         16'h12d8, 16'h12d9, 16'h12da, 16'h12db, 16'h12dc, 16'h12dd, 16'h12de, 16'h12df 	:	val_out <= 16'hb91c;
         16'h12e0, 16'h12e1, 16'h12e2, 16'h12e3, 16'h12e4, 16'h12e5, 16'h12e6, 16'h12e7 	:	val_out <= 16'hb932;
         16'h12e8, 16'h12e9, 16'h12ea, 16'h12eb, 16'h12ec, 16'h12ed, 16'h12ee, 16'h12ef 	:	val_out <= 16'hb949;
         16'h12f0, 16'h12f1, 16'h12f2, 16'h12f3, 16'h12f4, 16'h12f5, 16'h12f6, 16'h12f7 	:	val_out <= 16'hb95f;
         16'h12f8, 16'h12f9, 16'h12fa, 16'h12fb, 16'h12fc, 16'h12fd, 16'h12fe, 16'h12ff 	:	val_out <= 16'hb976;
         16'h1300, 16'h1301, 16'h1302, 16'h1303, 16'h1304, 16'h1305, 16'h1306, 16'h1307 	:	val_out <= 16'hb98c;
         16'h1308, 16'h1309, 16'h130a, 16'h130b, 16'h130c, 16'h130d, 16'h130e, 16'h130f 	:	val_out <= 16'hb9a3;
         16'h1310, 16'h1311, 16'h1312, 16'h1313, 16'h1314, 16'h1315, 16'h1316, 16'h1317 	:	val_out <= 16'hb9b9;
         16'h1318, 16'h1319, 16'h131a, 16'h131b, 16'h131c, 16'h131d, 16'h131e, 16'h131f 	:	val_out <= 16'hb9d0;
         16'h1320, 16'h1321, 16'h1322, 16'h1323, 16'h1324, 16'h1325, 16'h1326, 16'h1327 	:	val_out <= 16'hb9e6;
         16'h1328, 16'h1329, 16'h132a, 16'h132b, 16'h132c, 16'h132d, 16'h132e, 16'h132f 	:	val_out <= 16'hb9fd;
         16'h1330, 16'h1331, 16'h1332, 16'h1333, 16'h1334, 16'h1335, 16'h1336, 16'h1337 	:	val_out <= 16'hba13;
         16'h1338, 16'h1339, 16'h133a, 16'h133b, 16'h133c, 16'h133d, 16'h133e, 16'h133f 	:	val_out <= 16'hba29;
         16'h1340, 16'h1341, 16'h1342, 16'h1343, 16'h1344, 16'h1345, 16'h1346, 16'h1347 	:	val_out <= 16'hba40;
         16'h1348, 16'h1349, 16'h134a, 16'h134b, 16'h134c, 16'h134d, 16'h134e, 16'h134f 	:	val_out <= 16'hba56;
         16'h1350, 16'h1351, 16'h1352, 16'h1353, 16'h1354, 16'h1355, 16'h1356, 16'h1357 	:	val_out <= 16'hba6c;
         16'h1358, 16'h1359, 16'h135a, 16'h135b, 16'h135c, 16'h135d, 16'h135e, 16'h135f 	:	val_out <= 16'hba83;
         16'h1360, 16'h1361, 16'h1362, 16'h1363, 16'h1364, 16'h1365, 16'h1366, 16'h1367 	:	val_out <= 16'hba99;
         16'h1368, 16'h1369, 16'h136a, 16'h136b, 16'h136c, 16'h136d, 16'h136e, 16'h136f 	:	val_out <= 16'hbaaf;
         16'h1370, 16'h1371, 16'h1372, 16'h1373, 16'h1374, 16'h1375, 16'h1376, 16'h1377 	:	val_out <= 16'hbac6;
         16'h1378, 16'h1379, 16'h137a, 16'h137b, 16'h137c, 16'h137d, 16'h137e, 16'h137f 	:	val_out <= 16'hbadc;
         16'h1380, 16'h1381, 16'h1382, 16'h1383, 16'h1384, 16'h1385, 16'h1386, 16'h1387 	:	val_out <= 16'hbaf2;
         16'h1388, 16'h1389, 16'h138a, 16'h138b, 16'h138c, 16'h138d, 16'h138e, 16'h138f 	:	val_out <= 16'hbb09;
         16'h1390, 16'h1391, 16'h1392, 16'h1393, 16'h1394, 16'h1395, 16'h1396, 16'h1397 	:	val_out <= 16'hbb1f;
         16'h1398, 16'h1399, 16'h139a, 16'h139b, 16'h139c, 16'h139d, 16'h139e, 16'h139f 	:	val_out <= 16'hbb35;
         16'h13a0, 16'h13a1, 16'h13a2, 16'h13a3, 16'h13a4, 16'h13a5, 16'h13a6, 16'h13a7 	:	val_out <= 16'hbb4c;
         16'h13a8, 16'h13a9, 16'h13aa, 16'h13ab, 16'h13ac, 16'h13ad, 16'h13ae, 16'h13af 	:	val_out <= 16'hbb62;
         16'h13b0, 16'h13b1, 16'h13b2, 16'h13b3, 16'h13b4, 16'h13b5, 16'h13b6, 16'h13b7 	:	val_out <= 16'hbb78;
         16'h13b8, 16'h13b9, 16'h13ba, 16'h13bb, 16'h13bc, 16'h13bd, 16'h13be, 16'h13bf 	:	val_out <= 16'hbb8e;
         16'h13c0, 16'h13c1, 16'h13c2, 16'h13c3, 16'h13c4, 16'h13c5, 16'h13c6, 16'h13c7 	:	val_out <= 16'hbba5;
         16'h13c8, 16'h13c9, 16'h13ca, 16'h13cb, 16'h13cc, 16'h13cd, 16'h13ce, 16'h13cf 	:	val_out <= 16'hbbbb;
         16'h13d0, 16'h13d1, 16'h13d2, 16'h13d3, 16'h13d4, 16'h13d5, 16'h13d6, 16'h13d7 	:	val_out <= 16'hbbd1;
         16'h13d8, 16'h13d9, 16'h13da, 16'h13db, 16'h13dc, 16'h13dd, 16'h13de, 16'h13df 	:	val_out <= 16'hbbe7;
         16'h13e0, 16'h13e1, 16'h13e2, 16'h13e3, 16'h13e4, 16'h13e5, 16'h13e6, 16'h13e7 	:	val_out <= 16'hbbfd;
         16'h13e8, 16'h13e9, 16'h13ea, 16'h13eb, 16'h13ec, 16'h13ed, 16'h13ee, 16'h13ef 	:	val_out <= 16'hbc14;
         16'h13f0, 16'h13f1, 16'h13f2, 16'h13f3, 16'h13f4, 16'h13f5, 16'h13f6, 16'h13f7 	:	val_out <= 16'hbc2a;
         16'h13f8, 16'h13f9, 16'h13fa, 16'h13fb, 16'h13fc, 16'h13fd, 16'h13fe, 16'h13ff 	:	val_out <= 16'hbc40;
         16'h1400, 16'h1401, 16'h1402, 16'h1403, 16'h1404, 16'h1405, 16'h1406, 16'h1407 	:	val_out <= 16'hbc56;
         16'h1408, 16'h1409, 16'h140a, 16'h140b, 16'h140c, 16'h140d, 16'h140e, 16'h140f 	:	val_out <= 16'hbc6c;
         16'h1410, 16'h1411, 16'h1412, 16'h1413, 16'h1414, 16'h1415, 16'h1416, 16'h1417 	:	val_out <= 16'hbc83;
         16'h1418, 16'h1419, 16'h141a, 16'h141b, 16'h141c, 16'h141d, 16'h141e, 16'h141f 	:	val_out <= 16'hbc99;
         16'h1420, 16'h1421, 16'h1422, 16'h1423, 16'h1424, 16'h1425, 16'h1426, 16'h1427 	:	val_out <= 16'hbcaf;
         16'h1428, 16'h1429, 16'h142a, 16'h142b, 16'h142c, 16'h142d, 16'h142e, 16'h142f 	:	val_out <= 16'hbcc5;
         16'h1430, 16'h1431, 16'h1432, 16'h1433, 16'h1434, 16'h1435, 16'h1436, 16'h1437 	:	val_out <= 16'hbcdb;
         16'h1438, 16'h1439, 16'h143a, 16'h143b, 16'h143c, 16'h143d, 16'h143e, 16'h143f 	:	val_out <= 16'hbcf1;
         16'h1440, 16'h1441, 16'h1442, 16'h1443, 16'h1444, 16'h1445, 16'h1446, 16'h1447 	:	val_out <= 16'hbd07;
         16'h1448, 16'h1449, 16'h144a, 16'h144b, 16'h144c, 16'h144d, 16'h144e, 16'h144f 	:	val_out <= 16'hbd1d;
         16'h1450, 16'h1451, 16'h1452, 16'h1453, 16'h1454, 16'h1455, 16'h1456, 16'h1457 	:	val_out <= 16'hbd33;
         16'h1458, 16'h1459, 16'h145a, 16'h145b, 16'h145c, 16'h145d, 16'h145e, 16'h145f 	:	val_out <= 16'hbd49;
         16'h1460, 16'h1461, 16'h1462, 16'h1463, 16'h1464, 16'h1465, 16'h1466, 16'h1467 	:	val_out <= 16'hbd60;
         16'h1468, 16'h1469, 16'h146a, 16'h146b, 16'h146c, 16'h146d, 16'h146e, 16'h146f 	:	val_out <= 16'hbd76;
         16'h1470, 16'h1471, 16'h1472, 16'h1473, 16'h1474, 16'h1475, 16'h1476, 16'h1477 	:	val_out <= 16'hbd8c;
         16'h1478, 16'h1479, 16'h147a, 16'h147b, 16'h147c, 16'h147d, 16'h147e, 16'h147f 	:	val_out <= 16'hbda2;
         16'h1480, 16'h1481, 16'h1482, 16'h1483, 16'h1484, 16'h1485, 16'h1486, 16'h1487 	:	val_out <= 16'hbdb8;
         16'h1488, 16'h1489, 16'h148a, 16'h148b, 16'h148c, 16'h148d, 16'h148e, 16'h148f 	:	val_out <= 16'hbdce;
         16'h1490, 16'h1491, 16'h1492, 16'h1493, 16'h1494, 16'h1495, 16'h1496, 16'h1497 	:	val_out <= 16'hbde4;
         16'h1498, 16'h1499, 16'h149a, 16'h149b, 16'h149c, 16'h149d, 16'h149e, 16'h149f 	:	val_out <= 16'hbdfa;
         16'h14a0, 16'h14a1, 16'h14a2, 16'h14a3, 16'h14a4, 16'h14a5, 16'h14a6, 16'h14a7 	:	val_out <= 16'hbe10;
         16'h14a8, 16'h14a9, 16'h14aa, 16'h14ab, 16'h14ac, 16'h14ad, 16'h14ae, 16'h14af 	:	val_out <= 16'hbe26;
         16'h14b0, 16'h14b1, 16'h14b2, 16'h14b3, 16'h14b4, 16'h14b5, 16'h14b6, 16'h14b7 	:	val_out <= 16'hbe3c;
         16'h14b8, 16'h14b9, 16'h14ba, 16'h14bb, 16'h14bc, 16'h14bd, 16'h14be, 16'h14bf 	:	val_out <= 16'hbe52;
         16'h14c0, 16'h14c1, 16'h14c2, 16'h14c3, 16'h14c4, 16'h14c5, 16'h14c6, 16'h14c7 	:	val_out <= 16'hbe68;
         16'h14c8, 16'h14c9, 16'h14ca, 16'h14cb, 16'h14cc, 16'h14cd, 16'h14ce, 16'h14cf 	:	val_out <= 16'hbe7d;
         16'h14d0, 16'h14d1, 16'h14d2, 16'h14d3, 16'h14d4, 16'h14d5, 16'h14d6, 16'h14d7 	:	val_out <= 16'hbe93;
         16'h14d8, 16'h14d9, 16'h14da, 16'h14db, 16'h14dc, 16'h14dd, 16'h14de, 16'h14df 	:	val_out <= 16'hbea9;
         16'h14e0, 16'h14e1, 16'h14e2, 16'h14e3, 16'h14e4, 16'h14e5, 16'h14e6, 16'h14e7 	:	val_out <= 16'hbebf;
         16'h14e8, 16'h14e9, 16'h14ea, 16'h14eb, 16'h14ec, 16'h14ed, 16'h14ee, 16'h14ef 	:	val_out <= 16'hbed5;
         16'h14f0, 16'h14f1, 16'h14f2, 16'h14f3, 16'h14f4, 16'h14f5, 16'h14f6, 16'h14f7 	:	val_out <= 16'hbeeb;
         16'h14f8, 16'h14f9, 16'h14fa, 16'h14fb, 16'h14fc, 16'h14fd, 16'h14fe, 16'h14ff 	:	val_out <= 16'hbf01;
         16'h1500, 16'h1501, 16'h1502, 16'h1503, 16'h1504, 16'h1505, 16'h1506, 16'h1507 	:	val_out <= 16'hbf17;
         16'h1508, 16'h1509, 16'h150a, 16'h150b, 16'h150c, 16'h150d, 16'h150e, 16'h150f 	:	val_out <= 16'hbf2d;
         16'h1510, 16'h1511, 16'h1512, 16'h1513, 16'h1514, 16'h1515, 16'h1516, 16'h1517 	:	val_out <= 16'hbf43;
         16'h1518, 16'h1519, 16'h151a, 16'h151b, 16'h151c, 16'h151d, 16'h151e, 16'h151f 	:	val_out <= 16'hbf58;
         16'h1520, 16'h1521, 16'h1522, 16'h1523, 16'h1524, 16'h1525, 16'h1526, 16'h1527 	:	val_out <= 16'hbf6e;
         16'h1528, 16'h1529, 16'h152a, 16'h152b, 16'h152c, 16'h152d, 16'h152e, 16'h152f 	:	val_out <= 16'hbf84;
         16'h1530, 16'h1531, 16'h1532, 16'h1533, 16'h1534, 16'h1535, 16'h1536, 16'h1537 	:	val_out <= 16'hbf9a;
         16'h1538, 16'h1539, 16'h153a, 16'h153b, 16'h153c, 16'h153d, 16'h153e, 16'h153f 	:	val_out <= 16'hbfb0;
         16'h1540, 16'h1541, 16'h1542, 16'h1543, 16'h1544, 16'h1545, 16'h1546, 16'h1547 	:	val_out <= 16'hbfc5;
         16'h1548, 16'h1549, 16'h154a, 16'h154b, 16'h154c, 16'h154d, 16'h154e, 16'h154f 	:	val_out <= 16'hbfdb;
         16'h1550, 16'h1551, 16'h1552, 16'h1553, 16'h1554, 16'h1555, 16'h1556, 16'h1557 	:	val_out <= 16'hbff1;
         16'h1558, 16'h1559, 16'h155a, 16'h155b, 16'h155c, 16'h155d, 16'h155e, 16'h155f 	:	val_out <= 16'hc007;
         16'h1560, 16'h1561, 16'h1562, 16'h1563, 16'h1564, 16'h1565, 16'h1566, 16'h1567 	:	val_out <= 16'hc01d;
         16'h1568, 16'h1569, 16'h156a, 16'h156b, 16'h156c, 16'h156d, 16'h156e, 16'h156f 	:	val_out <= 16'hc032;
         16'h1570, 16'h1571, 16'h1572, 16'h1573, 16'h1574, 16'h1575, 16'h1576, 16'h1577 	:	val_out <= 16'hc048;
         16'h1578, 16'h1579, 16'h157a, 16'h157b, 16'h157c, 16'h157d, 16'h157e, 16'h157f 	:	val_out <= 16'hc05e;
         16'h1580, 16'h1581, 16'h1582, 16'h1583, 16'h1584, 16'h1585, 16'h1586, 16'h1587 	:	val_out <= 16'hc073;
         16'h1588, 16'h1589, 16'h158a, 16'h158b, 16'h158c, 16'h158d, 16'h158e, 16'h158f 	:	val_out <= 16'hc089;
         16'h1590, 16'h1591, 16'h1592, 16'h1593, 16'h1594, 16'h1595, 16'h1596, 16'h1597 	:	val_out <= 16'hc09f;
         16'h1598, 16'h1599, 16'h159a, 16'h159b, 16'h159c, 16'h159d, 16'h159e, 16'h159f 	:	val_out <= 16'hc0b5;
         16'h15a0, 16'h15a1, 16'h15a2, 16'h15a3, 16'h15a4, 16'h15a5, 16'h15a6, 16'h15a7 	:	val_out <= 16'hc0ca;
         16'h15a8, 16'h15a9, 16'h15aa, 16'h15ab, 16'h15ac, 16'h15ad, 16'h15ae, 16'h15af 	:	val_out <= 16'hc0e0;
         16'h15b0, 16'h15b1, 16'h15b2, 16'h15b3, 16'h15b4, 16'h15b5, 16'h15b6, 16'h15b7 	:	val_out <= 16'hc0f6;
         16'h15b8, 16'h15b9, 16'h15ba, 16'h15bb, 16'h15bc, 16'h15bd, 16'h15be, 16'h15bf 	:	val_out <= 16'hc10b;
         16'h15c0, 16'h15c1, 16'h15c2, 16'h15c3, 16'h15c4, 16'h15c5, 16'h15c6, 16'h15c7 	:	val_out <= 16'hc121;
         16'h15c8, 16'h15c9, 16'h15ca, 16'h15cb, 16'h15cc, 16'h15cd, 16'h15ce, 16'h15cf 	:	val_out <= 16'hc136;
         16'h15d0, 16'h15d1, 16'h15d2, 16'h15d3, 16'h15d4, 16'h15d5, 16'h15d6, 16'h15d7 	:	val_out <= 16'hc14c;
         16'h15d8, 16'h15d9, 16'h15da, 16'h15db, 16'h15dc, 16'h15dd, 16'h15de, 16'h15df 	:	val_out <= 16'hc162;
         16'h15e0, 16'h15e1, 16'h15e2, 16'h15e3, 16'h15e4, 16'h15e5, 16'h15e6, 16'h15e7 	:	val_out <= 16'hc177;
         16'h15e8, 16'h15e9, 16'h15ea, 16'h15eb, 16'h15ec, 16'h15ed, 16'h15ee, 16'h15ef 	:	val_out <= 16'hc18d;
         16'h15f0, 16'h15f1, 16'h15f2, 16'h15f3, 16'h15f4, 16'h15f5, 16'h15f6, 16'h15f7 	:	val_out <= 16'hc1a2;
         16'h15f8, 16'h15f9, 16'h15fa, 16'h15fb, 16'h15fc, 16'h15fd, 16'h15fe, 16'h15ff 	:	val_out <= 16'hc1b8;
         16'h1600, 16'h1601, 16'h1602, 16'h1603, 16'h1604, 16'h1605, 16'h1606, 16'h1607 	:	val_out <= 16'hc1ce;
         16'h1608, 16'h1609, 16'h160a, 16'h160b, 16'h160c, 16'h160d, 16'h160e, 16'h160f 	:	val_out <= 16'hc1e3;
         16'h1610, 16'h1611, 16'h1612, 16'h1613, 16'h1614, 16'h1615, 16'h1616, 16'h1617 	:	val_out <= 16'hc1f9;
         16'h1618, 16'h1619, 16'h161a, 16'h161b, 16'h161c, 16'h161d, 16'h161e, 16'h161f 	:	val_out <= 16'hc20e;
         16'h1620, 16'h1621, 16'h1622, 16'h1623, 16'h1624, 16'h1625, 16'h1626, 16'h1627 	:	val_out <= 16'hc224;
         16'h1628, 16'h1629, 16'h162a, 16'h162b, 16'h162c, 16'h162d, 16'h162e, 16'h162f 	:	val_out <= 16'hc239;
         16'h1630, 16'h1631, 16'h1632, 16'h1633, 16'h1634, 16'h1635, 16'h1636, 16'h1637 	:	val_out <= 16'hc24f;
         16'h1638, 16'h1639, 16'h163a, 16'h163b, 16'h163c, 16'h163d, 16'h163e, 16'h163f 	:	val_out <= 16'hc264;
         16'h1640, 16'h1641, 16'h1642, 16'h1643, 16'h1644, 16'h1645, 16'h1646, 16'h1647 	:	val_out <= 16'hc27a;
         16'h1648, 16'h1649, 16'h164a, 16'h164b, 16'h164c, 16'h164d, 16'h164e, 16'h164f 	:	val_out <= 16'hc28f;
         16'h1650, 16'h1651, 16'h1652, 16'h1653, 16'h1654, 16'h1655, 16'h1656, 16'h1657 	:	val_out <= 16'hc2a5;
         16'h1658, 16'h1659, 16'h165a, 16'h165b, 16'h165c, 16'h165d, 16'h165e, 16'h165f 	:	val_out <= 16'hc2ba;
         16'h1660, 16'h1661, 16'h1662, 16'h1663, 16'h1664, 16'h1665, 16'h1666, 16'h1667 	:	val_out <= 16'hc2d0;
         16'h1668, 16'h1669, 16'h166a, 16'h166b, 16'h166c, 16'h166d, 16'h166e, 16'h166f 	:	val_out <= 16'hc2e5;
         16'h1670, 16'h1671, 16'h1672, 16'h1673, 16'h1674, 16'h1675, 16'h1676, 16'h1677 	:	val_out <= 16'hc2fa;
         16'h1678, 16'h1679, 16'h167a, 16'h167b, 16'h167c, 16'h167d, 16'h167e, 16'h167f 	:	val_out <= 16'hc310;
         16'h1680, 16'h1681, 16'h1682, 16'h1683, 16'h1684, 16'h1685, 16'h1686, 16'h1687 	:	val_out <= 16'hc325;
         16'h1688, 16'h1689, 16'h168a, 16'h168b, 16'h168c, 16'h168d, 16'h168e, 16'h168f 	:	val_out <= 16'hc33b;
         16'h1690, 16'h1691, 16'h1692, 16'h1693, 16'h1694, 16'h1695, 16'h1696, 16'h1697 	:	val_out <= 16'hc350;
         16'h1698, 16'h1699, 16'h169a, 16'h169b, 16'h169c, 16'h169d, 16'h169e, 16'h169f 	:	val_out <= 16'hc365;
         16'h16a0, 16'h16a1, 16'h16a2, 16'h16a3, 16'h16a4, 16'h16a5, 16'h16a6, 16'h16a7 	:	val_out <= 16'hc37b;
         16'h16a8, 16'h16a9, 16'h16aa, 16'h16ab, 16'h16ac, 16'h16ad, 16'h16ae, 16'h16af 	:	val_out <= 16'hc390;
         16'h16b0, 16'h16b1, 16'h16b2, 16'h16b3, 16'h16b4, 16'h16b5, 16'h16b6, 16'h16b7 	:	val_out <= 16'hc3a5;
         16'h16b8, 16'h16b9, 16'h16ba, 16'h16bb, 16'h16bc, 16'h16bd, 16'h16be, 16'h16bf 	:	val_out <= 16'hc3bb;
         16'h16c0, 16'h16c1, 16'h16c2, 16'h16c3, 16'h16c4, 16'h16c5, 16'h16c6, 16'h16c7 	:	val_out <= 16'hc3d0;
         16'h16c8, 16'h16c9, 16'h16ca, 16'h16cb, 16'h16cc, 16'h16cd, 16'h16ce, 16'h16cf 	:	val_out <= 16'hc3e5;
         16'h16d0, 16'h16d1, 16'h16d2, 16'h16d3, 16'h16d4, 16'h16d5, 16'h16d6, 16'h16d7 	:	val_out <= 16'hc3fb;
         16'h16d8, 16'h16d9, 16'h16da, 16'h16db, 16'h16dc, 16'h16dd, 16'h16de, 16'h16df 	:	val_out <= 16'hc410;
         16'h16e0, 16'h16e1, 16'h16e2, 16'h16e3, 16'h16e4, 16'h16e5, 16'h16e6, 16'h16e7 	:	val_out <= 16'hc425;
         16'h16e8, 16'h16e9, 16'h16ea, 16'h16eb, 16'h16ec, 16'h16ed, 16'h16ee, 16'h16ef 	:	val_out <= 16'hc43b;
         16'h16f0, 16'h16f1, 16'h16f2, 16'h16f3, 16'h16f4, 16'h16f5, 16'h16f6, 16'h16f7 	:	val_out <= 16'hc450;
         16'h16f8, 16'h16f9, 16'h16fa, 16'h16fb, 16'h16fc, 16'h16fd, 16'h16fe, 16'h16ff 	:	val_out <= 16'hc465;
         16'h1700, 16'h1701, 16'h1702, 16'h1703, 16'h1704, 16'h1705, 16'h1706, 16'h1707 	:	val_out <= 16'hc47a;
         16'h1708, 16'h1709, 16'h170a, 16'h170b, 16'h170c, 16'h170d, 16'h170e, 16'h170f 	:	val_out <= 16'hc490;
         16'h1710, 16'h1711, 16'h1712, 16'h1713, 16'h1714, 16'h1715, 16'h1716, 16'h1717 	:	val_out <= 16'hc4a5;
         16'h1718, 16'h1719, 16'h171a, 16'h171b, 16'h171c, 16'h171d, 16'h171e, 16'h171f 	:	val_out <= 16'hc4ba;
         16'h1720, 16'h1721, 16'h1722, 16'h1723, 16'h1724, 16'h1725, 16'h1726, 16'h1727 	:	val_out <= 16'hc4cf;
         16'h1728, 16'h1729, 16'h172a, 16'h172b, 16'h172c, 16'h172d, 16'h172e, 16'h172f 	:	val_out <= 16'hc4e4;
         16'h1730, 16'h1731, 16'h1732, 16'h1733, 16'h1734, 16'h1735, 16'h1736, 16'h1737 	:	val_out <= 16'hc4fa;
         16'h1738, 16'h1739, 16'h173a, 16'h173b, 16'h173c, 16'h173d, 16'h173e, 16'h173f 	:	val_out <= 16'hc50f;
         16'h1740, 16'h1741, 16'h1742, 16'h1743, 16'h1744, 16'h1745, 16'h1746, 16'h1747 	:	val_out <= 16'hc524;
         16'h1748, 16'h1749, 16'h174a, 16'h174b, 16'h174c, 16'h174d, 16'h174e, 16'h174f 	:	val_out <= 16'hc539;
         16'h1750, 16'h1751, 16'h1752, 16'h1753, 16'h1754, 16'h1755, 16'h1756, 16'h1757 	:	val_out <= 16'hc54e;
         16'h1758, 16'h1759, 16'h175a, 16'h175b, 16'h175c, 16'h175d, 16'h175e, 16'h175f 	:	val_out <= 16'hc563;
         16'h1760, 16'h1761, 16'h1762, 16'h1763, 16'h1764, 16'h1765, 16'h1766, 16'h1767 	:	val_out <= 16'hc578;
         16'h1768, 16'h1769, 16'h176a, 16'h176b, 16'h176c, 16'h176d, 16'h176e, 16'h176f 	:	val_out <= 16'hc58d;
         16'h1770, 16'h1771, 16'h1772, 16'h1773, 16'h1774, 16'h1775, 16'h1776, 16'h1777 	:	val_out <= 16'hc5a3;
         16'h1778, 16'h1779, 16'h177a, 16'h177b, 16'h177c, 16'h177d, 16'h177e, 16'h177f 	:	val_out <= 16'hc5b8;
         16'h1780, 16'h1781, 16'h1782, 16'h1783, 16'h1784, 16'h1785, 16'h1786, 16'h1787 	:	val_out <= 16'hc5cd;
         16'h1788, 16'h1789, 16'h178a, 16'h178b, 16'h178c, 16'h178d, 16'h178e, 16'h178f 	:	val_out <= 16'hc5e2;
         16'h1790, 16'h1791, 16'h1792, 16'h1793, 16'h1794, 16'h1795, 16'h1796, 16'h1797 	:	val_out <= 16'hc5f7;
         16'h1798, 16'h1799, 16'h179a, 16'h179b, 16'h179c, 16'h179d, 16'h179e, 16'h179f 	:	val_out <= 16'hc60c;
         16'h17a0, 16'h17a1, 16'h17a2, 16'h17a3, 16'h17a4, 16'h17a5, 16'h17a6, 16'h17a7 	:	val_out <= 16'hc621;
         16'h17a8, 16'h17a9, 16'h17aa, 16'h17ab, 16'h17ac, 16'h17ad, 16'h17ae, 16'h17af 	:	val_out <= 16'hc636;
         16'h17b0, 16'h17b1, 16'h17b2, 16'h17b3, 16'h17b4, 16'h17b5, 16'h17b6, 16'h17b7 	:	val_out <= 16'hc64b;
         16'h17b8, 16'h17b9, 16'h17ba, 16'h17bb, 16'h17bc, 16'h17bd, 16'h17be, 16'h17bf 	:	val_out <= 16'hc660;
         16'h17c0, 16'h17c1, 16'h17c2, 16'h17c3, 16'h17c4, 16'h17c5, 16'h17c6, 16'h17c7 	:	val_out <= 16'hc675;
         16'h17c8, 16'h17c9, 16'h17ca, 16'h17cb, 16'h17cc, 16'h17cd, 16'h17ce, 16'h17cf 	:	val_out <= 16'hc68a;
         16'h17d0, 16'h17d1, 16'h17d2, 16'h17d3, 16'h17d4, 16'h17d5, 16'h17d6, 16'h17d7 	:	val_out <= 16'hc69f;
         16'h17d8, 16'h17d9, 16'h17da, 16'h17db, 16'h17dc, 16'h17dd, 16'h17de, 16'h17df 	:	val_out <= 16'hc6b4;
         16'h17e0, 16'h17e1, 16'h17e2, 16'h17e3, 16'h17e4, 16'h17e5, 16'h17e6, 16'h17e7 	:	val_out <= 16'hc6c9;
         16'h17e8, 16'h17e9, 16'h17ea, 16'h17eb, 16'h17ec, 16'h17ed, 16'h17ee, 16'h17ef 	:	val_out <= 16'hc6de;
         16'h17f0, 16'h17f1, 16'h17f2, 16'h17f3, 16'h17f4, 16'h17f5, 16'h17f6, 16'h17f7 	:	val_out <= 16'hc6f3;
         16'h17f8, 16'h17f9, 16'h17fa, 16'h17fb, 16'h17fc, 16'h17fd, 16'h17fe, 16'h17ff 	:	val_out <= 16'hc708;
         16'h1800, 16'h1801, 16'h1802, 16'h1803, 16'h1804, 16'h1805, 16'h1806, 16'h1807 	:	val_out <= 16'hc71c;
         16'h1808, 16'h1809, 16'h180a, 16'h180b, 16'h180c, 16'h180d, 16'h180e, 16'h180f 	:	val_out <= 16'hc731;
         16'h1810, 16'h1811, 16'h1812, 16'h1813, 16'h1814, 16'h1815, 16'h1816, 16'h1817 	:	val_out <= 16'hc746;
         16'h1818, 16'h1819, 16'h181a, 16'h181b, 16'h181c, 16'h181d, 16'h181e, 16'h181f 	:	val_out <= 16'hc75b;
         16'h1820, 16'h1821, 16'h1822, 16'h1823, 16'h1824, 16'h1825, 16'h1826, 16'h1827 	:	val_out <= 16'hc770;
         16'h1828, 16'h1829, 16'h182a, 16'h182b, 16'h182c, 16'h182d, 16'h182e, 16'h182f 	:	val_out <= 16'hc785;
         16'h1830, 16'h1831, 16'h1832, 16'h1833, 16'h1834, 16'h1835, 16'h1836, 16'h1837 	:	val_out <= 16'hc79a;
         16'h1838, 16'h1839, 16'h183a, 16'h183b, 16'h183c, 16'h183d, 16'h183e, 16'h183f 	:	val_out <= 16'hc7ae;
         16'h1840, 16'h1841, 16'h1842, 16'h1843, 16'h1844, 16'h1845, 16'h1846, 16'h1847 	:	val_out <= 16'hc7c3;
         16'h1848, 16'h1849, 16'h184a, 16'h184b, 16'h184c, 16'h184d, 16'h184e, 16'h184f 	:	val_out <= 16'hc7d8;
         16'h1850, 16'h1851, 16'h1852, 16'h1853, 16'h1854, 16'h1855, 16'h1856, 16'h1857 	:	val_out <= 16'hc7ed;
         16'h1858, 16'h1859, 16'h185a, 16'h185b, 16'h185c, 16'h185d, 16'h185e, 16'h185f 	:	val_out <= 16'hc802;
         16'h1860, 16'h1861, 16'h1862, 16'h1863, 16'h1864, 16'h1865, 16'h1866, 16'h1867 	:	val_out <= 16'hc816;
         16'h1868, 16'h1869, 16'h186a, 16'h186b, 16'h186c, 16'h186d, 16'h186e, 16'h186f 	:	val_out <= 16'hc82b;
         16'h1870, 16'h1871, 16'h1872, 16'h1873, 16'h1874, 16'h1875, 16'h1876, 16'h1877 	:	val_out <= 16'hc840;
         16'h1878, 16'h1879, 16'h187a, 16'h187b, 16'h187c, 16'h187d, 16'h187e, 16'h187f 	:	val_out <= 16'hc855;
         16'h1880, 16'h1881, 16'h1882, 16'h1883, 16'h1884, 16'h1885, 16'h1886, 16'h1887 	:	val_out <= 16'hc869;
         16'h1888, 16'h1889, 16'h188a, 16'h188b, 16'h188c, 16'h188d, 16'h188e, 16'h188f 	:	val_out <= 16'hc87e;
         16'h1890, 16'h1891, 16'h1892, 16'h1893, 16'h1894, 16'h1895, 16'h1896, 16'h1897 	:	val_out <= 16'hc893;
         16'h1898, 16'h1899, 16'h189a, 16'h189b, 16'h189c, 16'h189d, 16'h189e, 16'h189f 	:	val_out <= 16'hc8a8;
         16'h18a0, 16'h18a1, 16'h18a2, 16'h18a3, 16'h18a4, 16'h18a5, 16'h18a6, 16'h18a7 	:	val_out <= 16'hc8bc;
         16'h18a8, 16'h18a9, 16'h18aa, 16'h18ab, 16'h18ac, 16'h18ad, 16'h18ae, 16'h18af 	:	val_out <= 16'hc8d1;
         16'h18b0, 16'h18b1, 16'h18b2, 16'h18b3, 16'h18b4, 16'h18b5, 16'h18b6, 16'h18b7 	:	val_out <= 16'hc8e6;
         16'h18b8, 16'h18b9, 16'h18ba, 16'h18bb, 16'h18bc, 16'h18bd, 16'h18be, 16'h18bf 	:	val_out <= 16'hc8fa;
         16'h18c0, 16'h18c1, 16'h18c2, 16'h18c3, 16'h18c4, 16'h18c5, 16'h18c6, 16'h18c7 	:	val_out <= 16'hc90f;
         16'h18c8, 16'h18c9, 16'h18ca, 16'h18cb, 16'h18cc, 16'h18cd, 16'h18ce, 16'h18cf 	:	val_out <= 16'hc923;
         16'h18d0, 16'h18d1, 16'h18d2, 16'h18d3, 16'h18d4, 16'h18d5, 16'h18d6, 16'h18d7 	:	val_out <= 16'hc938;
         16'h18d8, 16'h18d9, 16'h18da, 16'h18db, 16'h18dc, 16'h18dd, 16'h18de, 16'h18df 	:	val_out <= 16'hc94d;
         16'h18e0, 16'h18e1, 16'h18e2, 16'h18e3, 16'h18e4, 16'h18e5, 16'h18e6, 16'h18e7 	:	val_out <= 16'hc961;
         16'h18e8, 16'h18e9, 16'h18ea, 16'h18eb, 16'h18ec, 16'h18ed, 16'h18ee, 16'h18ef 	:	val_out <= 16'hc976;
         16'h18f0, 16'h18f1, 16'h18f2, 16'h18f3, 16'h18f4, 16'h18f5, 16'h18f6, 16'h18f7 	:	val_out <= 16'hc98a;
         16'h18f8, 16'h18f9, 16'h18fa, 16'h18fb, 16'h18fc, 16'h18fd, 16'h18fe, 16'h18ff 	:	val_out <= 16'hc99f;
         16'h1900, 16'h1901, 16'h1902, 16'h1903, 16'h1904, 16'h1905, 16'h1906, 16'h1907 	:	val_out <= 16'hc9b4;
         16'h1908, 16'h1909, 16'h190a, 16'h190b, 16'h190c, 16'h190d, 16'h190e, 16'h190f 	:	val_out <= 16'hc9c8;
         16'h1910, 16'h1911, 16'h1912, 16'h1913, 16'h1914, 16'h1915, 16'h1916, 16'h1917 	:	val_out <= 16'hc9dd;
         16'h1918, 16'h1919, 16'h191a, 16'h191b, 16'h191c, 16'h191d, 16'h191e, 16'h191f 	:	val_out <= 16'hc9f1;
         16'h1920, 16'h1921, 16'h1922, 16'h1923, 16'h1924, 16'h1925, 16'h1926, 16'h1927 	:	val_out <= 16'hca06;
         16'h1928, 16'h1929, 16'h192a, 16'h192b, 16'h192c, 16'h192d, 16'h192e, 16'h192f 	:	val_out <= 16'hca1a;
         16'h1930, 16'h1931, 16'h1932, 16'h1933, 16'h1934, 16'h1935, 16'h1936, 16'h1937 	:	val_out <= 16'hca2f;
         16'h1938, 16'h1939, 16'h193a, 16'h193b, 16'h193c, 16'h193d, 16'h193e, 16'h193f 	:	val_out <= 16'hca43;
         16'h1940, 16'h1941, 16'h1942, 16'h1943, 16'h1944, 16'h1945, 16'h1946, 16'h1947 	:	val_out <= 16'hca58;
         16'h1948, 16'h1949, 16'h194a, 16'h194b, 16'h194c, 16'h194d, 16'h194e, 16'h194f 	:	val_out <= 16'hca6c;
         16'h1950, 16'h1951, 16'h1952, 16'h1953, 16'h1954, 16'h1955, 16'h1956, 16'h1957 	:	val_out <= 16'hca81;
         16'h1958, 16'h1959, 16'h195a, 16'h195b, 16'h195c, 16'h195d, 16'h195e, 16'h195f 	:	val_out <= 16'hca95;
         16'h1960, 16'h1961, 16'h1962, 16'h1963, 16'h1964, 16'h1965, 16'h1966, 16'h1967 	:	val_out <= 16'hcaa9;
         16'h1968, 16'h1969, 16'h196a, 16'h196b, 16'h196c, 16'h196d, 16'h196e, 16'h196f 	:	val_out <= 16'hcabe;
         16'h1970, 16'h1971, 16'h1972, 16'h1973, 16'h1974, 16'h1975, 16'h1976, 16'h1977 	:	val_out <= 16'hcad2;
         16'h1978, 16'h1979, 16'h197a, 16'h197b, 16'h197c, 16'h197d, 16'h197e, 16'h197f 	:	val_out <= 16'hcae7;
         16'h1980, 16'h1981, 16'h1982, 16'h1983, 16'h1984, 16'h1985, 16'h1986, 16'h1987 	:	val_out <= 16'hcafb;
         16'h1988, 16'h1989, 16'h198a, 16'h198b, 16'h198c, 16'h198d, 16'h198e, 16'h198f 	:	val_out <= 16'hcb0f;
         16'h1990, 16'h1991, 16'h1992, 16'h1993, 16'h1994, 16'h1995, 16'h1996, 16'h1997 	:	val_out <= 16'hcb24;
         16'h1998, 16'h1999, 16'h199a, 16'h199b, 16'h199c, 16'h199d, 16'h199e, 16'h199f 	:	val_out <= 16'hcb38;
         16'h19a0, 16'h19a1, 16'h19a2, 16'h19a3, 16'h19a4, 16'h19a5, 16'h19a6, 16'h19a7 	:	val_out <= 16'hcb4c;
         16'h19a8, 16'h19a9, 16'h19aa, 16'h19ab, 16'h19ac, 16'h19ad, 16'h19ae, 16'h19af 	:	val_out <= 16'hcb61;
         16'h19b0, 16'h19b1, 16'h19b2, 16'h19b3, 16'h19b4, 16'h19b5, 16'h19b6, 16'h19b7 	:	val_out <= 16'hcb75;
         16'h19b8, 16'h19b9, 16'h19ba, 16'h19bb, 16'h19bc, 16'h19bd, 16'h19be, 16'h19bf 	:	val_out <= 16'hcb89;
         16'h19c0, 16'h19c1, 16'h19c2, 16'h19c3, 16'h19c4, 16'h19c5, 16'h19c6, 16'h19c7 	:	val_out <= 16'hcb9e;
         16'h19c8, 16'h19c9, 16'h19ca, 16'h19cb, 16'h19cc, 16'h19cd, 16'h19ce, 16'h19cf 	:	val_out <= 16'hcbb2;
         16'h19d0, 16'h19d1, 16'h19d2, 16'h19d3, 16'h19d4, 16'h19d5, 16'h19d6, 16'h19d7 	:	val_out <= 16'hcbc6;
         16'h19d8, 16'h19d9, 16'h19da, 16'h19db, 16'h19dc, 16'h19dd, 16'h19de, 16'h19df 	:	val_out <= 16'hcbda;
         16'h19e0, 16'h19e1, 16'h19e2, 16'h19e3, 16'h19e4, 16'h19e5, 16'h19e6, 16'h19e7 	:	val_out <= 16'hcbef;
         16'h19e8, 16'h19e9, 16'h19ea, 16'h19eb, 16'h19ec, 16'h19ed, 16'h19ee, 16'h19ef 	:	val_out <= 16'hcc03;
         16'h19f0, 16'h19f1, 16'h19f2, 16'h19f3, 16'h19f4, 16'h19f5, 16'h19f6, 16'h19f7 	:	val_out <= 16'hcc17;
         16'h19f8, 16'h19f9, 16'h19fa, 16'h19fb, 16'h19fc, 16'h19fd, 16'h19fe, 16'h19ff 	:	val_out <= 16'hcc2b;
         16'h1a00, 16'h1a01, 16'h1a02, 16'h1a03, 16'h1a04, 16'h1a05, 16'h1a06, 16'h1a07 	:	val_out <= 16'hcc3f;
         16'h1a08, 16'h1a09, 16'h1a0a, 16'h1a0b, 16'h1a0c, 16'h1a0d, 16'h1a0e, 16'h1a0f 	:	val_out <= 16'hcc54;
         16'h1a10, 16'h1a11, 16'h1a12, 16'h1a13, 16'h1a14, 16'h1a15, 16'h1a16, 16'h1a17 	:	val_out <= 16'hcc68;
         16'h1a18, 16'h1a19, 16'h1a1a, 16'h1a1b, 16'h1a1c, 16'h1a1d, 16'h1a1e, 16'h1a1f 	:	val_out <= 16'hcc7c;
         16'h1a20, 16'h1a21, 16'h1a22, 16'h1a23, 16'h1a24, 16'h1a25, 16'h1a26, 16'h1a27 	:	val_out <= 16'hcc90;
         16'h1a28, 16'h1a29, 16'h1a2a, 16'h1a2b, 16'h1a2c, 16'h1a2d, 16'h1a2e, 16'h1a2f 	:	val_out <= 16'hcca4;
         16'h1a30, 16'h1a31, 16'h1a32, 16'h1a33, 16'h1a34, 16'h1a35, 16'h1a36, 16'h1a37 	:	val_out <= 16'hccb8;
         16'h1a38, 16'h1a39, 16'h1a3a, 16'h1a3b, 16'h1a3c, 16'h1a3d, 16'h1a3e, 16'h1a3f 	:	val_out <= 16'hcccc;
         16'h1a40, 16'h1a41, 16'h1a42, 16'h1a43, 16'h1a44, 16'h1a45, 16'h1a46, 16'h1a47 	:	val_out <= 16'hcce1;
         16'h1a48, 16'h1a49, 16'h1a4a, 16'h1a4b, 16'h1a4c, 16'h1a4d, 16'h1a4e, 16'h1a4f 	:	val_out <= 16'hccf5;
         16'h1a50, 16'h1a51, 16'h1a52, 16'h1a53, 16'h1a54, 16'h1a55, 16'h1a56, 16'h1a57 	:	val_out <= 16'hcd09;
         16'h1a58, 16'h1a59, 16'h1a5a, 16'h1a5b, 16'h1a5c, 16'h1a5d, 16'h1a5e, 16'h1a5f 	:	val_out <= 16'hcd1d;
         16'h1a60, 16'h1a61, 16'h1a62, 16'h1a63, 16'h1a64, 16'h1a65, 16'h1a66, 16'h1a67 	:	val_out <= 16'hcd31;
         16'h1a68, 16'h1a69, 16'h1a6a, 16'h1a6b, 16'h1a6c, 16'h1a6d, 16'h1a6e, 16'h1a6f 	:	val_out <= 16'hcd45;
         16'h1a70, 16'h1a71, 16'h1a72, 16'h1a73, 16'h1a74, 16'h1a75, 16'h1a76, 16'h1a77 	:	val_out <= 16'hcd59;
         16'h1a78, 16'h1a79, 16'h1a7a, 16'h1a7b, 16'h1a7c, 16'h1a7d, 16'h1a7e, 16'h1a7f 	:	val_out <= 16'hcd6d;
         16'h1a80, 16'h1a81, 16'h1a82, 16'h1a83, 16'h1a84, 16'h1a85, 16'h1a86, 16'h1a87 	:	val_out <= 16'hcd81;
         16'h1a88, 16'h1a89, 16'h1a8a, 16'h1a8b, 16'h1a8c, 16'h1a8d, 16'h1a8e, 16'h1a8f 	:	val_out <= 16'hcd95;
         16'h1a90, 16'h1a91, 16'h1a92, 16'h1a93, 16'h1a94, 16'h1a95, 16'h1a96, 16'h1a97 	:	val_out <= 16'hcda9;
         16'h1a98, 16'h1a99, 16'h1a9a, 16'h1a9b, 16'h1a9c, 16'h1a9d, 16'h1a9e, 16'h1a9f 	:	val_out <= 16'hcdbd;
         16'h1aa0, 16'h1aa1, 16'h1aa2, 16'h1aa3, 16'h1aa4, 16'h1aa5, 16'h1aa6, 16'h1aa7 	:	val_out <= 16'hcdd1;
         16'h1aa8, 16'h1aa9, 16'h1aaa, 16'h1aab, 16'h1aac, 16'h1aad, 16'h1aae, 16'h1aaf 	:	val_out <= 16'hcde5;
         16'h1ab0, 16'h1ab1, 16'h1ab2, 16'h1ab3, 16'h1ab4, 16'h1ab5, 16'h1ab6, 16'h1ab7 	:	val_out <= 16'hcdf9;
         16'h1ab8, 16'h1ab9, 16'h1aba, 16'h1abb, 16'h1abc, 16'h1abd, 16'h1abe, 16'h1abf 	:	val_out <= 16'hce0d;
         16'h1ac0, 16'h1ac1, 16'h1ac2, 16'h1ac3, 16'h1ac4, 16'h1ac5, 16'h1ac6, 16'h1ac7 	:	val_out <= 16'hce21;
         16'h1ac8, 16'h1ac9, 16'h1aca, 16'h1acb, 16'h1acc, 16'h1acd, 16'h1ace, 16'h1acf 	:	val_out <= 16'hce34;
         16'h1ad0, 16'h1ad1, 16'h1ad2, 16'h1ad3, 16'h1ad4, 16'h1ad5, 16'h1ad6, 16'h1ad7 	:	val_out <= 16'hce48;
         16'h1ad8, 16'h1ad9, 16'h1ada, 16'h1adb, 16'h1adc, 16'h1add, 16'h1ade, 16'h1adf 	:	val_out <= 16'hce5c;
         16'h1ae0, 16'h1ae1, 16'h1ae2, 16'h1ae3, 16'h1ae4, 16'h1ae5, 16'h1ae6, 16'h1ae7 	:	val_out <= 16'hce70;
         16'h1ae8, 16'h1ae9, 16'h1aea, 16'h1aeb, 16'h1aec, 16'h1aed, 16'h1aee, 16'h1aef 	:	val_out <= 16'hce84;
         16'h1af0, 16'h1af1, 16'h1af2, 16'h1af3, 16'h1af4, 16'h1af5, 16'h1af6, 16'h1af7 	:	val_out <= 16'hce98;
         16'h1af8, 16'h1af9, 16'h1afa, 16'h1afb, 16'h1afc, 16'h1afd, 16'h1afe, 16'h1aff 	:	val_out <= 16'hceac;
         16'h1b00, 16'h1b01, 16'h1b02, 16'h1b03, 16'h1b04, 16'h1b05, 16'h1b06, 16'h1b07 	:	val_out <= 16'hcebf;
         16'h1b08, 16'h1b09, 16'h1b0a, 16'h1b0b, 16'h1b0c, 16'h1b0d, 16'h1b0e, 16'h1b0f 	:	val_out <= 16'hced3;
         16'h1b10, 16'h1b11, 16'h1b12, 16'h1b13, 16'h1b14, 16'h1b15, 16'h1b16, 16'h1b17 	:	val_out <= 16'hcee7;
         16'h1b18, 16'h1b19, 16'h1b1a, 16'h1b1b, 16'h1b1c, 16'h1b1d, 16'h1b1e, 16'h1b1f 	:	val_out <= 16'hcefb;
         16'h1b20, 16'h1b21, 16'h1b22, 16'h1b23, 16'h1b24, 16'h1b25, 16'h1b26, 16'h1b27 	:	val_out <= 16'hcf0f;
         16'h1b28, 16'h1b29, 16'h1b2a, 16'h1b2b, 16'h1b2c, 16'h1b2d, 16'h1b2e, 16'h1b2f 	:	val_out <= 16'hcf22;
         16'h1b30, 16'h1b31, 16'h1b32, 16'h1b33, 16'h1b34, 16'h1b35, 16'h1b36, 16'h1b37 	:	val_out <= 16'hcf36;
         16'h1b38, 16'h1b39, 16'h1b3a, 16'h1b3b, 16'h1b3c, 16'h1b3d, 16'h1b3e, 16'h1b3f 	:	val_out <= 16'hcf4a;
         16'h1b40, 16'h1b41, 16'h1b42, 16'h1b43, 16'h1b44, 16'h1b45, 16'h1b46, 16'h1b47 	:	val_out <= 16'hcf5e;
         16'h1b48, 16'h1b49, 16'h1b4a, 16'h1b4b, 16'h1b4c, 16'h1b4d, 16'h1b4e, 16'h1b4f 	:	val_out <= 16'hcf71;
         16'h1b50, 16'h1b51, 16'h1b52, 16'h1b53, 16'h1b54, 16'h1b55, 16'h1b56, 16'h1b57 	:	val_out <= 16'hcf85;
         16'h1b58, 16'h1b59, 16'h1b5a, 16'h1b5b, 16'h1b5c, 16'h1b5d, 16'h1b5e, 16'h1b5f 	:	val_out <= 16'hcf99;
         16'h1b60, 16'h1b61, 16'h1b62, 16'h1b63, 16'h1b64, 16'h1b65, 16'h1b66, 16'h1b67 	:	val_out <= 16'hcfac;
         16'h1b68, 16'h1b69, 16'h1b6a, 16'h1b6b, 16'h1b6c, 16'h1b6d, 16'h1b6e, 16'h1b6f 	:	val_out <= 16'hcfc0;
         16'h1b70, 16'h1b71, 16'h1b72, 16'h1b73, 16'h1b74, 16'h1b75, 16'h1b76, 16'h1b77 	:	val_out <= 16'hcfd4;
         16'h1b78, 16'h1b79, 16'h1b7a, 16'h1b7b, 16'h1b7c, 16'h1b7d, 16'h1b7e, 16'h1b7f 	:	val_out <= 16'hcfe7;
         16'h1b80, 16'h1b81, 16'h1b82, 16'h1b83, 16'h1b84, 16'h1b85, 16'h1b86, 16'h1b87 	:	val_out <= 16'hcffb;
         16'h1b88, 16'h1b89, 16'h1b8a, 16'h1b8b, 16'h1b8c, 16'h1b8d, 16'h1b8e, 16'h1b8f 	:	val_out <= 16'hd00f;
         16'h1b90, 16'h1b91, 16'h1b92, 16'h1b93, 16'h1b94, 16'h1b95, 16'h1b96, 16'h1b97 	:	val_out <= 16'hd022;
         16'h1b98, 16'h1b99, 16'h1b9a, 16'h1b9b, 16'h1b9c, 16'h1b9d, 16'h1b9e, 16'h1b9f 	:	val_out <= 16'hd036;
         16'h1ba0, 16'h1ba1, 16'h1ba2, 16'h1ba3, 16'h1ba4, 16'h1ba5, 16'h1ba6, 16'h1ba7 	:	val_out <= 16'hd049;
         16'h1ba8, 16'h1ba9, 16'h1baa, 16'h1bab, 16'h1bac, 16'h1bad, 16'h1bae, 16'h1baf 	:	val_out <= 16'hd05d;
         16'h1bb0, 16'h1bb1, 16'h1bb2, 16'h1bb3, 16'h1bb4, 16'h1bb5, 16'h1bb6, 16'h1bb7 	:	val_out <= 16'hd070;
         16'h1bb8, 16'h1bb9, 16'h1bba, 16'h1bbb, 16'h1bbc, 16'h1bbd, 16'h1bbe, 16'h1bbf 	:	val_out <= 16'hd084;
         16'h1bc0, 16'h1bc1, 16'h1bc2, 16'h1bc3, 16'h1bc4, 16'h1bc5, 16'h1bc6, 16'h1bc7 	:	val_out <= 16'hd097;
         16'h1bc8, 16'h1bc9, 16'h1bca, 16'h1bcb, 16'h1bcc, 16'h1bcd, 16'h1bce, 16'h1bcf 	:	val_out <= 16'hd0ab;
         16'h1bd0, 16'h1bd1, 16'h1bd2, 16'h1bd3, 16'h1bd4, 16'h1bd5, 16'h1bd6, 16'h1bd7 	:	val_out <= 16'hd0bf;
         16'h1bd8, 16'h1bd9, 16'h1bda, 16'h1bdb, 16'h1bdc, 16'h1bdd, 16'h1bde, 16'h1bdf 	:	val_out <= 16'hd0d2;
         16'h1be0, 16'h1be1, 16'h1be2, 16'h1be3, 16'h1be4, 16'h1be5, 16'h1be6, 16'h1be7 	:	val_out <= 16'hd0e5;
         16'h1be8, 16'h1be9, 16'h1bea, 16'h1beb, 16'h1bec, 16'h1bed, 16'h1bee, 16'h1bef 	:	val_out <= 16'hd0f9;
         16'h1bf0, 16'h1bf1, 16'h1bf2, 16'h1bf3, 16'h1bf4, 16'h1bf5, 16'h1bf6, 16'h1bf7 	:	val_out <= 16'hd10c;
         16'h1bf8, 16'h1bf9, 16'h1bfa, 16'h1bfb, 16'h1bfc, 16'h1bfd, 16'h1bfe, 16'h1bff 	:	val_out <= 16'hd120;
         16'h1c00, 16'h1c01, 16'h1c02, 16'h1c03, 16'h1c04, 16'h1c05, 16'h1c06, 16'h1c07 	:	val_out <= 16'hd133;
         16'h1c08, 16'h1c09, 16'h1c0a, 16'h1c0b, 16'h1c0c, 16'h1c0d, 16'h1c0e, 16'h1c0f 	:	val_out <= 16'hd147;
         16'h1c10, 16'h1c11, 16'h1c12, 16'h1c13, 16'h1c14, 16'h1c15, 16'h1c16, 16'h1c17 	:	val_out <= 16'hd15a;
         16'h1c18, 16'h1c19, 16'h1c1a, 16'h1c1b, 16'h1c1c, 16'h1c1d, 16'h1c1e, 16'h1c1f 	:	val_out <= 16'hd16e;
         16'h1c20, 16'h1c21, 16'h1c22, 16'h1c23, 16'h1c24, 16'h1c25, 16'h1c26, 16'h1c27 	:	val_out <= 16'hd181;
         16'h1c28, 16'h1c29, 16'h1c2a, 16'h1c2b, 16'h1c2c, 16'h1c2d, 16'h1c2e, 16'h1c2f 	:	val_out <= 16'hd194;
         16'h1c30, 16'h1c31, 16'h1c32, 16'h1c33, 16'h1c34, 16'h1c35, 16'h1c36, 16'h1c37 	:	val_out <= 16'hd1a8;
         16'h1c38, 16'h1c39, 16'h1c3a, 16'h1c3b, 16'h1c3c, 16'h1c3d, 16'h1c3e, 16'h1c3f 	:	val_out <= 16'hd1bb;
         16'h1c40, 16'h1c41, 16'h1c42, 16'h1c43, 16'h1c44, 16'h1c45, 16'h1c46, 16'h1c47 	:	val_out <= 16'hd1ce;
         16'h1c48, 16'h1c49, 16'h1c4a, 16'h1c4b, 16'h1c4c, 16'h1c4d, 16'h1c4e, 16'h1c4f 	:	val_out <= 16'hd1e2;
         16'h1c50, 16'h1c51, 16'h1c52, 16'h1c53, 16'h1c54, 16'h1c55, 16'h1c56, 16'h1c57 	:	val_out <= 16'hd1f5;
         16'h1c58, 16'h1c59, 16'h1c5a, 16'h1c5b, 16'h1c5c, 16'h1c5d, 16'h1c5e, 16'h1c5f 	:	val_out <= 16'hd208;
         16'h1c60, 16'h1c61, 16'h1c62, 16'h1c63, 16'h1c64, 16'h1c65, 16'h1c66, 16'h1c67 	:	val_out <= 16'hd21c;
         16'h1c68, 16'h1c69, 16'h1c6a, 16'h1c6b, 16'h1c6c, 16'h1c6d, 16'h1c6e, 16'h1c6f 	:	val_out <= 16'hd22f;
         16'h1c70, 16'h1c71, 16'h1c72, 16'h1c73, 16'h1c74, 16'h1c75, 16'h1c76, 16'h1c77 	:	val_out <= 16'hd242;
         16'h1c78, 16'h1c79, 16'h1c7a, 16'h1c7b, 16'h1c7c, 16'h1c7d, 16'h1c7e, 16'h1c7f 	:	val_out <= 16'hd255;
         16'h1c80, 16'h1c81, 16'h1c82, 16'h1c83, 16'h1c84, 16'h1c85, 16'h1c86, 16'h1c87 	:	val_out <= 16'hd269;
         16'h1c88, 16'h1c89, 16'h1c8a, 16'h1c8b, 16'h1c8c, 16'h1c8d, 16'h1c8e, 16'h1c8f 	:	val_out <= 16'hd27c;
         16'h1c90, 16'h1c91, 16'h1c92, 16'h1c93, 16'h1c94, 16'h1c95, 16'h1c96, 16'h1c97 	:	val_out <= 16'hd28f;
         16'h1c98, 16'h1c99, 16'h1c9a, 16'h1c9b, 16'h1c9c, 16'h1c9d, 16'h1c9e, 16'h1c9f 	:	val_out <= 16'hd2a2;
         16'h1ca0, 16'h1ca1, 16'h1ca2, 16'h1ca3, 16'h1ca4, 16'h1ca5, 16'h1ca6, 16'h1ca7 	:	val_out <= 16'hd2b5;
         16'h1ca8, 16'h1ca9, 16'h1caa, 16'h1cab, 16'h1cac, 16'h1cad, 16'h1cae, 16'h1caf 	:	val_out <= 16'hd2c9;
         16'h1cb0, 16'h1cb1, 16'h1cb2, 16'h1cb3, 16'h1cb4, 16'h1cb5, 16'h1cb6, 16'h1cb7 	:	val_out <= 16'hd2dc;
         16'h1cb8, 16'h1cb9, 16'h1cba, 16'h1cbb, 16'h1cbc, 16'h1cbd, 16'h1cbe, 16'h1cbf 	:	val_out <= 16'hd2ef;
         16'h1cc0, 16'h1cc1, 16'h1cc2, 16'h1cc3, 16'h1cc4, 16'h1cc5, 16'h1cc6, 16'h1cc7 	:	val_out <= 16'hd302;
         16'h1cc8, 16'h1cc9, 16'h1cca, 16'h1ccb, 16'h1ccc, 16'h1ccd, 16'h1cce, 16'h1ccf 	:	val_out <= 16'hd315;
         16'h1cd0, 16'h1cd1, 16'h1cd2, 16'h1cd3, 16'h1cd4, 16'h1cd5, 16'h1cd6, 16'h1cd7 	:	val_out <= 16'hd328;
         16'h1cd8, 16'h1cd9, 16'h1cda, 16'h1cdb, 16'h1cdc, 16'h1cdd, 16'h1cde, 16'h1cdf 	:	val_out <= 16'hd33b;
         16'h1ce0, 16'h1ce1, 16'h1ce2, 16'h1ce3, 16'h1ce4, 16'h1ce5, 16'h1ce6, 16'h1ce7 	:	val_out <= 16'hd34e;
         16'h1ce8, 16'h1ce9, 16'h1cea, 16'h1ceb, 16'h1cec, 16'h1ced, 16'h1cee, 16'h1cef 	:	val_out <= 16'hd362;
         16'h1cf0, 16'h1cf1, 16'h1cf2, 16'h1cf3, 16'h1cf4, 16'h1cf5, 16'h1cf6, 16'h1cf7 	:	val_out <= 16'hd375;
         16'h1cf8, 16'h1cf9, 16'h1cfa, 16'h1cfb, 16'h1cfc, 16'h1cfd, 16'h1cfe, 16'h1cff 	:	val_out <= 16'hd388;
         16'h1d00, 16'h1d01, 16'h1d02, 16'h1d03, 16'h1d04, 16'h1d05, 16'h1d06, 16'h1d07 	:	val_out <= 16'hd39b;
         16'h1d08, 16'h1d09, 16'h1d0a, 16'h1d0b, 16'h1d0c, 16'h1d0d, 16'h1d0e, 16'h1d0f 	:	val_out <= 16'hd3ae;
         16'h1d10, 16'h1d11, 16'h1d12, 16'h1d13, 16'h1d14, 16'h1d15, 16'h1d16, 16'h1d17 	:	val_out <= 16'hd3c1;
         16'h1d18, 16'h1d19, 16'h1d1a, 16'h1d1b, 16'h1d1c, 16'h1d1d, 16'h1d1e, 16'h1d1f 	:	val_out <= 16'hd3d4;
         16'h1d20, 16'h1d21, 16'h1d22, 16'h1d23, 16'h1d24, 16'h1d25, 16'h1d26, 16'h1d27 	:	val_out <= 16'hd3e7;
         16'h1d28, 16'h1d29, 16'h1d2a, 16'h1d2b, 16'h1d2c, 16'h1d2d, 16'h1d2e, 16'h1d2f 	:	val_out <= 16'hd3fa;
         16'h1d30, 16'h1d31, 16'h1d32, 16'h1d33, 16'h1d34, 16'h1d35, 16'h1d36, 16'h1d37 	:	val_out <= 16'hd40d;
         16'h1d38, 16'h1d39, 16'h1d3a, 16'h1d3b, 16'h1d3c, 16'h1d3d, 16'h1d3e, 16'h1d3f 	:	val_out <= 16'hd420;
         16'h1d40, 16'h1d41, 16'h1d42, 16'h1d43, 16'h1d44, 16'h1d45, 16'h1d46, 16'h1d47 	:	val_out <= 16'hd433;
         16'h1d48, 16'h1d49, 16'h1d4a, 16'h1d4b, 16'h1d4c, 16'h1d4d, 16'h1d4e, 16'h1d4f 	:	val_out <= 16'hd445;
         16'h1d50, 16'h1d51, 16'h1d52, 16'h1d53, 16'h1d54, 16'h1d55, 16'h1d56, 16'h1d57 	:	val_out <= 16'hd458;
         16'h1d58, 16'h1d59, 16'h1d5a, 16'h1d5b, 16'h1d5c, 16'h1d5d, 16'h1d5e, 16'h1d5f 	:	val_out <= 16'hd46b;
         16'h1d60, 16'h1d61, 16'h1d62, 16'h1d63, 16'h1d64, 16'h1d65, 16'h1d66, 16'h1d67 	:	val_out <= 16'hd47e;
         16'h1d68, 16'h1d69, 16'h1d6a, 16'h1d6b, 16'h1d6c, 16'h1d6d, 16'h1d6e, 16'h1d6f 	:	val_out <= 16'hd491;
         16'h1d70, 16'h1d71, 16'h1d72, 16'h1d73, 16'h1d74, 16'h1d75, 16'h1d76, 16'h1d77 	:	val_out <= 16'hd4a4;
         16'h1d78, 16'h1d79, 16'h1d7a, 16'h1d7b, 16'h1d7c, 16'h1d7d, 16'h1d7e, 16'h1d7f 	:	val_out <= 16'hd4b7;
         16'h1d80, 16'h1d81, 16'h1d82, 16'h1d83, 16'h1d84, 16'h1d85, 16'h1d86, 16'h1d87 	:	val_out <= 16'hd4ca;
         16'h1d88, 16'h1d89, 16'h1d8a, 16'h1d8b, 16'h1d8c, 16'h1d8d, 16'h1d8e, 16'h1d8f 	:	val_out <= 16'hd4dc;
         16'h1d90, 16'h1d91, 16'h1d92, 16'h1d93, 16'h1d94, 16'h1d95, 16'h1d96, 16'h1d97 	:	val_out <= 16'hd4ef;
         16'h1d98, 16'h1d99, 16'h1d9a, 16'h1d9b, 16'h1d9c, 16'h1d9d, 16'h1d9e, 16'h1d9f 	:	val_out <= 16'hd502;
         16'h1da0, 16'h1da1, 16'h1da2, 16'h1da3, 16'h1da4, 16'h1da5, 16'h1da6, 16'h1da7 	:	val_out <= 16'hd515;
         16'h1da8, 16'h1da9, 16'h1daa, 16'h1dab, 16'h1dac, 16'h1dad, 16'h1dae, 16'h1daf 	:	val_out <= 16'hd528;
         16'h1db0, 16'h1db1, 16'h1db2, 16'h1db3, 16'h1db4, 16'h1db5, 16'h1db6, 16'h1db7 	:	val_out <= 16'hd53a;
         16'h1db8, 16'h1db9, 16'h1dba, 16'h1dbb, 16'h1dbc, 16'h1dbd, 16'h1dbe, 16'h1dbf 	:	val_out <= 16'hd54d;
         16'h1dc0, 16'h1dc1, 16'h1dc2, 16'h1dc3, 16'h1dc4, 16'h1dc5, 16'h1dc6, 16'h1dc7 	:	val_out <= 16'hd560;
         16'h1dc8, 16'h1dc9, 16'h1dca, 16'h1dcb, 16'h1dcc, 16'h1dcd, 16'h1dce, 16'h1dcf 	:	val_out <= 16'hd572;
         16'h1dd0, 16'h1dd1, 16'h1dd2, 16'h1dd3, 16'h1dd4, 16'h1dd5, 16'h1dd6, 16'h1dd7 	:	val_out <= 16'hd585;
         16'h1dd8, 16'h1dd9, 16'h1dda, 16'h1ddb, 16'h1ddc, 16'h1ddd, 16'h1dde, 16'h1ddf 	:	val_out <= 16'hd598;
         16'h1de0, 16'h1de1, 16'h1de2, 16'h1de3, 16'h1de4, 16'h1de5, 16'h1de6, 16'h1de7 	:	val_out <= 16'hd5ab;
         16'h1de8, 16'h1de9, 16'h1dea, 16'h1deb, 16'h1dec, 16'h1ded, 16'h1dee, 16'h1def 	:	val_out <= 16'hd5bd;
         16'h1df0, 16'h1df1, 16'h1df2, 16'h1df3, 16'h1df4, 16'h1df5, 16'h1df6, 16'h1df7 	:	val_out <= 16'hd5d0;
         16'h1df8, 16'h1df9, 16'h1dfa, 16'h1dfb, 16'h1dfc, 16'h1dfd, 16'h1dfe, 16'h1dff 	:	val_out <= 16'hd5e3;
         16'h1e00, 16'h1e01, 16'h1e02, 16'h1e03, 16'h1e04, 16'h1e05, 16'h1e06, 16'h1e07 	:	val_out <= 16'hd5f5;
         16'h1e08, 16'h1e09, 16'h1e0a, 16'h1e0b, 16'h1e0c, 16'h1e0d, 16'h1e0e, 16'h1e0f 	:	val_out <= 16'hd608;
         16'h1e10, 16'h1e11, 16'h1e12, 16'h1e13, 16'h1e14, 16'h1e15, 16'h1e16, 16'h1e17 	:	val_out <= 16'hd61a;
         16'h1e18, 16'h1e19, 16'h1e1a, 16'h1e1b, 16'h1e1c, 16'h1e1d, 16'h1e1e, 16'h1e1f 	:	val_out <= 16'hd62d;
         16'h1e20, 16'h1e21, 16'h1e22, 16'h1e23, 16'h1e24, 16'h1e25, 16'h1e26, 16'h1e27 	:	val_out <= 16'hd640;
         16'h1e28, 16'h1e29, 16'h1e2a, 16'h1e2b, 16'h1e2c, 16'h1e2d, 16'h1e2e, 16'h1e2f 	:	val_out <= 16'hd652;
         16'h1e30, 16'h1e31, 16'h1e32, 16'h1e33, 16'h1e34, 16'h1e35, 16'h1e36, 16'h1e37 	:	val_out <= 16'hd665;
         16'h1e38, 16'h1e39, 16'h1e3a, 16'h1e3b, 16'h1e3c, 16'h1e3d, 16'h1e3e, 16'h1e3f 	:	val_out <= 16'hd677;
         16'h1e40, 16'h1e41, 16'h1e42, 16'h1e43, 16'h1e44, 16'h1e45, 16'h1e46, 16'h1e47 	:	val_out <= 16'hd68a;
         16'h1e48, 16'h1e49, 16'h1e4a, 16'h1e4b, 16'h1e4c, 16'h1e4d, 16'h1e4e, 16'h1e4f 	:	val_out <= 16'hd69c;
         16'h1e50, 16'h1e51, 16'h1e52, 16'h1e53, 16'h1e54, 16'h1e55, 16'h1e56, 16'h1e57 	:	val_out <= 16'hd6af;
         16'h1e58, 16'h1e59, 16'h1e5a, 16'h1e5b, 16'h1e5c, 16'h1e5d, 16'h1e5e, 16'h1e5f 	:	val_out <= 16'hd6c1;
         16'h1e60, 16'h1e61, 16'h1e62, 16'h1e63, 16'h1e64, 16'h1e65, 16'h1e66, 16'h1e67 	:	val_out <= 16'hd6d4;
         16'h1e68, 16'h1e69, 16'h1e6a, 16'h1e6b, 16'h1e6c, 16'h1e6d, 16'h1e6e, 16'h1e6f 	:	val_out <= 16'hd6e6;
         16'h1e70, 16'h1e71, 16'h1e72, 16'h1e73, 16'h1e74, 16'h1e75, 16'h1e76, 16'h1e77 	:	val_out <= 16'hd6f9;
         16'h1e78, 16'h1e79, 16'h1e7a, 16'h1e7b, 16'h1e7c, 16'h1e7d, 16'h1e7e, 16'h1e7f 	:	val_out <= 16'hd70b;
         16'h1e80, 16'h1e81, 16'h1e82, 16'h1e83, 16'h1e84, 16'h1e85, 16'h1e86, 16'h1e87 	:	val_out <= 16'hd71d;
         16'h1e88, 16'h1e89, 16'h1e8a, 16'h1e8b, 16'h1e8c, 16'h1e8d, 16'h1e8e, 16'h1e8f 	:	val_out <= 16'hd730;
         16'h1e90, 16'h1e91, 16'h1e92, 16'h1e93, 16'h1e94, 16'h1e95, 16'h1e96, 16'h1e97 	:	val_out <= 16'hd742;
         16'h1e98, 16'h1e99, 16'h1e9a, 16'h1e9b, 16'h1e9c, 16'h1e9d, 16'h1e9e, 16'h1e9f 	:	val_out <= 16'hd755;
         16'h1ea0, 16'h1ea1, 16'h1ea2, 16'h1ea3, 16'h1ea4, 16'h1ea5, 16'h1ea6, 16'h1ea7 	:	val_out <= 16'hd767;
         16'h1ea8, 16'h1ea9, 16'h1eaa, 16'h1eab, 16'h1eac, 16'h1ead, 16'h1eae, 16'h1eaf 	:	val_out <= 16'hd779;
         16'h1eb0, 16'h1eb1, 16'h1eb2, 16'h1eb3, 16'h1eb4, 16'h1eb5, 16'h1eb6, 16'h1eb7 	:	val_out <= 16'hd78c;
         16'h1eb8, 16'h1eb9, 16'h1eba, 16'h1ebb, 16'h1ebc, 16'h1ebd, 16'h1ebe, 16'h1ebf 	:	val_out <= 16'hd79e;
         16'h1ec0, 16'h1ec1, 16'h1ec2, 16'h1ec3, 16'h1ec4, 16'h1ec5, 16'h1ec6, 16'h1ec7 	:	val_out <= 16'hd7b0;
         16'h1ec8, 16'h1ec9, 16'h1eca, 16'h1ecb, 16'h1ecc, 16'h1ecd, 16'h1ece, 16'h1ecf 	:	val_out <= 16'hd7c3;
         16'h1ed0, 16'h1ed1, 16'h1ed2, 16'h1ed3, 16'h1ed4, 16'h1ed5, 16'h1ed6, 16'h1ed7 	:	val_out <= 16'hd7d5;
         16'h1ed8, 16'h1ed9, 16'h1eda, 16'h1edb, 16'h1edc, 16'h1edd, 16'h1ede, 16'h1edf 	:	val_out <= 16'hd7e7;
         16'h1ee0, 16'h1ee1, 16'h1ee2, 16'h1ee3, 16'h1ee4, 16'h1ee5, 16'h1ee6, 16'h1ee7 	:	val_out <= 16'hd7f9;
         16'h1ee8, 16'h1ee9, 16'h1eea, 16'h1eeb, 16'h1eec, 16'h1eed, 16'h1eee, 16'h1eef 	:	val_out <= 16'hd80c;
         16'h1ef0, 16'h1ef1, 16'h1ef2, 16'h1ef3, 16'h1ef4, 16'h1ef5, 16'h1ef6, 16'h1ef7 	:	val_out <= 16'hd81e;
         16'h1ef8, 16'h1ef9, 16'h1efa, 16'h1efb, 16'h1efc, 16'h1efd, 16'h1efe, 16'h1eff 	:	val_out <= 16'hd830;
         16'h1f00, 16'h1f01, 16'h1f02, 16'h1f03, 16'h1f04, 16'h1f05, 16'h1f06, 16'h1f07 	:	val_out <= 16'hd842;
         16'h1f08, 16'h1f09, 16'h1f0a, 16'h1f0b, 16'h1f0c, 16'h1f0d, 16'h1f0e, 16'h1f0f 	:	val_out <= 16'hd855;
         16'h1f10, 16'h1f11, 16'h1f12, 16'h1f13, 16'h1f14, 16'h1f15, 16'h1f16, 16'h1f17 	:	val_out <= 16'hd867;
         16'h1f18, 16'h1f19, 16'h1f1a, 16'h1f1b, 16'h1f1c, 16'h1f1d, 16'h1f1e, 16'h1f1f 	:	val_out <= 16'hd879;
         16'h1f20, 16'h1f21, 16'h1f22, 16'h1f23, 16'h1f24, 16'h1f25, 16'h1f26, 16'h1f27 	:	val_out <= 16'hd88b;
         16'h1f28, 16'h1f29, 16'h1f2a, 16'h1f2b, 16'h1f2c, 16'h1f2d, 16'h1f2e, 16'h1f2f 	:	val_out <= 16'hd89d;
         16'h1f30, 16'h1f31, 16'h1f32, 16'h1f33, 16'h1f34, 16'h1f35, 16'h1f36, 16'h1f37 	:	val_out <= 16'hd8af;
         16'h1f38, 16'h1f39, 16'h1f3a, 16'h1f3b, 16'h1f3c, 16'h1f3d, 16'h1f3e, 16'h1f3f 	:	val_out <= 16'hd8c1;
         16'h1f40, 16'h1f41, 16'h1f42, 16'h1f43, 16'h1f44, 16'h1f45, 16'h1f46, 16'h1f47 	:	val_out <= 16'hd8d4;
         16'h1f48, 16'h1f49, 16'h1f4a, 16'h1f4b, 16'h1f4c, 16'h1f4d, 16'h1f4e, 16'h1f4f 	:	val_out <= 16'hd8e6;
         16'h1f50, 16'h1f51, 16'h1f52, 16'h1f53, 16'h1f54, 16'h1f55, 16'h1f56, 16'h1f57 	:	val_out <= 16'hd8f8;
         16'h1f58, 16'h1f59, 16'h1f5a, 16'h1f5b, 16'h1f5c, 16'h1f5d, 16'h1f5e, 16'h1f5f 	:	val_out <= 16'hd90a;
         16'h1f60, 16'h1f61, 16'h1f62, 16'h1f63, 16'h1f64, 16'h1f65, 16'h1f66, 16'h1f67 	:	val_out <= 16'hd91c;
         16'h1f68, 16'h1f69, 16'h1f6a, 16'h1f6b, 16'h1f6c, 16'h1f6d, 16'h1f6e, 16'h1f6f 	:	val_out <= 16'hd92e;
         16'h1f70, 16'h1f71, 16'h1f72, 16'h1f73, 16'h1f74, 16'h1f75, 16'h1f76, 16'h1f77 	:	val_out <= 16'hd940;
         16'h1f78, 16'h1f79, 16'h1f7a, 16'h1f7b, 16'h1f7c, 16'h1f7d, 16'h1f7e, 16'h1f7f 	:	val_out <= 16'hd952;
         16'h1f80, 16'h1f81, 16'h1f82, 16'h1f83, 16'h1f84, 16'h1f85, 16'h1f86, 16'h1f87 	:	val_out <= 16'hd964;
         16'h1f88, 16'h1f89, 16'h1f8a, 16'h1f8b, 16'h1f8c, 16'h1f8d, 16'h1f8e, 16'h1f8f 	:	val_out <= 16'hd976;
         16'h1f90, 16'h1f91, 16'h1f92, 16'h1f93, 16'h1f94, 16'h1f95, 16'h1f96, 16'h1f97 	:	val_out <= 16'hd988;
         16'h1f98, 16'h1f99, 16'h1f9a, 16'h1f9b, 16'h1f9c, 16'h1f9d, 16'h1f9e, 16'h1f9f 	:	val_out <= 16'hd99a;
         16'h1fa0, 16'h1fa1, 16'h1fa2, 16'h1fa3, 16'h1fa4, 16'h1fa5, 16'h1fa6, 16'h1fa7 	:	val_out <= 16'hd9ac;
         16'h1fa8, 16'h1fa9, 16'h1faa, 16'h1fab, 16'h1fac, 16'h1fad, 16'h1fae, 16'h1faf 	:	val_out <= 16'hd9be;
         16'h1fb0, 16'h1fb1, 16'h1fb2, 16'h1fb3, 16'h1fb4, 16'h1fb5, 16'h1fb6, 16'h1fb7 	:	val_out <= 16'hd9d0;
         16'h1fb8, 16'h1fb9, 16'h1fba, 16'h1fbb, 16'h1fbc, 16'h1fbd, 16'h1fbe, 16'h1fbf 	:	val_out <= 16'hd9e1;
         16'h1fc0, 16'h1fc1, 16'h1fc2, 16'h1fc3, 16'h1fc4, 16'h1fc5, 16'h1fc6, 16'h1fc7 	:	val_out <= 16'hd9f3;
         16'h1fc8, 16'h1fc9, 16'h1fca, 16'h1fcb, 16'h1fcc, 16'h1fcd, 16'h1fce, 16'h1fcf 	:	val_out <= 16'hda05;
         16'h1fd0, 16'h1fd1, 16'h1fd2, 16'h1fd3, 16'h1fd4, 16'h1fd5, 16'h1fd6, 16'h1fd7 	:	val_out <= 16'hda17;
         16'h1fd8, 16'h1fd9, 16'h1fda, 16'h1fdb, 16'h1fdc, 16'h1fdd, 16'h1fde, 16'h1fdf 	:	val_out <= 16'hda29;
         16'h1fe0, 16'h1fe1, 16'h1fe2, 16'h1fe3, 16'h1fe4, 16'h1fe5, 16'h1fe6, 16'h1fe7 	:	val_out <= 16'hda3b;
         16'h1fe8, 16'h1fe9, 16'h1fea, 16'h1feb, 16'h1fec, 16'h1fed, 16'h1fee, 16'h1fef 	:	val_out <= 16'hda4d;
         16'h1ff0, 16'h1ff1, 16'h1ff2, 16'h1ff3, 16'h1ff4, 16'h1ff5, 16'h1ff6, 16'h1ff7 	:	val_out <= 16'hda5e;
         16'h1ff8, 16'h1ff9, 16'h1ffa, 16'h1ffb, 16'h1ffc, 16'h1ffd, 16'h1ffe, 16'h1fff 	:	val_out <= 16'hda70;
         16'h2000, 16'h2001, 16'h2002, 16'h2003, 16'h2004, 16'h2005, 16'h2006, 16'h2007 	:	val_out <= 16'hda82;
         16'h2008, 16'h2009, 16'h200a, 16'h200b, 16'h200c, 16'h200d, 16'h200e, 16'h200f 	:	val_out <= 16'hda94;
         16'h2010, 16'h2011, 16'h2012, 16'h2013, 16'h2014, 16'h2015, 16'h2016, 16'h2017 	:	val_out <= 16'hdaa5;
         16'h2018, 16'h2019, 16'h201a, 16'h201b, 16'h201c, 16'h201d, 16'h201e, 16'h201f 	:	val_out <= 16'hdab7;
         16'h2020, 16'h2021, 16'h2022, 16'h2023, 16'h2024, 16'h2025, 16'h2026, 16'h2027 	:	val_out <= 16'hdac9;
         16'h2028, 16'h2029, 16'h202a, 16'h202b, 16'h202c, 16'h202d, 16'h202e, 16'h202f 	:	val_out <= 16'hdadb;
         16'h2030, 16'h2031, 16'h2032, 16'h2033, 16'h2034, 16'h2035, 16'h2036, 16'h2037 	:	val_out <= 16'hdaec;
         16'h2038, 16'h2039, 16'h203a, 16'h203b, 16'h203c, 16'h203d, 16'h203e, 16'h203f 	:	val_out <= 16'hdafe;
         16'h2040, 16'h2041, 16'h2042, 16'h2043, 16'h2044, 16'h2045, 16'h2046, 16'h2047 	:	val_out <= 16'hdb10;
         16'h2048, 16'h2049, 16'h204a, 16'h204b, 16'h204c, 16'h204d, 16'h204e, 16'h204f 	:	val_out <= 16'hdb21;
         16'h2050, 16'h2051, 16'h2052, 16'h2053, 16'h2054, 16'h2055, 16'h2056, 16'h2057 	:	val_out <= 16'hdb33;
         16'h2058, 16'h2059, 16'h205a, 16'h205b, 16'h205c, 16'h205d, 16'h205e, 16'h205f 	:	val_out <= 16'hdb45;
         16'h2060, 16'h2061, 16'h2062, 16'h2063, 16'h2064, 16'h2065, 16'h2066, 16'h2067 	:	val_out <= 16'hdb56;
         16'h2068, 16'h2069, 16'h206a, 16'h206b, 16'h206c, 16'h206d, 16'h206e, 16'h206f 	:	val_out <= 16'hdb68;
         16'h2070, 16'h2071, 16'h2072, 16'h2073, 16'h2074, 16'h2075, 16'h2076, 16'h2077 	:	val_out <= 16'hdb79;
         16'h2078, 16'h2079, 16'h207a, 16'h207b, 16'h207c, 16'h207d, 16'h207e, 16'h207f 	:	val_out <= 16'hdb8b;
         16'h2080, 16'h2081, 16'h2082, 16'h2083, 16'h2084, 16'h2085, 16'h2086, 16'h2087 	:	val_out <= 16'hdb9d;
         16'h2088, 16'h2089, 16'h208a, 16'h208b, 16'h208c, 16'h208d, 16'h208e, 16'h208f 	:	val_out <= 16'hdbae;
         16'h2090, 16'h2091, 16'h2092, 16'h2093, 16'h2094, 16'h2095, 16'h2096, 16'h2097 	:	val_out <= 16'hdbc0;
         16'h2098, 16'h2099, 16'h209a, 16'h209b, 16'h209c, 16'h209d, 16'h209e, 16'h209f 	:	val_out <= 16'hdbd1;
         16'h20a0, 16'h20a1, 16'h20a2, 16'h20a3, 16'h20a4, 16'h20a5, 16'h20a6, 16'h20a7 	:	val_out <= 16'hdbe3;
         16'h20a8, 16'h20a9, 16'h20aa, 16'h20ab, 16'h20ac, 16'h20ad, 16'h20ae, 16'h20af 	:	val_out <= 16'hdbf4;
         16'h20b0, 16'h20b1, 16'h20b2, 16'h20b3, 16'h20b4, 16'h20b5, 16'h20b6, 16'h20b7 	:	val_out <= 16'hdc06;
         16'h20b8, 16'h20b9, 16'h20ba, 16'h20bb, 16'h20bc, 16'h20bd, 16'h20be, 16'h20bf 	:	val_out <= 16'hdc17;
         16'h20c0, 16'h20c1, 16'h20c2, 16'h20c3, 16'h20c4, 16'h20c5, 16'h20c6, 16'h20c7 	:	val_out <= 16'hdc29;
         16'h20c8, 16'h20c9, 16'h20ca, 16'h20cb, 16'h20cc, 16'h20cd, 16'h20ce, 16'h20cf 	:	val_out <= 16'hdc3a;
         16'h20d0, 16'h20d1, 16'h20d2, 16'h20d3, 16'h20d4, 16'h20d5, 16'h20d6, 16'h20d7 	:	val_out <= 16'hdc4b;
         16'h20d8, 16'h20d9, 16'h20da, 16'h20db, 16'h20dc, 16'h20dd, 16'h20de, 16'h20df 	:	val_out <= 16'hdc5d;
         16'h20e0, 16'h20e1, 16'h20e2, 16'h20e3, 16'h20e4, 16'h20e5, 16'h20e6, 16'h20e7 	:	val_out <= 16'hdc6e;
         16'h20e8, 16'h20e9, 16'h20ea, 16'h20eb, 16'h20ec, 16'h20ed, 16'h20ee, 16'h20ef 	:	val_out <= 16'hdc80;
         16'h20f0, 16'h20f1, 16'h20f2, 16'h20f3, 16'h20f4, 16'h20f5, 16'h20f6, 16'h20f7 	:	val_out <= 16'hdc91;
         16'h20f8, 16'h20f9, 16'h20fa, 16'h20fb, 16'h20fc, 16'h20fd, 16'h20fe, 16'h20ff 	:	val_out <= 16'hdca2;
         16'h2100, 16'h2101, 16'h2102, 16'h2103, 16'h2104, 16'h2105, 16'h2106, 16'h2107 	:	val_out <= 16'hdcb4;
         16'h2108, 16'h2109, 16'h210a, 16'h210b, 16'h210c, 16'h210d, 16'h210e, 16'h210f 	:	val_out <= 16'hdcc5;
         16'h2110, 16'h2111, 16'h2112, 16'h2113, 16'h2114, 16'h2115, 16'h2116, 16'h2117 	:	val_out <= 16'hdcd6;
         16'h2118, 16'h2119, 16'h211a, 16'h211b, 16'h211c, 16'h211d, 16'h211e, 16'h211f 	:	val_out <= 16'hdce8;
         16'h2120, 16'h2121, 16'h2122, 16'h2123, 16'h2124, 16'h2125, 16'h2126, 16'h2127 	:	val_out <= 16'hdcf9;
         16'h2128, 16'h2129, 16'h212a, 16'h212b, 16'h212c, 16'h212d, 16'h212e, 16'h212f 	:	val_out <= 16'hdd0a;
         16'h2130, 16'h2131, 16'h2132, 16'h2133, 16'h2134, 16'h2135, 16'h2136, 16'h2137 	:	val_out <= 16'hdd1b;
         16'h2138, 16'h2139, 16'h213a, 16'h213b, 16'h213c, 16'h213d, 16'h213e, 16'h213f 	:	val_out <= 16'hdd2d;
         16'h2140, 16'h2141, 16'h2142, 16'h2143, 16'h2144, 16'h2145, 16'h2146, 16'h2147 	:	val_out <= 16'hdd3e;
         16'h2148, 16'h2149, 16'h214a, 16'h214b, 16'h214c, 16'h214d, 16'h214e, 16'h214f 	:	val_out <= 16'hdd4f;
         16'h2150, 16'h2151, 16'h2152, 16'h2153, 16'h2154, 16'h2155, 16'h2156, 16'h2157 	:	val_out <= 16'hdd60;
         16'h2158, 16'h2159, 16'h215a, 16'h215b, 16'h215c, 16'h215d, 16'h215e, 16'h215f 	:	val_out <= 16'hdd71;
         16'h2160, 16'h2161, 16'h2162, 16'h2163, 16'h2164, 16'h2165, 16'h2166, 16'h2167 	:	val_out <= 16'hdd83;
         16'h2168, 16'h2169, 16'h216a, 16'h216b, 16'h216c, 16'h216d, 16'h216e, 16'h216f 	:	val_out <= 16'hdd94;
         16'h2170, 16'h2171, 16'h2172, 16'h2173, 16'h2174, 16'h2175, 16'h2176, 16'h2177 	:	val_out <= 16'hdda5;
         16'h2178, 16'h2179, 16'h217a, 16'h217b, 16'h217c, 16'h217d, 16'h217e, 16'h217f 	:	val_out <= 16'hddb6;
         16'h2180, 16'h2181, 16'h2182, 16'h2183, 16'h2184, 16'h2185, 16'h2186, 16'h2187 	:	val_out <= 16'hddc7;
         16'h2188, 16'h2189, 16'h218a, 16'h218b, 16'h218c, 16'h218d, 16'h218e, 16'h218f 	:	val_out <= 16'hddd8;
         16'h2190, 16'h2191, 16'h2192, 16'h2193, 16'h2194, 16'h2195, 16'h2196, 16'h2197 	:	val_out <= 16'hdde9;
         16'h2198, 16'h2199, 16'h219a, 16'h219b, 16'h219c, 16'h219d, 16'h219e, 16'h219f 	:	val_out <= 16'hddfa;
         16'h21a0, 16'h21a1, 16'h21a2, 16'h21a3, 16'h21a4, 16'h21a5, 16'h21a6, 16'h21a7 	:	val_out <= 16'hde0b;
         16'h21a8, 16'h21a9, 16'h21aa, 16'h21ab, 16'h21ac, 16'h21ad, 16'h21ae, 16'h21af 	:	val_out <= 16'hde1c;
         16'h21b0, 16'h21b1, 16'h21b2, 16'h21b3, 16'h21b4, 16'h21b5, 16'h21b6, 16'h21b7 	:	val_out <= 16'hde2d;
         16'h21b8, 16'h21b9, 16'h21ba, 16'h21bb, 16'h21bc, 16'h21bd, 16'h21be, 16'h21bf 	:	val_out <= 16'hde3f;
         16'h21c0, 16'h21c1, 16'h21c2, 16'h21c3, 16'h21c4, 16'h21c5, 16'h21c6, 16'h21c7 	:	val_out <= 16'hde50;
         16'h21c8, 16'h21c9, 16'h21ca, 16'h21cb, 16'h21cc, 16'h21cd, 16'h21ce, 16'h21cf 	:	val_out <= 16'hde60;
         16'h21d0, 16'h21d1, 16'h21d2, 16'h21d3, 16'h21d4, 16'h21d5, 16'h21d6, 16'h21d7 	:	val_out <= 16'hde71;
         16'h21d8, 16'h21d9, 16'h21da, 16'h21db, 16'h21dc, 16'h21dd, 16'h21de, 16'h21df 	:	val_out <= 16'hde82;
         16'h21e0, 16'h21e1, 16'h21e2, 16'h21e3, 16'h21e4, 16'h21e5, 16'h21e6, 16'h21e7 	:	val_out <= 16'hde93;
         16'h21e8, 16'h21e9, 16'h21ea, 16'h21eb, 16'h21ec, 16'h21ed, 16'h21ee, 16'h21ef 	:	val_out <= 16'hdea4;
         16'h21f0, 16'h21f1, 16'h21f2, 16'h21f3, 16'h21f4, 16'h21f5, 16'h21f6, 16'h21f7 	:	val_out <= 16'hdeb5;
         16'h21f8, 16'h21f9, 16'h21fa, 16'h21fb, 16'h21fc, 16'h21fd, 16'h21fe, 16'h21ff 	:	val_out <= 16'hdec6;
         16'h2200, 16'h2201, 16'h2202, 16'h2203, 16'h2204, 16'h2205, 16'h2206, 16'h2207 	:	val_out <= 16'hded7;
         16'h2208, 16'h2209, 16'h220a, 16'h220b, 16'h220c, 16'h220d, 16'h220e, 16'h220f 	:	val_out <= 16'hdee8;
         16'h2210, 16'h2211, 16'h2212, 16'h2213, 16'h2214, 16'h2215, 16'h2216, 16'h2217 	:	val_out <= 16'hdef9;
         16'h2218, 16'h2219, 16'h221a, 16'h221b, 16'h221c, 16'h221d, 16'h221e, 16'h221f 	:	val_out <= 16'hdf0a;
         16'h2220, 16'h2221, 16'h2222, 16'h2223, 16'h2224, 16'h2225, 16'h2226, 16'h2227 	:	val_out <= 16'hdf1a;
         16'h2228, 16'h2229, 16'h222a, 16'h222b, 16'h222c, 16'h222d, 16'h222e, 16'h222f 	:	val_out <= 16'hdf2b;
         16'h2230, 16'h2231, 16'h2232, 16'h2233, 16'h2234, 16'h2235, 16'h2236, 16'h2237 	:	val_out <= 16'hdf3c;
         16'h2238, 16'h2239, 16'h223a, 16'h223b, 16'h223c, 16'h223d, 16'h223e, 16'h223f 	:	val_out <= 16'hdf4d;
         16'h2240, 16'h2241, 16'h2242, 16'h2243, 16'h2244, 16'h2245, 16'h2246, 16'h2247 	:	val_out <= 16'hdf5e;
         16'h2248, 16'h2249, 16'h224a, 16'h224b, 16'h224c, 16'h224d, 16'h224e, 16'h224f 	:	val_out <= 16'hdf6e;
         16'h2250, 16'h2251, 16'h2252, 16'h2253, 16'h2254, 16'h2255, 16'h2256, 16'h2257 	:	val_out <= 16'hdf7f;
         16'h2258, 16'h2259, 16'h225a, 16'h225b, 16'h225c, 16'h225d, 16'h225e, 16'h225f 	:	val_out <= 16'hdf90;
         16'h2260, 16'h2261, 16'h2262, 16'h2263, 16'h2264, 16'h2265, 16'h2266, 16'h2267 	:	val_out <= 16'hdfa0;
         16'h2268, 16'h2269, 16'h226a, 16'h226b, 16'h226c, 16'h226d, 16'h226e, 16'h226f 	:	val_out <= 16'hdfb1;
         16'h2270, 16'h2271, 16'h2272, 16'h2273, 16'h2274, 16'h2275, 16'h2276, 16'h2277 	:	val_out <= 16'hdfc2;
         16'h2278, 16'h2279, 16'h227a, 16'h227b, 16'h227c, 16'h227d, 16'h227e, 16'h227f 	:	val_out <= 16'hdfd3;
         16'h2280, 16'h2281, 16'h2282, 16'h2283, 16'h2284, 16'h2285, 16'h2286, 16'h2287 	:	val_out <= 16'hdfe3;
         16'h2288, 16'h2289, 16'h228a, 16'h228b, 16'h228c, 16'h228d, 16'h228e, 16'h228f 	:	val_out <= 16'hdff4;
         16'h2290, 16'h2291, 16'h2292, 16'h2293, 16'h2294, 16'h2295, 16'h2296, 16'h2297 	:	val_out <= 16'he004;
         16'h2298, 16'h2299, 16'h229a, 16'h229b, 16'h229c, 16'h229d, 16'h229e, 16'h229f 	:	val_out <= 16'he015;
         16'h22a0, 16'h22a1, 16'h22a2, 16'h22a3, 16'h22a4, 16'h22a5, 16'h22a6, 16'h22a7 	:	val_out <= 16'he026;
         16'h22a8, 16'h22a9, 16'h22aa, 16'h22ab, 16'h22ac, 16'h22ad, 16'h22ae, 16'h22af 	:	val_out <= 16'he036;
         16'h22b0, 16'h22b1, 16'h22b2, 16'h22b3, 16'h22b4, 16'h22b5, 16'h22b6, 16'h22b7 	:	val_out <= 16'he047;
         16'h22b8, 16'h22b9, 16'h22ba, 16'h22bb, 16'h22bc, 16'h22bd, 16'h22be, 16'h22bf 	:	val_out <= 16'he057;
         16'h22c0, 16'h22c1, 16'h22c2, 16'h22c3, 16'h22c4, 16'h22c5, 16'h22c6, 16'h22c7 	:	val_out <= 16'he068;
         16'h22c8, 16'h22c9, 16'h22ca, 16'h22cb, 16'h22cc, 16'h22cd, 16'h22ce, 16'h22cf 	:	val_out <= 16'he078;
         16'h22d0, 16'h22d1, 16'h22d2, 16'h22d3, 16'h22d4, 16'h22d5, 16'h22d6, 16'h22d7 	:	val_out <= 16'he089;
         16'h22d8, 16'h22d9, 16'h22da, 16'h22db, 16'h22dc, 16'h22dd, 16'h22de, 16'h22df 	:	val_out <= 16'he099;
         16'h22e0, 16'h22e1, 16'h22e2, 16'h22e3, 16'h22e4, 16'h22e5, 16'h22e6, 16'h22e7 	:	val_out <= 16'he0aa;
         16'h22e8, 16'h22e9, 16'h22ea, 16'h22eb, 16'h22ec, 16'h22ed, 16'h22ee, 16'h22ef 	:	val_out <= 16'he0ba;
         16'h22f0, 16'h22f1, 16'h22f2, 16'h22f3, 16'h22f4, 16'h22f5, 16'h22f6, 16'h22f7 	:	val_out <= 16'he0cb;
         16'h22f8, 16'h22f9, 16'h22fa, 16'h22fb, 16'h22fc, 16'h22fd, 16'h22fe, 16'h22ff 	:	val_out <= 16'he0db;
         16'h2300, 16'h2301, 16'h2302, 16'h2303, 16'h2304, 16'h2305, 16'h2306, 16'h2307 	:	val_out <= 16'he0ec;
         16'h2308, 16'h2309, 16'h230a, 16'h230b, 16'h230c, 16'h230d, 16'h230e, 16'h230f 	:	val_out <= 16'he0fc;
         16'h2310, 16'h2311, 16'h2312, 16'h2313, 16'h2314, 16'h2315, 16'h2316, 16'h2317 	:	val_out <= 16'he10d;
         16'h2318, 16'h2319, 16'h231a, 16'h231b, 16'h231c, 16'h231d, 16'h231e, 16'h231f 	:	val_out <= 16'he11d;
         16'h2320, 16'h2321, 16'h2322, 16'h2323, 16'h2324, 16'h2325, 16'h2326, 16'h2327 	:	val_out <= 16'he12d;
         16'h2328, 16'h2329, 16'h232a, 16'h232b, 16'h232c, 16'h232d, 16'h232e, 16'h232f 	:	val_out <= 16'he13e;
         16'h2330, 16'h2331, 16'h2332, 16'h2333, 16'h2334, 16'h2335, 16'h2336, 16'h2337 	:	val_out <= 16'he14e;
         16'h2338, 16'h2339, 16'h233a, 16'h233b, 16'h233c, 16'h233d, 16'h233e, 16'h233f 	:	val_out <= 16'he15e;
         16'h2340, 16'h2341, 16'h2342, 16'h2343, 16'h2344, 16'h2345, 16'h2346, 16'h2347 	:	val_out <= 16'he16f;
         16'h2348, 16'h2349, 16'h234a, 16'h234b, 16'h234c, 16'h234d, 16'h234e, 16'h234f 	:	val_out <= 16'he17f;
         16'h2350, 16'h2351, 16'h2352, 16'h2353, 16'h2354, 16'h2355, 16'h2356, 16'h2357 	:	val_out <= 16'he18f;
         16'h2358, 16'h2359, 16'h235a, 16'h235b, 16'h235c, 16'h235d, 16'h235e, 16'h235f 	:	val_out <= 16'he19f;
         16'h2360, 16'h2361, 16'h2362, 16'h2363, 16'h2364, 16'h2365, 16'h2366, 16'h2367 	:	val_out <= 16'he1b0;
         16'h2368, 16'h2369, 16'h236a, 16'h236b, 16'h236c, 16'h236d, 16'h236e, 16'h236f 	:	val_out <= 16'he1c0;
         16'h2370, 16'h2371, 16'h2372, 16'h2373, 16'h2374, 16'h2375, 16'h2376, 16'h2377 	:	val_out <= 16'he1d0;
         16'h2378, 16'h2379, 16'h237a, 16'h237b, 16'h237c, 16'h237d, 16'h237e, 16'h237f 	:	val_out <= 16'he1e0;
         16'h2380, 16'h2381, 16'h2382, 16'h2383, 16'h2384, 16'h2385, 16'h2386, 16'h2387 	:	val_out <= 16'he1f1;
         16'h2388, 16'h2389, 16'h238a, 16'h238b, 16'h238c, 16'h238d, 16'h238e, 16'h238f 	:	val_out <= 16'he201;
         16'h2390, 16'h2391, 16'h2392, 16'h2393, 16'h2394, 16'h2395, 16'h2396, 16'h2397 	:	val_out <= 16'he211;
         16'h2398, 16'h2399, 16'h239a, 16'h239b, 16'h239c, 16'h239d, 16'h239e, 16'h239f 	:	val_out <= 16'he221;
         16'h23a0, 16'h23a1, 16'h23a2, 16'h23a3, 16'h23a4, 16'h23a5, 16'h23a6, 16'h23a7 	:	val_out <= 16'he231;
         16'h23a8, 16'h23a9, 16'h23aa, 16'h23ab, 16'h23ac, 16'h23ad, 16'h23ae, 16'h23af 	:	val_out <= 16'he241;
         16'h23b0, 16'h23b1, 16'h23b2, 16'h23b3, 16'h23b4, 16'h23b5, 16'h23b6, 16'h23b7 	:	val_out <= 16'he251;
         16'h23b8, 16'h23b9, 16'h23ba, 16'h23bb, 16'h23bc, 16'h23bd, 16'h23be, 16'h23bf 	:	val_out <= 16'he261;
         16'h23c0, 16'h23c1, 16'h23c2, 16'h23c3, 16'h23c4, 16'h23c5, 16'h23c6, 16'h23c7 	:	val_out <= 16'he271;
         16'h23c8, 16'h23c9, 16'h23ca, 16'h23cb, 16'h23cc, 16'h23cd, 16'h23ce, 16'h23cf 	:	val_out <= 16'he282;
         16'h23d0, 16'h23d1, 16'h23d2, 16'h23d3, 16'h23d4, 16'h23d5, 16'h23d6, 16'h23d7 	:	val_out <= 16'he292;
         16'h23d8, 16'h23d9, 16'h23da, 16'h23db, 16'h23dc, 16'h23dd, 16'h23de, 16'h23df 	:	val_out <= 16'he2a2;
         16'h23e0, 16'h23e1, 16'h23e2, 16'h23e3, 16'h23e4, 16'h23e5, 16'h23e6, 16'h23e7 	:	val_out <= 16'he2b2;
         16'h23e8, 16'h23e9, 16'h23ea, 16'h23eb, 16'h23ec, 16'h23ed, 16'h23ee, 16'h23ef 	:	val_out <= 16'he2c2;
         16'h23f0, 16'h23f1, 16'h23f2, 16'h23f3, 16'h23f4, 16'h23f5, 16'h23f6, 16'h23f7 	:	val_out <= 16'he2d2;
         16'h23f8, 16'h23f9, 16'h23fa, 16'h23fb, 16'h23fc, 16'h23fd, 16'h23fe, 16'h23ff 	:	val_out <= 16'he2e2;
         16'h2400, 16'h2401, 16'h2402, 16'h2403, 16'h2404, 16'h2405, 16'h2406, 16'h2407 	:	val_out <= 16'he2f2;
         16'h2408, 16'h2409, 16'h240a, 16'h240b, 16'h240c, 16'h240d, 16'h240e, 16'h240f 	:	val_out <= 16'he301;
         16'h2410, 16'h2411, 16'h2412, 16'h2413, 16'h2414, 16'h2415, 16'h2416, 16'h2417 	:	val_out <= 16'he311;
         16'h2418, 16'h2419, 16'h241a, 16'h241b, 16'h241c, 16'h241d, 16'h241e, 16'h241f 	:	val_out <= 16'he321;
         16'h2420, 16'h2421, 16'h2422, 16'h2423, 16'h2424, 16'h2425, 16'h2426, 16'h2427 	:	val_out <= 16'he331;
         16'h2428, 16'h2429, 16'h242a, 16'h242b, 16'h242c, 16'h242d, 16'h242e, 16'h242f 	:	val_out <= 16'he341;
         16'h2430, 16'h2431, 16'h2432, 16'h2433, 16'h2434, 16'h2435, 16'h2436, 16'h2437 	:	val_out <= 16'he351;
         16'h2438, 16'h2439, 16'h243a, 16'h243b, 16'h243c, 16'h243d, 16'h243e, 16'h243f 	:	val_out <= 16'he361;
         16'h2440, 16'h2441, 16'h2442, 16'h2443, 16'h2444, 16'h2445, 16'h2446, 16'h2447 	:	val_out <= 16'he371;
         16'h2448, 16'h2449, 16'h244a, 16'h244b, 16'h244c, 16'h244d, 16'h244e, 16'h244f 	:	val_out <= 16'he380;
         16'h2450, 16'h2451, 16'h2452, 16'h2453, 16'h2454, 16'h2455, 16'h2456, 16'h2457 	:	val_out <= 16'he390;
         16'h2458, 16'h2459, 16'h245a, 16'h245b, 16'h245c, 16'h245d, 16'h245e, 16'h245f 	:	val_out <= 16'he3a0;
         16'h2460, 16'h2461, 16'h2462, 16'h2463, 16'h2464, 16'h2465, 16'h2466, 16'h2467 	:	val_out <= 16'he3b0;
         16'h2468, 16'h2469, 16'h246a, 16'h246b, 16'h246c, 16'h246d, 16'h246e, 16'h246f 	:	val_out <= 16'he3c0;
         16'h2470, 16'h2471, 16'h2472, 16'h2473, 16'h2474, 16'h2475, 16'h2476, 16'h2477 	:	val_out <= 16'he3cf;
         16'h2478, 16'h2479, 16'h247a, 16'h247b, 16'h247c, 16'h247d, 16'h247e, 16'h247f 	:	val_out <= 16'he3df;
         16'h2480, 16'h2481, 16'h2482, 16'h2483, 16'h2484, 16'h2485, 16'h2486, 16'h2487 	:	val_out <= 16'he3ef;
         16'h2488, 16'h2489, 16'h248a, 16'h248b, 16'h248c, 16'h248d, 16'h248e, 16'h248f 	:	val_out <= 16'he3fe;
         16'h2490, 16'h2491, 16'h2492, 16'h2493, 16'h2494, 16'h2495, 16'h2496, 16'h2497 	:	val_out <= 16'he40e;
         16'h2498, 16'h2499, 16'h249a, 16'h249b, 16'h249c, 16'h249d, 16'h249e, 16'h249f 	:	val_out <= 16'he41e;
         16'h24a0, 16'h24a1, 16'h24a2, 16'h24a3, 16'h24a4, 16'h24a5, 16'h24a6, 16'h24a7 	:	val_out <= 16'he42d;
         16'h24a8, 16'h24a9, 16'h24aa, 16'h24ab, 16'h24ac, 16'h24ad, 16'h24ae, 16'h24af 	:	val_out <= 16'he43d;
         16'h24b0, 16'h24b1, 16'h24b2, 16'h24b3, 16'h24b4, 16'h24b5, 16'h24b6, 16'h24b7 	:	val_out <= 16'he44d;
         16'h24b8, 16'h24b9, 16'h24ba, 16'h24bb, 16'h24bc, 16'h24bd, 16'h24be, 16'h24bf 	:	val_out <= 16'he45c;
         16'h24c0, 16'h24c1, 16'h24c2, 16'h24c3, 16'h24c4, 16'h24c5, 16'h24c6, 16'h24c7 	:	val_out <= 16'he46c;
         16'h24c8, 16'h24c9, 16'h24ca, 16'h24cb, 16'h24cc, 16'h24cd, 16'h24ce, 16'h24cf 	:	val_out <= 16'he47b;
         16'h24d0, 16'h24d1, 16'h24d2, 16'h24d3, 16'h24d4, 16'h24d5, 16'h24d6, 16'h24d7 	:	val_out <= 16'he48b;
         16'h24d8, 16'h24d9, 16'h24da, 16'h24db, 16'h24dc, 16'h24dd, 16'h24de, 16'h24df 	:	val_out <= 16'he49b;
         16'h24e0, 16'h24e1, 16'h24e2, 16'h24e3, 16'h24e4, 16'h24e5, 16'h24e6, 16'h24e7 	:	val_out <= 16'he4aa;
         16'h24e8, 16'h24e9, 16'h24ea, 16'h24eb, 16'h24ec, 16'h24ed, 16'h24ee, 16'h24ef 	:	val_out <= 16'he4ba;
         16'h24f0, 16'h24f1, 16'h24f2, 16'h24f3, 16'h24f4, 16'h24f5, 16'h24f6, 16'h24f7 	:	val_out <= 16'he4c9;
         16'h24f8, 16'h24f9, 16'h24fa, 16'h24fb, 16'h24fc, 16'h24fd, 16'h24fe, 16'h24ff 	:	val_out <= 16'he4d9;
         16'h2500, 16'h2501, 16'h2502, 16'h2503, 16'h2504, 16'h2505, 16'h2506, 16'h2507 	:	val_out <= 16'he4e8;
         16'h2508, 16'h2509, 16'h250a, 16'h250b, 16'h250c, 16'h250d, 16'h250e, 16'h250f 	:	val_out <= 16'he4f7;
         16'h2510, 16'h2511, 16'h2512, 16'h2513, 16'h2514, 16'h2515, 16'h2516, 16'h2517 	:	val_out <= 16'he507;
         16'h2518, 16'h2519, 16'h251a, 16'h251b, 16'h251c, 16'h251d, 16'h251e, 16'h251f 	:	val_out <= 16'he516;
         16'h2520, 16'h2521, 16'h2522, 16'h2523, 16'h2524, 16'h2525, 16'h2526, 16'h2527 	:	val_out <= 16'he526;
         16'h2528, 16'h2529, 16'h252a, 16'h252b, 16'h252c, 16'h252d, 16'h252e, 16'h252f 	:	val_out <= 16'he535;
         16'h2530, 16'h2531, 16'h2532, 16'h2533, 16'h2534, 16'h2535, 16'h2536, 16'h2537 	:	val_out <= 16'he545;
         16'h2538, 16'h2539, 16'h253a, 16'h253b, 16'h253c, 16'h253d, 16'h253e, 16'h253f 	:	val_out <= 16'he554;
         16'h2540, 16'h2541, 16'h2542, 16'h2543, 16'h2544, 16'h2545, 16'h2546, 16'h2547 	:	val_out <= 16'he563;
         16'h2548, 16'h2549, 16'h254a, 16'h254b, 16'h254c, 16'h254d, 16'h254e, 16'h254f 	:	val_out <= 16'he573;
         16'h2550, 16'h2551, 16'h2552, 16'h2553, 16'h2554, 16'h2555, 16'h2556, 16'h2557 	:	val_out <= 16'he582;
         16'h2558, 16'h2559, 16'h255a, 16'h255b, 16'h255c, 16'h255d, 16'h255e, 16'h255f 	:	val_out <= 16'he591;
         16'h2560, 16'h2561, 16'h2562, 16'h2563, 16'h2564, 16'h2565, 16'h2566, 16'h2567 	:	val_out <= 16'he5a0;
         16'h2568, 16'h2569, 16'h256a, 16'h256b, 16'h256c, 16'h256d, 16'h256e, 16'h256f 	:	val_out <= 16'he5b0;
         16'h2570, 16'h2571, 16'h2572, 16'h2573, 16'h2574, 16'h2575, 16'h2576, 16'h2577 	:	val_out <= 16'he5bf;
         16'h2578, 16'h2579, 16'h257a, 16'h257b, 16'h257c, 16'h257d, 16'h257e, 16'h257f 	:	val_out <= 16'he5ce;
         16'h2580, 16'h2581, 16'h2582, 16'h2583, 16'h2584, 16'h2585, 16'h2586, 16'h2587 	:	val_out <= 16'he5dd;
         16'h2588, 16'h2589, 16'h258a, 16'h258b, 16'h258c, 16'h258d, 16'h258e, 16'h258f 	:	val_out <= 16'he5ed;
         16'h2590, 16'h2591, 16'h2592, 16'h2593, 16'h2594, 16'h2595, 16'h2596, 16'h2597 	:	val_out <= 16'he5fc;
         16'h2598, 16'h2599, 16'h259a, 16'h259b, 16'h259c, 16'h259d, 16'h259e, 16'h259f 	:	val_out <= 16'he60b;
         16'h25a0, 16'h25a1, 16'h25a2, 16'h25a3, 16'h25a4, 16'h25a5, 16'h25a6, 16'h25a7 	:	val_out <= 16'he61a;
         16'h25a8, 16'h25a9, 16'h25aa, 16'h25ab, 16'h25ac, 16'h25ad, 16'h25ae, 16'h25af 	:	val_out <= 16'he629;
         16'h25b0, 16'h25b1, 16'h25b2, 16'h25b3, 16'h25b4, 16'h25b5, 16'h25b6, 16'h25b7 	:	val_out <= 16'he639;
         16'h25b8, 16'h25b9, 16'h25ba, 16'h25bb, 16'h25bc, 16'h25bd, 16'h25be, 16'h25bf 	:	val_out <= 16'he648;
         16'h25c0, 16'h25c1, 16'h25c2, 16'h25c3, 16'h25c4, 16'h25c5, 16'h25c6, 16'h25c7 	:	val_out <= 16'he657;
         16'h25c8, 16'h25c9, 16'h25ca, 16'h25cb, 16'h25cc, 16'h25cd, 16'h25ce, 16'h25cf 	:	val_out <= 16'he666;
         16'h25d0, 16'h25d1, 16'h25d2, 16'h25d3, 16'h25d4, 16'h25d5, 16'h25d6, 16'h25d7 	:	val_out <= 16'he675;
         16'h25d8, 16'h25d9, 16'h25da, 16'h25db, 16'h25dc, 16'h25dd, 16'h25de, 16'h25df 	:	val_out <= 16'he684;
         16'h25e0, 16'h25e1, 16'h25e2, 16'h25e3, 16'h25e4, 16'h25e5, 16'h25e6, 16'h25e7 	:	val_out <= 16'he693;
         16'h25e8, 16'h25e9, 16'h25ea, 16'h25eb, 16'h25ec, 16'h25ed, 16'h25ee, 16'h25ef 	:	val_out <= 16'he6a2;
         16'h25f0, 16'h25f1, 16'h25f2, 16'h25f3, 16'h25f4, 16'h25f5, 16'h25f6, 16'h25f7 	:	val_out <= 16'he6b1;
         16'h25f8, 16'h25f9, 16'h25fa, 16'h25fb, 16'h25fc, 16'h25fd, 16'h25fe, 16'h25ff 	:	val_out <= 16'he6c0;
         16'h2600, 16'h2601, 16'h2602, 16'h2603, 16'h2604, 16'h2605, 16'h2606, 16'h2607 	:	val_out <= 16'he6cf;
         16'h2608, 16'h2609, 16'h260a, 16'h260b, 16'h260c, 16'h260d, 16'h260e, 16'h260f 	:	val_out <= 16'he6de;
         16'h2610, 16'h2611, 16'h2612, 16'h2613, 16'h2614, 16'h2615, 16'h2616, 16'h2617 	:	val_out <= 16'he6ed;
         16'h2618, 16'h2619, 16'h261a, 16'h261b, 16'h261c, 16'h261d, 16'h261e, 16'h261f 	:	val_out <= 16'he6fc;
         16'h2620, 16'h2621, 16'h2622, 16'h2623, 16'h2624, 16'h2625, 16'h2626, 16'h2627 	:	val_out <= 16'he70b;
         16'h2628, 16'h2629, 16'h262a, 16'h262b, 16'h262c, 16'h262d, 16'h262e, 16'h262f 	:	val_out <= 16'he71a;
         16'h2630, 16'h2631, 16'h2632, 16'h2633, 16'h2634, 16'h2635, 16'h2636, 16'h2637 	:	val_out <= 16'he729;
         16'h2638, 16'h2639, 16'h263a, 16'h263b, 16'h263c, 16'h263d, 16'h263e, 16'h263f 	:	val_out <= 16'he737;
         16'h2640, 16'h2641, 16'h2642, 16'h2643, 16'h2644, 16'h2645, 16'h2646, 16'h2647 	:	val_out <= 16'he746;
         16'h2648, 16'h2649, 16'h264a, 16'h264b, 16'h264c, 16'h264d, 16'h264e, 16'h264f 	:	val_out <= 16'he755;
         16'h2650, 16'h2651, 16'h2652, 16'h2653, 16'h2654, 16'h2655, 16'h2656, 16'h2657 	:	val_out <= 16'he764;
         16'h2658, 16'h2659, 16'h265a, 16'h265b, 16'h265c, 16'h265d, 16'h265e, 16'h265f 	:	val_out <= 16'he773;
         16'h2660, 16'h2661, 16'h2662, 16'h2663, 16'h2664, 16'h2665, 16'h2666, 16'h2667 	:	val_out <= 16'he782;
         16'h2668, 16'h2669, 16'h266a, 16'h266b, 16'h266c, 16'h266d, 16'h266e, 16'h266f 	:	val_out <= 16'he790;
         16'h2670, 16'h2671, 16'h2672, 16'h2673, 16'h2674, 16'h2675, 16'h2676, 16'h2677 	:	val_out <= 16'he79f;
         16'h2678, 16'h2679, 16'h267a, 16'h267b, 16'h267c, 16'h267d, 16'h267e, 16'h267f 	:	val_out <= 16'he7ae;
         16'h2680, 16'h2681, 16'h2682, 16'h2683, 16'h2684, 16'h2685, 16'h2686, 16'h2687 	:	val_out <= 16'he7bd;
         16'h2688, 16'h2689, 16'h268a, 16'h268b, 16'h268c, 16'h268d, 16'h268e, 16'h268f 	:	val_out <= 16'he7cb;
         16'h2690, 16'h2691, 16'h2692, 16'h2693, 16'h2694, 16'h2695, 16'h2696, 16'h2697 	:	val_out <= 16'he7da;
         16'h2698, 16'h2699, 16'h269a, 16'h269b, 16'h269c, 16'h269d, 16'h269e, 16'h269f 	:	val_out <= 16'he7e9;
         16'h26a0, 16'h26a1, 16'h26a2, 16'h26a3, 16'h26a4, 16'h26a5, 16'h26a6, 16'h26a7 	:	val_out <= 16'he7f7;
         16'h26a8, 16'h26a9, 16'h26aa, 16'h26ab, 16'h26ac, 16'h26ad, 16'h26ae, 16'h26af 	:	val_out <= 16'he806;
         16'h26b0, 16'h26b1, 16'h26b2, 16'h26b3, 16'h26b4, 16'h26b5, 16'h26b6, 16'h26b7 	:	val_out <= 16'he815;
         16'h26b8, 16'h26b9, 16'h26ba, 16'h26bb, 16'h26bc, 16'h26bd, 16'h26be, 16'h26bf 	:	val_out <= 16'he823;
         16'h26c0, 16'h26c1, 16'h26c2, 16'h26c3, 16'h26c4, 16'h26c5, 16'h26c6, 16'h26c7 	:	val_out <= 16'he832;
         16'h26c8, 16'h26c9, 16'h26ca, 16'h26cb, 16'h26cc, 16'h26cd, 16'h26ce, 16'h26cf 	:	val_out <= 16'he840;
         16'h26d0, 16'h26d1, 16'h26d2, 16'h26d3, 16'h26d4, 16'h26d5, 16'h26d6, 16'h26d7 	:	val_out <= 16'he84f;
         16'h26d8, 16'h26d9, 16'h26da, 16'h26db, 16'h26dc, 16'h26dd, 16'h26de, 16'h26df 	:	val_out <= 16'he85e;
         16'h26e0, 16'h26e1, 16'h26e2, 16'h26e3, 16'h26e4, 16'h26e5, 16'h26e6, 16'h26e7 	:	val_out <= 16'he86c;
         16'h26e8, 16'h26e9, 16'h26ea, 16'h26eb, 16'h26ec, 16'h26ed, 16'h26ee, 16'h26ef 	:	val_out <= 16'he87b;
         16'h26f0, 16'h26f1, 16'h26f2, 16'h26f3, 16'h26f4, 16'h26f5, 16'h26f6, 16'h26f7 	:	val_out <= 16'he889;
         16'h26f8, 16'h26f9, 16'h26fa, 16'h26fb, 16'h26fc, 16'h26fd, 16'h26fe, 16'h26ff 	:	val_out <= 16'he898;
         16'h2700, 16'h2701, 16'h2702, 16'h2703, 16'h2704, 16'h2705, 16'h2706, 16'h2707 	:	val_out <= 16'he8a6;
         16'h2708, 16'h2709, 16'h270a, 16'h270b, 16'h270c, 16'h270d, 16'h270e, 16'h270f 	:	val_out <= 16'he8b5;
         16'h2710, 16'h2711, 16'h2712, 16'h2713, 16'h2714, 16'h2715, 16'h2716, 16'h2717 	:	val_out <= 16'he8c3;
         16'h2718, 16'h2719, 16'h271a, 16'h271b, 16'h271c, 16'h271d, 16'h271e, 16'h271f 	:	val_out <= 16'he8d1;
         16'h2720, 16'h2721, 16'h2722, 16'h2723, 16'h2724, 16'h2725, 16'h2726, 16'h2727 	:	val_out <= 16'he8e0;
         16'h2728, 16'h2729, 16'h272a, 16'h272b, 16'h272c, 16'h272d, 16'h272e, 16'h272f 	:	val_out <= 16'he8ee;
         16'h2730, 16'h2731, 16'h2732, 16'h2733, 16'h2734, 16'h2735, 16'h2736, 16'h2737 	:	val_out <= 16'he8fd;
         16'h2738, 16'h2739, 16'h273a, 16'h273b, 16'h273c, 16'h273d, 16'h273e, 16'h273f 	:	val_out <= 16'he90b;
         16'h2740, 16'h2741, 16'h2742, 16'h2743, 16'h2744, 16'h2745, 16'h2746, 16'h2747 	:	val_out <= 16'he919;
         16'h2748, 16'h2749, 16'h274a, 16'h274b, 16'h274c, 16'h274d, 16'h274e, 16'h274f 	:	val_out <= 16'he928;
         16'h2750, 16'h2751, 16'h2752, 16'h2753, 16'h2754, 16'h2755, 16'h2756, 16'h2757 	:	val_out <= 16'he936;
         16'h2758, 16'h2759, 16'h275a, 16'h275b, 16'h275c, 16'h275d, 16'h275e, 16'h275f 	:	val_out <= 16'he944;
         16'h2760, 16'h2761, 16'h2762, 16'h2763, 16'h2764, 16'h2765, 16'h2766, 16'h2767 	:	val_out <= 16'he953;
         16'h2768, 16'h2769, 16'h276a, 16'h276b, 16'h276c, 16'h276d, 16'h276e, 16'h276f 	:	val_out <= 16'he961;
         16'h2770, 16'h2771, 16'h2772, 16'h2773, 16'h2774, 16'h2775, 16'h2776, 16'h2777 	:	val_out <= 16'he96f;
         16'h2778, 16'h2779, 16'h277a, 16'h277b, 16'h277c, 16'h277d, 16'h277e, 16'h277f 	:	val_out <= 16'he97d;
         16'h2780, 16'h2781, 16'h2782, 16'h2783, 16'h2784, 16'h2785, 16'h2786, 16'h2787 	:	val_out <= 16'he98c;
         16'h2788, 16'h2789, 16'h278a, 16'h278b, 16'h278c, 16'h278d, 16'h278e, 16'h278f 	:	val_out <= 16'he99a;
         16'h2790, 16'h2791, 16'h2792, 16'h2793, 16'h2794, 16'h2795, 16'h2796, 16'h2797 	:	val_out <= 16'he9a8;
         16'h2798, 16'h2799, 16'h279a, 16'h279b, 16'h279c, 16'h279d, 16'h279e, 16'h279f 	:	val_out <= 16'he9b6;
         16'h27a0, 16'h27a1, 16'h27a2, 16'h27a3, 16'h27a4, 16'h27a5, 16'h27a6, 16'h27a7 	:	val_out <= 16'he9c4;
         16'h27a8, 16'h27a9, 16'h27aa, 16'h27ab, 16'h27ac, 16'h27ad, 16'h27ae, 16'h27af 	:	val_out <= 16'he9d3;
         16'h27b0, 16'h27b1, 16'h27b2, 16'h27b3, 16'h27b4, 16'h27b5, 16'h27b6, 16'h27b7 	:	val_out <= 16'he9e1;
         16'h27b8, 16'h27b9, 16'h27ba, 16'h27bb, 16'h27bc, 16'h27bd, 16'h27be, 16'h27bf 	:	val_out <= 16'he9ef;
         16'h27c0, 16'h27c1, 16'h27c2, 16'h27c3, 16'h27c4, 16'h27c5, 16'h27c6, 16'h27c7 	:	val_out <= 16'he9fd;
         16'h27c8, 16'h27c9, 16'h27ca, 16'h27cb, 16'h27cc, 16'h27cd, 16'h27ce, 16'h27cf 	:	val_out <= 16'hea0b;
         16'h27d0, 16'h27d1, 16'h27d2, 16'h27d3, 16'h27d4, 16'h27d5, 16'h27d6, 16'h27d7 	:	val_out <= 16'hea19;
         16'h27d8, 16'h27d9, 16'h27da, 16'h27db, 16'h27dc, 16'h27dd, 16'h27de, 16'h27df 	:	val_out <= 16'hea27;
         16'h27e0, 16'h27e1, 16'h27e2, 16'h27e3, 16'h27e4, 16'h27e5, 16'h27e6, 16'h27e7 	:	val_out <= 16'hea35;
         16'h27e8, 16'h27e9, 16'h27ea, 16'h27eb, 16'h27ec, 16'h27ed, 16'h27ee, 16'h27ef 	:	val_out <= 16'hea43;
         16'h27f0, 16'h27f1, 16'h27f2, 16'h27f3, 16'h27f4, 16'h27f5, 16'h27f6, 16'h27f7 	:	val_out <= 16'hea51;
         16'h27f8, 16'h27f9, 16'h27fa, 16'h27fb, 16'h27fc, 16'h27fd, 16'h27fe, 16'h27ff 	:	val_out <= 16'hea5f;
         16'h2800, 16'h2801, 16'h2802, 16'h2803, 16'h2804, 16'h2805, 16'h2806, 16'h2807 	:	val_out <= 16'hea6d;
         16'h2808, 16'h2809, 16'h280a, 16'h280b, 16'h280c, 16'h280d, 16'h280e, 16'h280f 	:	val_out <= 16'hea7b;
         16'h2810, 16'h2811, 16'h2812, 16'h2813, 16'h2814, 16'h2815, 16'h2816, 16'h2817 	:	val_out <= 16'hea89;
         16'h2818, 16'h2819, 16'h281a, 16'h281b, 16'h281c, 16'h281d, 16'h281e, 16'h281f 	:	val_out <= 16'hea97;
         16'h2820, 16'h2821, 16'h2822, 16'h2823, 16'h2824, 16'h2825, 16'h2826, 16'h2827 	:	val_out <= 16'heaa5;
         16'h2828, 16'h2829, 16'h282a, 16'h282b, 16'h282c, 16'h282d, 16'h282e, 16'h282f 	:	val_out <= 16'heab3;
         16'h2830, 16'h2831, 16'h2832, 16'h2833, 16'h2834, 16'h2835, 16'h2836, 16'h2837 	:	val_out <= 16'heac1;
         16'h2838, 16'h2839, 16'h283a, 16'h283b, 16'h283c, 16'h283d, 16'h283e, 16'h283f 	:	val_out <= 16'heace;
         16'h2840, 16'h2841, 16'h2842, 16'h2843, 16'h2844, 16'h2845, 16'h2846, 16'h2847 	:	val_out <= 16'headc;
         16'h2848, 16'h2849, 16'h284a, 16'h284b, 16'h284c, 16'h284d, 16'h284e, 16'h284f 	:	val_out <= 16'heaea;
         16'h2850, 16'h2851, 16'h2852, 16'h2853, 16'h2854, 16'h2855, 16'h2856, 16'h2857 	:	val_out <= 16'heaf8;
         16'h2858, 16'h2859, 16'h285a, 16'h285b, 16'h285c, 16'h285d, 16'h285e, 16'h285f 	:	val_out <= 16'heb06;
         16'h2860, 16'h2861, 16'h2862, 16'h2863, 16'h2864, 16'h2865, 16'h2866, 16'h2867 	:	val_out <= 16'heb13;
         16'h2868, 16'h2869, 16'h286a, 16'h286b, 16'h286c, 16'h286d, 16'h286e, 16'h286f 	:	val_out <= 16'heb21;
         16'h2870, 16'h2871, 16'h2872, 16'h2873, 16'h2874, 16'h2875, 16'h2876, 16'h2877 	:	val_out <= 16'heb2f;
         16'h2878, 16'h2879, 16'h287a, 16'h287b, 16'h287c, 16'h287d, 16'h287e, 16'h287f 	:	val_out <= 16'heb3d;
         16'h2880, 16'h2881, 16'h2882, 16'h2883, 16'h2884, 16'h2885, 16'h2886, 16'h2887 	:	val_out <= 16'heb4a;
         16'h2888, 16'h2889, 16'h288a, 16'h288b, 16'h288c, 16'h288d, 16'h288e, 16'h288f 	:	val_out <= 16'heb58;
         16'h2890, 16'h2891, 16'h2892, 16'h2893, 16'h2894, 16'h2895, 16'h2896, 16'h2897 	:	val_out <= 16'heb66;
         16'h2898, 16'h2899, 16'h289a, 16'h289b, 16'h289c, 16'h289d, 16'h289e, 16'h289f 	:	val_out <= 16'heb73;
         16'h28a0, 16'h28a1, 16'h28a2, 16'h28a3, 16'h28a4, 16'h28a5, 16'h28a6, 16'h28a7 	:	val_out <= 16'heb81;
         16'h28a8, 16'h28a9, 16'h28aa, 16'h28ab, 16'h28ac, 16'h28ad, 16'h28ae, 16'h28af 	:	val_out <= 16'heb8f;
         16'h28b0, 16'h28b1, 16'h28b2, 16'h28b3, 16'h28b4, 16'h28b5, 16'h28b6, 16'h28b7 	:	val_out <= 16'heb9c;
         16'h28b8, 16'h28b9, 16'h28ba, 16'h28bb, 16'h28bc, 16'h28bd, 16'h28be, 16'h28bf 	:	val_out <= 16'hebaa;
         16'h28c0, 16'h28c1, 16'h28c2, 16'h28c3, 16'h28c4, 16'h28c5, 16'h28c6, 16'h28c7 	:	val_out <= 16'hebb8;
         16'h28c8, 16'h28c9, 16'h28ca, 16'h28cb, 16'h28cc, 16'h28cd, 16'h28ce, 16'h28cf 	:	val_out <= 16'hebc5;
         16'h28d0, 16'h28d1, 16'h28d2, 16'h28d3, 16'h28d4, 16'h28d5, 16'h28d6, 16'h28d7 	:	val_out <= 16'hebd3;
         16'h28d8, 16'h28d9, 16'h28da, 16'h28db, 16'h28dc, 16'h28dd, 16'h28de, 16'h28df 	:	val_out <= 16'hebe0;
         16'h28e0, 16'h28e1, 16'h28e2, 16'h28e3, 16'h28e4, 16'h28e5, 16'h28e6, 16'h28e7 	:	val_out <= 16'hebee;
         16'h28e8, 16'h28e9, 16'h28ea, 16'h28eb, 16'h28ec, 16'h28ed, 16'h28ee, 16'h28ef 	:	val_out <= 16'hebfb;
         16'h28f0, 16'h28f1, 16'h28f2, 16'h28f3, 16'h28f4, 16'h28f5, 16'h28f6, 16'h28f7 	:	val_out <= 16'hec09;
         16'h28f8, 16'h28f9, 16'h28fa, 16'h28fb, 16'h28fc, 16'h28fd, 16'h28fe, 16'h28ff 	:	val_out <= 16'hec16;
         16'h2900, 16'h2901, 16'h2902, 16'h2903, 16'h2904, 16'h2905, 16'h2906, 16'h2907 	:	val_out <= 16'hec24;
         16'h2908, 16'h2909, 16'h290a, 16'h290b, 16'h290c, 16'h290d, 16'h290e, 16'h290f 	:	val_out <= 16'hec31;
         16'h2910, 16'h2911, 16'h2912, 16'h2913, 16'h2914, 16'h2915, 16'h2916, 16'h2917 	:	val_out <= 16'hec3f;
         16'h2918, 16'h2919, 16'h291a, 16'h291b, 16'h291c, 16'h291d, 16'h291e, 16'h291f 	:	val_out <= 16'hec4c;
         16'h2920, 16'h2921, 16'h2922, 16'h2923, 16'h2924, 16'h2925, 16'h2926, 16'h2927 	:	val_out <= 16'hec59;
         16'h2928, 16'h2929, 16'h292a, 16'h292b, 16'h292c, 16'h292d, 16'h292e, 16'h292f 	:	val_out <= 16'hec67;
         16'h2930, 16'h2931, 16'h2932, 16'h2933, 16'h2934, 16'h2935, 16'h2936, 16'h2937 	:	val_out <= 16'hec74;
         16'h2938, 16'h2939, 16'h293a, 16'h293b, 16'h293c, 16'h293d, 16'h293e, 16'h293f 	:	val_out <= 16'hec81;
         16'h2940, 16'h2941, 16'h2942, 16'h2943, 16'h2944, 16'h2945, 16'h2946, 16'h2947 	:	val_out <= 16'hec8f;
         16'h2948, 16'h2949, 16'h294a, 16'h294b, 16'h294c, 16'h294d, 16'h294e, 16'h294f 	:	val_out <= 16'hec9c;
         16'h2950, 16'h2951, 16'h2952, 16'h2953, 16'h2954, 16'h2955, 16'h2956, 16'h2957 	:	val_out <= 16'heca9;
         16'h2958, 16'h2959, 16'h295a, 16'h295b, 16'h295c, 16'h295d, 16'h295e, 16'h295f 	:	val_out <= 16'hecb7;
         16'h2960, 16'h2961, 16'h2962, 16'h2963, 16'h2964, 16'h2965, 16'h2966, 16'h2967 	:	val_out <= 16'hecc4;
         16'h2968, 16'h2969, 16'h296a, 16'h296b, 16'h296c, 16'h296d, 16'h296e, 16'h296f 	:	val_out <= 16'hecd1;
         16'h2970, 16'h2971, 16'h2972, 16'h2973, 16'h2974, 16'h2975, 16'h2976, 16'h2977 	:	val_out <= 16'hecde;
         16'h2978, 16'h2979, 16'h297a, 16'h297b, 16'h297c, 16'h297d, 16'h297e, 16'h297f 	:	val_out <= 16'hecec;
         16'h2980, 16'h2981, 16'h2982, 16'h2983, 16'h2984, 16'h2985, 16'h2986, 16'h2987 	:	val_out <= 16'hecf9;
         16'h2988, 16'h2989, 16'h298a, 16'h298b, 16'h298c, 16'h298d, 16'h298e, 16'h298f 	:	val_out <= 16'hed06;
         16'h2990, 16'h2991, 16'h2992, 16'h2993, 16'h2994, 16'h2995, 16'h2996, 16'h2997 	:	val_out <= 16'hed13;
         16'h2998, 16'h2999, 16'h299a, 16'h299b, 16'h299c, 16'h299d, 16'h299e, 16'h299f 	:	val_out <= 16'hed20;
         16'h29a0, 16'h29a1, 16'h29a2, 16'h29a3, 16'h29a4, 16'h29a5, 16'h29a6, 16'h29a7 	:	val_out <= 16'hed2d;
         16'h29a8, 16'h29a9, 16'h29aa, 16'h29ab, 16'h29ac, 16'h29ad, 16'h29ae, 16'h29af 	:	val_out <= 16'hed3a;
         16'h29b0, 16'h29b1, 16'h29b2, 16'h29b3, 16'h29b4, 16'h29b5, 16'h29b6, 16'h29b7 	:	val_out <= 16'hed48;
         16'h29b8, 16'h29b9, 16'h29ba, 16'h29bb, 16'h29bc, 16'h29bd, 16'h29be, 16'h29bf 	:	val_out <= 16'hed55;
         16'h29c0, 16'h29c1, 16'h29c2, 16'h29c3, 16'h29c4, 16'h29c5, 16'h29c6, 16'h29c7 	:	val_out <= 16'hed62;
         16'h29c8, 16'h29c9, 16'h29ca, 16'h29cb, 16'h29cc, 16'h29cd, 16'h29ce, 16'h29cf 	:	val_out <= 16'hed6f;
         16'h29d0, 16'h29d1, 16'h29d2, 16'h29d3, 16'h29d4, 16'h29d5, 16'h29d6, 16'h29d7 	:	val_out <= 16'hed7c;
         16'h29d8, 16'h29d9, 16'h29da, 16'h29db, 16'h29dc, 16'h29dd, 16'h29de, 16'h29df 	:	val_out <= 16'hed89;
         16'h29e0, 16'h29e1, 16'h29e2, 16'h29e3, 16'h29e4, 16'h29e5, 16'h29e6, 16'h29e7 	:	val_out <= 16'hed96;
         16'h29e8, 16'h29e9, 16'h29ea, 16'h29eb, 16'h29ec, 16'h29ed, 16'h29ee, 16'h29ef 	:	val_out <= 16'heda3;
         16'h29f0, 16'h29f1, 16'h29f2, 16'h29f3, 16'h29f4, 16'h29f5, 16'h29f6, 16'h29f7 	:	val_out <= 16'hedb0;
         16'h29f8, 16'h29f9, 16'h29fa, 16'h29fb, 16'h29fc, 16'h29fd, 16'h29fe, 16'h29ff 	:	val_out <= 16'hedbd;
         16'h2a00, 16'h2a01, 16'h2a02, 16'h2a03, 16'h2a04, 16'h2a05, 16'h2a06, 16'h2a07 	:	val_out <= 16'hedca;
         16'h2a08, 16'h2a09, 16'h2a0a, 16'h2a0b, 16'h2a0c, 16'h2a0d, 16'h2a0e, 16'h2a0f 	:	val_out <= 16'hedd6;
         16'h2a10, 16'h2a11, 16'h2a12, 16'h2a13, 16'h2a14, 16'h2a15, 16'h2a16, 16'h2a17 	:	val_out <= 16'hede3;
         16'h2a18, 16'h2a19, 16'h2a1a, 16'h2a1b, 16'h2a1c, 16'h2a1d, 16'h2a1e, 16'h2a1f 	:	val_out <= 16'hedf0;
         16'h2a20, 16'h2a21, 16'h2a22, 16'h2a23, 16'h2a24, 16'h2a25, 16'h2a26, 16'h2a27 	:	val_out <= 16'hedfd;
         16'h2a28, 16'h2a29, 16'h2a2a, 16'h2a2b, 16'h2a2c, 16'h2a2d, 16'h2a2e, 16'h2a2f 	:	val_out <= 16'hee0a;
         16'h2a30, 16'h2a31, 16'h2a32, 16'h2a33, 16'h2a34, 16'h2a35, 16'h2a36, 16'h2a37 	:	val_out <= 16'hee17;
         16'h2a38, 16'h2a39, 16'h2a3a, 16'h2a3b, 16'h2a3c, 16'h2a3d, 16'h2a3e, 16'h2a3f 	:	val_out <= 16'hee24;
         16'h2a40, 16'h2a41, 16'h2a42, 16'h2a43, 16'h2a44, 16'h2a45, 16'h2a46, 16'h2a47 	:	val_out <= 16'hee30;
         16'h2a48, 16'h2a49, 16'h2a4a, 16'h2a4b, 16'h2a4c, 16'h2a4d, 16'h2a4e, 16'h2a4f 	:	val_out <= 16'hee3d;
         16'h2a50, 16'h2a51, 16'h2a52, 16'h2a53, 16'h2a54, 16'h2a55, 16'h2a56, 16'h2a57 	:	val_out <= 16'hee4a;
         16'h2a58, 16'h2a59, 16'h2a5a, 16'h2a5b, 16'h2a5c, 16'h2a5d, 16'h2a5e, 16'h2a5f 	:	val_out <= 16'hee57;
         16'h2a60, 16'h2a61, 16'h2a62, 16'h2a63, 16'h2a64, 16'h2a65, 16'h2a66, 16'h2a67 	:	val_out <= 16'hee63;
         16'h2a68, 16'h2a69, 16'h2a6a, 16'h2a6b, 16'h2a6c, 16'h2a6d, 16'h2a6e, 16'h2a6f 	:	val_out <= 16'hee70;
         16'h2a70, 16'h2a71, 16'h2a72, 16'h2a73, 16'h2a74, 16'h2a75, 16'h2a76, 16'h2a77 	:	val_out <= 16'hee7d;
         16'h2a78, 16'h2a79, 16'h2a7a, 16'h2a7b, 16'h2a7c, 16'h2a7d, 16'h2a7e, 16'h2a7f 	:	val_out <= 16'hee89;
         16'h2a80, 16'h2a81, 16'h2a82, 16'h2a83, 16'h2a84, 16'h2a85, 16'h2a86, 16'h2a87 	:	val_out <= 16'hee96;
         16'h2a88, 16'h2a89, 16'h2a8a, 16'h2a8b, 16'h2a8c, 16'h2a8d, 16'h2a8e, 16'h2a8f 	:	val_out <= 16'heea3;
         16'h2a90, 16'h2a91, 16'h2a92, 16'h2a93, 16'h2a94, 16'h2a95, 16'h2a96, 16'h2a97 	:	val_out <= 16'heeaf;
         16'h2a98, 16'h2a99, 16'h2a9a, 16'h2a9b, 16'h2a9c, 16'h2a9d, 16'h2a9e, 16'h2a9f 	:	val_out <= 16'heebc;
         16'h2aa0, 16'h2aa1, 16'h2aa2, 16'h2aa3, 16'h2aa4, 16'h2aa5, 16'h2aa6, 16'h2aa7 	:	val_out <= 16'heec9;
         16'h2aa8, 16'h2aa9, 16'h2aaa, 16'h2aab, 16'h2aac, 16'h2aad, 16'h2aae, 16'h2aaf 	:	val_out <= 16'heed5;
         16'h2ab0, 16'h2ab1, 16'h2ab2, 16'h2ab3, 16'h2ab4, 16'h2ab5, 16'h2ab6, 16'h2ab7 	:	val_out <= 16'heee2;
         16'h2ab8, 16'h2ab9, 16'h2aba, 16'h2abb, 16'h2abc, 16'h2abd, 16'h2abe, 16'h2abf 	:	val_out <= 16'heeee;
         16'h2ac0, 16'h2ac1, 16'h2ac2, 16'h2ac3, 16'h2ac4, 16'h2ac5, 16'h2ac6, 16'h2ac7 	:	val_out <= 16'heefb;
         16'h2ac8, 16'h2ac9, 16'h2aca, 16'h2acb, 16'h2acc, 16'h2acd, 16'h2ace, 16'h2acf 	:	val_out <= 16'hef07;
         16'h2ad0, 16'h2ad1, 16'h2ad2, 16'h2ad3, 16'h2ad4, 16'h2ad5, 16'h2ad6, 16'h2ad7 	:	val_out <= 16'hef14;
         16'h2ad8, 16'h2ad9, 16'h2ada, 16'h2adb, 16'h2adc, 16'h2add, 16'h2ade, 16'h2adf 	:	val_out <= 16'hef20;
         16'h2ae0, 16'h2ae1, 16'h2ae2, 16'h2ae3, 16'h2ae4, 16'h2ae5, 16'h2ae6, 16'h2ae7 	:	val_out <= 16'hef2d;
         16'h2ae8, 16'h2ae9, 16'h2aea, 16'h2aeb, 16'h2aec, 16'h2aed, 16'h2aee, 16'h2aef 	:	val_out <= 16'hef39;
         16'h2af0, 16'h2af1, 16'h2af2, 16'h2af3, 16'h2af4, 16'h2af5, 16'h2af6, 16'h2af7 	:	val_out <= 16'hef46;
         16'h2af8, 16'h2af9, 16'h2afa, 16'h2afb, 16'h2afc, 16'h2afd, 16'h2afe, 16'h2aff 	:	val_out <= 16'hef52;
         16'h2b00, 16'h2b01, 16'h2b02, 16'h2b03, 16'h2b04, 16'h2b05, 16'h2b06, 16'h2b07 	:	val_out <= 16'hef5f;
         16'h2b08, 16'h2b09, 16'h2b0a, 16'h2b0b, 16'h2b0c, 16'h2b0d, 16'h2b0e, 16'h2b0f 	:	val_out <= 16'hef6b;
         16'h2b10, 16'h2b11, 16'h2b12, 16'h2b13, 16'h2b14, 16'h2b15, 16'h2b16, 16'h2b17 	:	val_out <= 16'hef77;
         16'h2b18, 16'h2b19, 16'h2b1a, 16'h2b1b, 16'h2b1c, 16'h2b1d, 16'h2b1e, 16'h2b1f 	:	val_out <= 16'hef84;
         16'h2b20, 16'h2b21, 16'h2b22, 16'h2b23, 16'h2b24, 16'h2b25, 16'h2b26, 16'h2b27 	:	val_out <= 16'hef90;
         16'h2b28, 16'h2b29, 16'h2b2a, 16'h2b2b, 16'h2b2c, 16'h2b2d, 16'h2b2e, 16'h2b2f 	:	val_out <= 16'hef9c;
         16'h2b30, 16'h2b31, 16'h2b32, 16'h2b33, 16'h2b34, 16'h2b35, 16'h2b36, 16'h2b37 	:	val_out <= 16'hefa9;
         16'h2b38, 16'h2b39, 16'h2b3a, 16'h2b3b, 16'h2b3c, 16'h2b3d, 16'h2b3e, 16'h2b3f 	:	val_out <= 16'hefb5;
         16'h2b40, 16'h2b41, 16'h2b42, 16'h2b43, 16'h2b44, 16'h2b45, 16'h2b46, 16'h2b47 	:	val_out <= 16'hefc1;
         16'h2b48, 16'h2b49, 16'h2b4a, 16'h2b4b, 16'h2b4c, 16'h2b4d, 16'h2b4e, 16'h2b4f 	:	val_out <= 16'hefcd;
         16'h2b50, 16'h2b51, 16'h2b52, 16'h2b53, 16'h2b54, 16'h2b55, 16'h2b56, 16'h2b57 	:	val_out <= 16'hefda;
         16'h2b58, 16'h2b59, 16'h2b5a, 16'h2b5b, 16'h2b5c, 16'h2b5d, 16'h2b5e, 16'h2b5f 	:	val_out <= 16'hefe6;
         16'h2b60, 16'h2b61, 16'h2b62, 16'h2b63, 16'h2b64, 16'h2b65, 16'h2b66, 16'h2b67 	:	val_out <= 16'heff2;
         16'h2b68, 16'h2b69, 16'h2b6a, 16'h2b6b, 16'h2b6c, 16'h2b6d, 16'h2b6e, 16'h2b6f 	:	val_out <= 16'heffe;
         16'h2b70, 16'h2b71, 16'h2b72, 16'h2b73, 16'h2b74, 16'h2b75, 16'h2b76, 16'h2b77 	:	val_out <= 16'hf00a;
         16'h2b78, 16'h2b79, 16'h2b7a, 16'h2b7b, 16'h2b7c, 16'h2b7d, 16'h2b7e, 16'h2b7f 	:	val_out <= 16'hf016;
         16'h2b80, 16'h2b81, 16'h2b82, 16'h2b83, 16'h2b84, 16'h2b85, 16'h2b86, 16'h2b87 	:	val_out <= 16'hf023;
         16'h2b88, 16'h2b89, 16'h2b8a, 16'h2b8b, 16'h2b8c, 16'h2b8d, 16'h2b8e, 16'h2b8f 	:	val_out <= 16'hf02f;
         16'h2b90, 16'h2b91, 16'h2b92, 16'h2b93, 16'h2b94, 16'h2b95, 16'h2b96, 16'h2b97 	:	val_out <= 16'hf03b;
         16'h2b98, 16'h2b99, 16'h2b9a, 16'h2b9b, 16'h2b9c, 16'h2b9d, 16'h2b9e, 16'h2b9f 	:	val_out <= 16'hf047;
         16'h2ba0, 16'h2ba1, 16'h2ba2, 16'h2ba3, 16'h2ba4, 16'h2ba5, 16'h2ba6, 16'h2ba7 	:	val_out <= 16'hf053;
         16'h2ba8, 16'h2ba9, 16'h2baa, 16'h2bab, 16'h2bac, 16'h2bad, 16'h2bae, 16'h2baf 	:	val_out <= 16'hf05f;
         16'h2bb0, 16'h2bb1, 16'h2bb2, 16'h2bb3, 16'h2bb4, 16'h2bb5, 16'h2bb6, 16'h2bb7 	:	val_out <= 16'hf06b;
         16'h2bb8, 16'h2bb9, 16'h2bba, 16'h2bbb, 16'h2bbc, 16'h2bbd, 16'h2bbe, 16'h2bbf 	:	val_out <= 16'hf077;
         16'h2bc0, 16'h2bc1, 16'h2bc2, 16'h2bc3, 16'h2bc4, 16'h2bc5, 16'h2bc6, 16'h2bc7 	:	val_out <= 16'hf083;
         16'h2bc8, 16'h2bc9, 16'h2bca, 16'h2bcb, 16'h2bcc, 16'h2bcd, 16'h2bce, 16'h2bcf 	:	val_out <= 16'hf08f;
         16'h2bd0, 16'h2bd1, 16'h2bd2, 16'h2bd3, 16'h2bd4, 16'h2bd5, 16'h2bd6, 16'h2bd7 	:	val_out <= 16'hf09b;
         16'h2bd8, 16'h2bd9, 16'h2bda, 16'h2bdb, 16'h2bdc, 16'h2bdd, 16'h2bde, 16'h2bdf 	:	val_out <= 16'hf0a7;
         16'h2be0, 16'h2be1, 16'h2be2, 16'h2be3, 16'h2be4, 16'h2be5, 16'h2be6, 16'h2be7 	:	val_out <= 16'hf0b3;
         16'h2be8, 16'h2be9, 16'h2bea, 16'h2beb, 16'h2bec, 16'h2bed, 16'h2bee, 16'h2bef 	:	val_out <= 16'hf0bf;
         16'h2bf0, 16'h2bf1, 16'h2bf2, 16'h2bf3, 16'h2bf4, 16'h2bf5, 16'h2bf6, 16'h2bf7 	:	val_out <= 16'hf0cb;
         16'h2bf8, 16'h2bf9, 16'h2bfa, 16'h2bfb, 16'h2bfc, 16'h2bfd, 16'h2bfe, 16'h2bff 	:	val_out <= 16'hf0d6;
         16'h2c00, 16'h2c01, 16'h2c02, 16'h2c03, 16'h2c04, 16'h2c05, 16'h2c06, 16'h2c07 	:	val_out <= 16'hf0e2;
         16'h2c08, 16'h2c09, 16'h2c0a, 16'h2c0b, 16'h2c0c, 16'h2c0d, 16'h2c0e, 16'h2c0f 	:	val_out <= 16'hf0ee;
         16'h2c10, 16'h2c11, 16'h2c12, 16'h2c13, 16'h2c14, 16'h2c15, 16'h2c16, 16'h2c17 	:	val_out <= 16'hf0fa;
         16'h2c18, 16'h2c19, 16'h2c1a, 16'h2c1b, 16'h2c1c, 16'h2c1d, 16'h2c1e, 16'h2c1f 	:	val_out <= 16'hf106;
         16'h2c20, 16'h2c21, 16'h2c22, 16'h2c23, 16'h2c24, 16'h2c25, 16'h2c26, 16'h2c27 	:	val_out <= 16'hf112;
         16'h2c28, 16'h2c29, 16'h2c2a, 16'h2c2b, 16'h2c2c, 16'h2c2d, 16'h2c2e, 16'h2c2f 	:	val_out <= 16'hf11d;
         16'h2c30, 16'h2c31, 16'h2c32, 16'h2c33, 16'h2c34, 16'h2c35, 16'h2c36, 16'h2c37 	:	val_out <= 16'hf129;
         16'h2c38, 16'h2c39, 16'h2c3a, 16'h2c3b, 16'h2c3c, 16'h2c3d, 16'h2c3e, 16'h2c3f 	:	val_out <= 16'hf135;
         16'h2c40, 16'h2c41, 16'h2c42, 16'h2c43, 16'h2c44, 16'h2c45, 16'h2c46, 16'h2c47 	:	val_out <= 16'hf141;
         16'h2c48, 16'h2c49, 16'h2c4a, 16'h2c4b, 16'h2c4c, 16'h2c4d, 16'h2c4e, 16'h2c4f 	:	val_out <= 16'hf14c;
         16'h2c50, 16'h2c51, 16'h2c52, 16'h2c53, 16'h2c54, 16'h2c55, 16'h2c56, 16'h2c57 	:	val_out <= 16'hf158;
         16'h2c58, 16'h2c59, 16'h2c5a, 16'h2c5b, 16'h2c5c, 16'h2c5d, 16'h2c5e, 16'h2c5f 	:	val_out <= 16'hf164;
         16'h2c60, 16'h2c61, 16'h2c62, 16'h2c63, 16'h2c64, 16'h2c65, 16'h2c66, 16'h2c67 	:	val_out <= 16'hf16f;
         16'h2c68, 16'h2c69, 16'h2c6a, 16'h2c6b, 16'h2c6c, 16'h2c6d, 16'h2c6e, 16'h2c6f 	:	val_out <= 16'hf17b;
         16'h2c70, 16'h2c71, 16'h2c72, 16'h2c73, 16'h2c74, 16'h2c75, 16'h2c76, 16'h2c77 	:	val_out <= 16'hf186;
         16'h2c78, 16'h2c79, 16'h2c7a, 16'h2c7b, 16'h2c7c, 16'h2c7d, 16'h2c7e, 16'h2c7f 	:	val_out <= 16'hf192;
         16'h2c80, 16'h2c81, 16'h2c82, 16'h2c83, 16'h2c84, 16'h2c85, 16'h2c86, 16'h2c87 	:	val_out <= 16'hf19e;
         16'h2c88, 16'h2c89, 16'h2c8a, 16'h2c8b, 16'h2c8c, 16'h2c8d, 16'h2c8e, 16'h2c8f 	:	val_out <= 16'hf1a9;
         16'h2c90, 16'h2c91, 16'h2c92, 16'h2c93, 16'h2c94, 16'h2c95, 16'h2c96, 16'h2c97 	:	val_out <= 16'hf1b5;
         16'h2c98, 16'h2c99, 16'h2c9a, 16'h2c9b, 16'h2c9c, 16'h2c9d, 16'h2c9e, 16'h2c9f 	:	val_out <= 16'hf1c0;
         16'h2ca0, 16'h2ca1, 16'h2ca2, 16'h2ca3, 16'h2ca4, 16'h2ca5, 16'h2ca6, 16'h2ca7 	:	val_out <= 16'hf1cc;
         16'h2ca8, 16'h2ca9, 16'h2caa, 16'h2cab, 16'h2cac, 16'h2cad, 16'h2cae, 16'h2caf 	:	val_out <= 16'hf1d7;
         16'h2cb0, 16'h2cb1, 16'h2cb2, 16'h2cb3, 16'h2cb4, 16'h2cb5, 16'h2cb6, 16'h2cb7 	:	val_out <= 16'hf1e3;
         16'h2cb8, 16'h2cb9, 16'h2cba, 16'h2cbb, 16'h2cbc, 16'h2cbd, 16'h2cbe, 16'h2cbf 	:	val_out <= 16'hf1ee;
         16'h2cc0, 16'h2cc1, 16'h2cc2, 16'h2cc3, 16'h2cc4, 16'h2cc5, 16'h2cc6, 16'h2cc7 	:	val_out <= 16'hf1fa;
         16'h2cc8, 16'h2cc9, 16'h2cca, 16'h2ccb, 16'h2ccc, 16'h2ccd, 16'h2cce, 16'h2ccf 	:	val_out <= 16'hf205;
         16'h2cd0, 16'h2cd1, 16'h2cd2, 16'h2cd3, 16'h2cd4, 16'h2cd5, 16'h2cd6, 16'h2cd7 	:	val_out <= 16'hf211;
         16'h2cd8, 16'h2cd9, 16'h2cda, 16'h2cdb, 16'h2cdc, 16'h2cdd, 16'h2cde, 16'h2cdf 	:	val_out <= 16'hf21c;
         16'h2ce0, 16'h2ce1, 16'h2ce2, 16'h2ce3, 16'h2ce4, 16'h2ce5, 16'h2ce6, 16'h2ce7 	:	val_out <= 16'hf227;
         16'h2ce8, 16'h2ce9, 16'h2cea, 16'h2ceb, 16'h2cec, 16'h2ced, 16'h2cee, 16'h2cef 	:	val_out <= 16'hf233;
         16'h2cf0, 16'h2cf1, 16'h2cf2, 16'h2cf3, 16'h2cf4, 16'h2cf5, 16'h2cf6, 16'h2cf7 	:	val_out <= 16'hf23e;
         16'h2cf8, 16'h2cf9, 16'h2cfa, 16'h2cfb, 16'h2cfc, 16'h2cfd, 16'h2cfe, 16'h2cff 	:	val_out <= 16'hf249;
         16'h2d00, 16'h2d01, 16'h2d02, 16'h2d03, 16'h2d04, 16'h2d05, 16'h2d06, 16'h2d07 	:	val_out <= 16'hf255;
         16'h2d08, 16'h2d09, 16'h2d0a, 16'h2d0b, 16'h2d0c, 16'h2d0d, 16'h2d0e, 16'h2d0f 	:	val_out <= 16'hf260;
         16'h2d10, 16'h2d11, 16'h2d12, 16'h2d13, 16'h2d14, 16'h2d15, 16'h2d16, 16'h2d17 	:	val_out <= 16'hf26b;
         16'h2d18, 16'h2d19, 16'h2d1a, 16'h2d1b, 16'h2d1c, 16'h2d1d, 16'h2d1e, 16'h2d1f 	:	val_out <= 16'hf276;
         16'h2d20, 16'h2d21, 16'h2d22, 16'h2d23, 16'h2d24, 16'h2d25, 16'h2d26, 16'h2d27 	:	val_out <= 16'hf282;
         16'h2d28, 16'h2d29, 16'h2d2a, 16'h2d2b, 16'h2d2c, 16'h2d2d, 16'h2d2e, 16'h2d2f 	:	val_out <= 16'hf28d;
         16'h2d30, 16'h2d31, 16'h2d32, 16'h2d33, 16'h2d34, 16'h2d35, 16'h2d36, 16'h2d37 	:	val_out <= 16'hf298;
         16'h2d38, 16'h2d39, 16'h2d3a, 16'h2d3b, 16'h2d3c, 16'h2d3d, 16'h2d3e, 16'h2d3f 	:	val_out <= 16'hf2a3;
         16'h2d40, 16'h2d41, 16'h2d42, 16'h2d43, 16'h2d44, 16'h2d45, 16'h2d46, 16'h2d47 	:	val_out <= 16'hf2af;
         16'h2d48, 16'h2d49, 16'h2d4a, 16'h2d4b, 16'h2d4c, 16'h2d4d, 16'h2d4e, 16'h2d4f 	:	val_out <= 16'hf2ba;
         16'h2d50, 16'h2d51, 16'h2d52, 16'h2d53, 16'h2d54, 16'h2d55, 16'h2d56, 16'h2d57 	:	val_out <= 16'hf2c5;
         16'h2d58, 16'h2d59, 16'h2d5a, 16'h2d5b, 16'h2d5c, 16'h2d5d, 16'h2d5e, 16'h2d5f 	:	val_out <= 16'hf2d0;
         16'h2d60, 16'h2d61, 16'h2d62, 16'h2d63, 16'h2d64, 16'h2d65, 16'h2d66, 16'h2d67 	:	val_out <= 16'hf2db;
         16'h2d68, 16'h2d69, 16'h2d6a, 16'h2d6b, 16'h2d6c, 16'h2d6d, 16'h2d6e, 16'h2d6f 	:	val_out <= 16'hf2e6;
         16'h2d70, 16'h2d71, 16'h2d72, 16'h2d73, 16'h2d74, 16'h2d75, 16'h2d76, 16'h2d77 	:	val_out <= 16'hf2f1;
         16'h2d78, 16'h2d79, 16'h2d7a, 16'h2d7b, 16'h2d7c, 16'h2d7d, 16'h2d7e, 16'h2d7f 	:	val_out <= 16'hf2fc;
         16'h2d80, 16'h2d81, 16'h2d82, 16'h2d83, 16'h2d84, 16'h2d85, 16'h2d86, 16'h2d87 	:	val_out <= 16'hf307;
         16'h2d88, 16'h2d89, 16'h2d8a, 16'h2d8b, 16'h2d8c, 16'h2d8d, 16'h2d8e, 16'h2d8f 	:	val_out <= 16'hf312;
         16'h2d90, 16'h2d91, 16'h2d92, 16'h2d93, 16'h2d94, 16'h2d95, 16'h2d96, 16'h2d97 	:	val_out <= 16'hf31d;
         16'h2d98, 16'h2d99, 16'h2d9a, 16'h2d9b, 16'h2d9c, 16'h2d9d, 16'h2d9e, 16'h2d9f 	:	val_out <= 16'hf328;
         16'h2da0, 16'h2da1, 16'h2da2, 16'h2da3, 16'h2da4, 16'h2da5, 16'h2da6, 16'h2da7 	:	val_out <= 16'hf333;
         16'h2da8, 16'h2da9, 16'h2daa, 16'h2dab, 16'h2dac, 16'h2dad, 16'h2dae, 16'h2daf 	:	val_out <= 16'hf33e;
         16'h2db0, 16'h2db1, 16'h2db2, 16'h2db3, 16'h2db4, 16'h2db5, 16'h2db6, 16'h2db7 	:	val_out <= 16'hf349;
         16'h2db8, 16'h2db9, 16'h2dba, 16'h2dbb, 16'h2dbc, 16'h2dbd, 16'h2dbe, 16'h2dbf 	:	val_out <= 16'hf354;
         16'h2dc0, 16'h2dc1, 16'h2dc2, 16'h2dc3, 16'h2dc4, 16'h2dc5, 16'h2dc6, 16'h2dc7 	:	val_out <= 16'hf35f;
         16'h2dc8, 16'h2dc9, 16'h2dca, 16'h2dcb, 16'h2dcc, 16'h2dcd, 16'h2dce, 16'h2dcf 	:	val_out <= 16'hf36a;
         16'h2dd0, 16'h2dd1, 16'h2dd2, 16'h2dd3, 16'h2dd4, 16'h2dd5, 16'h2dd6, 16'h2dd7 	:	val_out <= 16'hf375;
         16'h2dd8, 16'h2dd9, 16'h2dda, 16'h2ddb, 16'h2ddc, 16'h2ddd, 16'h2dde, 16'h2ddf 	:	val_out <= 16'hf37f;
         16'h2de0, 16'h2de1, 16'h2de2, 16'h2de3, 16'h2de4, 16'h2de5, 16'h2de6, 16'h2de7 	:	val_out <= 16'hf38a;
         16'h2de8, 16'h2de9, 16'h2dea, 16'h2deb, 16'h2dec, 16'h2ded, 16'h2dee, 16'h2def 	:	val_out <= 16'hf395;
         16'h2df0, 16'h2df1, 16'h2df2, 16'h2df3, 16'h2df4, 16'h2df5, 16'h2df6, 16'h2df7 	:	val_out <= 16'hf3a0;
         16'h2df8, 16'h2df9, 16'h2dfa, 16'h2dfb, 16'h2dfc, 16'h2dfd, 16'h2dfe, 16'h2dff 	:	val_out <= 16'hf3ab;
         16'h2e00, 16'h2e01, 16'h2e02, 16'h2e03, 16'h2e04, 16'h2e05, 16'h2e06, 16'h2e07 	:	val_out <= 16'hf3b5;
         16'h2e08, 16'h2e09, 16'h2e0a, 16'h2e0b, 16'h2e0c, 16'h2e0d, 16'h2e0e, 16'h2e0f 	:	val_out <= 16'hf3c0;
         16'h2e10, 16'h2e11, 16'h2e12, 16'h2e13, 16'h2e14, 16'h2e15, 16'h2e16, 16'h2e17 	:	val_out <= 16'hf3cb;
         16'h2e18, 16'h2e19, 16'h2e1a, 16'h2e1b, 16'h2e1c, 16'h2e1d, 16'h2e1e, 16'h2e1f 	:	val_out <= 16'hf3d6;
         16'h2e20, 16'h2e21, 16'h2e22, 16'h2e23, 16'h2e24, 16'h2e25, 16'h2e26, 16'h2e27 	:	val_out <= 16'hf3e0;
         16'h2e28, 16'h2e29, 16'h2e2a, 16'h2e2b, 16'h2e2c, 16'h2e2d, 16'h2e2e, 16'h2e2f 	:	val_out <= 16'hf3eb;
         16'h2e30, 16'h2e31, 16'h2e32, 16'h2e33, 16'h2e34, 16'h2e35, 16'h2e36, 16'h2e37 	:	val_out <= 16'hf3f6;
         16'h2e38, 16'h2e39, 16'h2e3a, 16'h2e3b, 16'h2e3c, 16'h2e3d, 16'h2e3e, 16'h2e3f 	:	val_out <= 16'hf400;
         16'h2e40, 16'h2e41, 16'h2e42, 16'h2e43, 16'h2e44, 16'h2e45, 16'h2e46, 16'h2e47 	:	val_out <= 16'hf40b;
         16'h2e48, 16'h2e49, 16'h2e4a, 16'h2e4b, 16'h2e4c, 16'h2e4d, 16'h2e4e, 16'h2e4f 	:	val_out <= 16'hf415;
         16'h2e50, 16'h2e51, 16'h2e52, 16'h2e53, 16'h2e54, 16'h2e55, 16'h2e56, 16'h2e57 	:	val_out <= 16'hf420;
         16'h2e58, 16'h2e59, 16'h2e5a, 16'h2e5b, 16'h2e5c, 16'h2e5d, 16'h2e5e, 16'h2e5f 	:	val_out <= 16'hf42b;
         16'h2e60, 16'h2e61, 16'h2e62, 16'h2e63, 16'h2e64, 16'h2e65, 16'h2e66, 16'h2e67 	:	val_out <= 16'hf435;
         16'h2e68, 16'h2e69, 16'h2e6a, 16'h2e6b, 16'h2e6c, 16'h2e6d, 16'h2e6e, 16'h2e6f 	:	val_out <= 16'hf440;
         16'h2e70, 16'h2e71, 16'h2e72, 16'h2e73, 16'h2e74, 16'h2e75, 16'h2e76, 16'h2e77 	:	val_out <= 16'hf44a;
         16'h2e78, 16'h2e79, 16'h2e7a, 16'h2e7b, 16'h2e7c, 16'h2e7d, 16'h2e7e, 16'h2e7f 	:	val_out <= 16'hf455;
         16'h2e80, 16'h2e81, 16'h2e82, 16'h2e83, 16'h2e84, 16'h2e85, 16'h2e86, 16'h2e87 	:	val_out <= 16'hf45f;
         16'h2e88, 16'h2e89, 16'h2e8a, 16'h2e8b, 16'h2e8c, 16'h2e8d, 16'h2e8e, 16'h2e8f 	:	val_out <= 16'hf46a;
         16'h2e90, 16'h2e91, 16'h2e92, 16'h2e93, 16'h2e94, 16'h2e95, 16'h2e96, 16'h2e97 	:	val_out <= 16'hf474;
         16'h2e98, 16'h2e99, 16'h2e9a, 16'h2e9b, 16'h2e9c, 16'h2e9d, 16'h2e9e, 16'h2e9f 	:	val_out <= 16'hf47e;
         16'h2ea0, 16'h2ea1, 16'h2ea2, 16'h2ea3, 16'h2ea4, 16'h2ea5, 16'h2ea6, 16'h2ea7 	:	val_out <= 16'hf489;
         16'h2ea8, 16'h2ea9, 16'h2eaa, 16'h2eab, 16'h2eac, 16'h2ead, 16'h2eae, 16'h2eaf 	:	val_out <= 16'hf493;
         16'h2eb0, 16'h2eb1, 16'h2eb2, 16'h2eb3, 16'h2eb4, 16'h2eb5, 16'h2eb6, 16'h2eb7 	:	val_out <= 16'hf49e;
         16'h2eb8, 16'h2eb9, 16'h2eba, 16'h2ebb, 16'h2ebc, 16'h2ebd, 16'h2ebe, 16'h2ebf 	:	val_out <= 16'hf4a8;
         16'h2ec0, 16'h2ec1, 16'h2ec2, 16'h2ec3, 16'h2ec4, 16'h2ec5, 16'h2ec6, 16'h2ec7 	:	val_out <= 16'hf4b2;
         16'h2ec8, 16'h2ec9, 16'h2eca, 16'h2ecb, 16'h2ecc, 16'h2ecd, 16'h2ece, 16'h2ecf 	:	val_out <= 16'hf4bd;
         16'h2ed0, 16'h2ed1, 16'h2ed2, 16'h2ed3, 16'h2ed4, 16'h2ed5, 16'h2ed6, 16'h2ed7 	:	val_out <= 16'hf4c7;
         16'h2ed8, 16'h2ed9, 16'h2eda, 16'h2edb, 16'h2edc, 16'h2edd, 16'h2ede, 16'h2edf 	:	val_out <= 16'hf4d1;
         16'h2ee0, 16'h2ee1, 16'h2ee2, 16'h2ee3, 16'h2ee4, 16'h2ee5, 16'h2ee6, 16'h2ee7 	:	val_out <= 16'hf4db;
         16'h2ee8, 16'h2ee9, 16'h2eea, 16'h2eeb, 16'h2eec, 16'h2eed, 16'h2eee, 16'h2eef 	:	val_out <= 16'hf4e6;
         16'h2ef0, 16'h2ef1, 16'h2ef2, 16'h2ef3, 16'h2ef4, 16'h2ef5, 16'h2ef6, 16'h2ef7 	:	val_out <= 16'hf4f0;
         16'h2ef8, 16'h2ef9, 16'h2efa, 16'h2efb, 16'h2efc, 16'h2efd, 16'h2efe, 16'h2eff 	:	val_out <= 16'hf4fa;
         16'h2f00, 16'h2f01, 16'h2f02, 16'h2f03, 16'h2f04, 16'h2f05, 16'h2f06, 16'h2f07 	:	val_out <= 16'hf504;
         16'h2f08, 16'h2f09, 16'h2f0a, 16'h2f0b, 16'h2f0c, 16'h2f0d, 16'h2f0e, 16'h2f0f 	:	val_out <= 16'hf50f;
         16'h2f10, 16'h2f11, 16'h2f12, 16'h2f13, 16'h2f14, 16'h2f15, 16'h2f16, 16'h2f17 	:	val_out <= 16'hf519;
         16'h2f18, 16'h2f19, 16'h2f1a, 16'h2f1b, 16'h2f1c, 16'h2f1d, 16'h2f1e, 16'h2f1f 	:	val_out <= 16'hf523;
         16'h2f20, 16'h2f21, 16'h2f22, 16'h2f23, 16'h2f24, 16'h2f25, 16'h2f26, 16'h2f27 	:	val_out <= 16'hf52d;
         16'h2f28, 16'h2f29, 16'h2f2a, 16'h2f2b, 16'h2f2c, 16'h2f2d, 16'h2f2e, 16'h2f2f 	:	val_out <= 16'hf537;
         16'h2f30, 16'h2f31, 16'h2f32, 16'h2f33, 16'h2f34, 16'h2f35, 16'h2f36, 16'h2f37 	:	val_out <= 16'hf541;
         16'h2f38, 16'h2f39, 16'h2f3a, 16'h2f3b, 16'h2f3c, 16'h2f3d, 16'h2f3e, 16'h2f3f 	:	val_out <= 16'hf54b;
         16'h2f40, 16'h2f41, 16'h2f42, 16'h2f43, 16'h2f44, 16'h2f45, 16'h2f46, 16'h2f47 	:	val_out <= 16'hf555;
         16'h2f48, 16'h2f49, 16'h2f4a, 16'h2f4b, 16'h2f4c, 16'h2f4d, 16'h2f4e, 16'h2f4f 	:	val_out <= 16'hf55f;
         16'h2f50, 16'h2f51, 16'h2f52, 16'h2f53, 16'h2f54, 16'h2f55, 16'h2f56, 16'h2f57 	:	val_out <= 16'hf569;
         16'h2f58, 16'h2f59, 16'h2f5a, 16'h2f5b, 16'h2f5c, 16'h2f5d, 16'h2f5e, 16'h2f5f 	:	val_out <= 16'hf573;
         16'h2f60, 16'h2f61, 16'h2f62, 16'h2f63, 16'h2f64, 16'h2f65, 16'h2f66, 16'h2f67 	:	val_out <= 16'hf57d;
         16'h2f68, 16'h2f69, 16'h2f6a, 16'h2f6b, 16'h2f6c, 16'h2f6d, 16'h2f6e, 16'h2f6f 	:	val_out <= 16'hf587;
         16'h2f70, 16'h2f71, 16'h2f72, 16'h2f73, 16'h2f74, 16'h2f75, 16'h2f76, 16'h2f77 	:	val_out <= 16'hf591;
         16'h2f78, 16'h2f79, 16'h2f7a, 16'h2f7b, 16'h2f7c, 16'h2f7d, 16'h2f7e, 16'h2f7f 	:	val_out <= 16'hf59b;
         16'h2f80, 16'h2f81, 16'h2f82, 16'h2f83, 16'h2f84, 16'h2f85, 16'h2f86, 16'h2f87 	:	val_out <= 16'hf5a5;
         16'h2f88, 16'h2f89, 16'h2f8a, 16'h2f8b, 16'h2f8c, 16'h2f8d, 16'h2f8e, 16'h2f8f 	:	val_out <= 16'hf5af;
         16'h2f90, 16'h2f91, 16'h2f92, 16'h2f93, 16'h2f94, 16'h2f95, 16'h2f96, 16'h2f97 	:	val_out <= 16'hf5b9;
         16'h2f98, 16'h2f99, 16'h2f9a, 16'h2f9b, 16'h2f9c, 16'h2f9d, 16'h2f9e, 16'h2f9f 	:	val_out <= 16'hf5c3;
         16'h2fa0, 16'h2fa1, 16'h2fa2, 16'h2fa3, 16'h2fa4, 16'h2fa5, 16'h2fa6, 16'h2fa7 	:	val_out <= 16'hf5cc;
         16'h2fa8, 16'h2fa9, 16'h2faa, 16'h2fab, 16'h2fac, 16'h2fad, 16'h2fae, 16'h2faf 	:	val_out <= 16'hf5d6;
         16'h2fb0, 16'h2fb1, 16'h2fb2, 16'h2fb3, 16'h2fb4, 16'h2fb5, 16'h2fb6, 16'h2fb7 	:	val_out <= 16'hf5e0;
         16'h2fb8, 16'h2fb9, 16'h2fba, 16'h2fbb, 16'h2fbc, 16'h2fbd, 16'h2fbe, 16'h2fbf 	:	val_out <= 16'hf5ea;
         16'h2fc0, 16'h2fc1, 16'h2fc2, 16'h2fc3, 16'h2fc4, 16'h2fc5, 16'h2fc6, 16'h2fc7 	:	val_out <= 16'hf5f4;
         16'h2fc8, 16'h2fc9, 16'h2fca, 16'h2fcb, 16'h2fcc, 16'h2fcd, 16'h2fce, 16'h2fcf 	:	val_out <= 16'hf5fd;
         16'h2fd0, 16'h2fd1, 16'h2fd2, 16'h2fd3, 16'h2fd4, 16'h2fd5, 16'h2fd6, 16'h2fd7 	:	val_out <= 16'hf607;
         16'h2fd8, 16'h2fd9, 16'h2fda, 16'h2fdb, 16'h2fdc, 16'h2fdd, 16'h2fde, 16'h2fdf 	:	val_out <= 16'hf611;
         16'h2fe0, 16'h2fe1, 16'h2fe2, 16'h2fe3, 16'h2fe4, 16'h2fe5, 16'h2fe6, 16'h2fe7 	:	val_out <= 16'hf61b;
         16'h2fe8, 16'h2fe9, 16'h2fea, 16'h2feb, 16'h2fec, 16'h2fed, 16'h2fee, 16'h2fef 	:	val_out <= 16'hf624;
         16'h2ff0, 16'h2ff1, 16'h2ff2, 16'h2ff3, 16'h2ff4, 16'h2ff5, 16'h2ff6, 16'h2ff7 	:	val_out <= 16'hf62e;
         16'h2ff8, 16'h2ff9, 16'h2ffa, 16'h2ffb, 16'h2ffc, 16'h2ffd, 16'h2ffe, 16'h2fff 	:	val_out <= 16'hf638;
         16'h3000, 16'h3001, 16'h3002, 16'h3003, 16'h3004, 16'h3005, 16'h3006, 16'h3007 	:	val_out <= 16'hf641;
         16'h3008, 16'h3009, 16'h300a, 16'h300b, 16'h300c, 16'h300d, 16'h300e, 16'h300f 	:	val_out <= 16'hf64b;
         16'h3010, 16'h3011, 16'h3012, 16'h3013, 16'h3014, 16'h3015, 16'h3016, 16'h3017 	:	val_out <= 16'hf654;
         16'h3018, 16'h3019, 16'h301a, 16'h301b, 16'h301c, 16'h301d, 16'h301e, 16'h301f 	:	val_out <= 16'hf65e;
         16'h3020, 16'h3021, 16'h3022, 16'h3023, 16'h3024, 16'h3025, 16'h3026, 16'h3027 	:	val_out <= 16'hf668;
         16'h3028, 16'h3029, 16'h302a, 16'h302b, 16'h302c, 16'h302d, 16'h302e, 16'h302f 	:	val_out <= 16'hf671;
         16'h3030, 16'h3031, 16'h3032, 16'h3033, 16'h3034, 16'h3035, 16'h3036, 16'h3037 	:	val_out <= 16'hf67b;
         16'h3038, 16'h3039, 16'h303a, 16'h303b, 16'h303c, 16'h303d, 16'h303e, 16'h303f 	:	val_out <= 16'hf684;
         16'h3040, 16'h3041, 16'h3042, 16'h3043, 16'h3044, 16'h3045, 16'h3046, 16'h3047 	:	val_out <= 16'hf68e;
         16'h3048, 16'h3049, 16'h304a, 16'h304b, 16'h304c, 16'h304d, 16'h304e, 16'h304f 	:	val_out <= 16'hf697;
         16'h3050, 16'h3051, 16'h3052, 16'h3053, 16'h3054, 16'h3055, 16'h3056, 16'h3057 	:	val_out <= 16'hf6a0;
         16'h3058, 16'h3059, 16'h305a, 16'h305b, 16'h305c, 16'h305d, 16'h305e, 16'h305f 	:	val_out <= 16'hf6aa;
         16'h3060, 16'h3061, 16'h3062, 16'h3063, 16'h3064, 16'h3065, 16'h3066, 16'h3067 	:	val_out <= 16'hf6b3;
         16'h3068, 16'h3069, 16'h306a, 16'h306b, 16'h306c, 16'h306d, 16'h306e, 16'h306f 	:	val_out <= 16'hf6bd;
         16'h3070, 16'h3071, 16'h3072, 16'h3073, 16'h3074, 16'h3075, 16'h3076, 16'h3077 	:	val_out <= 16'hf6c6;
         16'h3078, 16'h3079, 16'h307a, 16'h307b, 16'h307c, 16'h307d, 16'h307e, 16'h307f 	:	val_out <= 16'hf6cf;
         16'h3080, 16'h3081, 16'h3082, 16'h3083, 16'h3084, 16'h3085, 16'h3086, 16'h3087 	:	val_out <= 16'hf6d9;
         16'h3088, 16'h3089, 16'h308a, 16'h308b, 16'h308c, 16'h308d, 16'h308e, 16'h308f 	:	val_out <= 16'hf6e2;
         16'h3090, 16'h3091, 16'h3092, 16'h3093, 16'h3094, 16'h3095, 16'h3096, 16'h3097 	:	val_out <= 16'hf6eb;
         16'h3098, 16'h3099, 16'h309a, 16'h309b, 16'h309c, 16'h309d, 16'h309e, 16'h309f 	:	val_out <= 16'hf6f5;
         16'h30a0, 16'h30a1, 16'h30a2, 16'h30a3, 16'h30a4, 16'h30a5, 16'h30a6, 16'h30a7 	:	val_out <= 16'hf6fe;
         16'h30a8, 16'h30a9, 16'h30aa, 16'h30ab, 16'h30ac, 16'h30ad, 16'h30ae, 16'h30af 	:	val_out <= 16'hf707;
         16'h30b0, 16'h30b1, 16'h30b2, 16'h30b3, 16'h30b4, 16'h30b5, 16'h30b6, 16'h30b7 	:	val_out <= 16'hf710;
         16'h30b8, 16'h30b9, 16'h30ba, 16'h30bb, 16'h30bc, 16'h30bd, 16'h30be, 16'h30bf 	:	val_out <= 16'hf71a;
         16'h30c0, 16'h30c1, 16'h30c2, 16'h30c3, 16'h30c4, 16'h30c5, 16'h30c6, 16'h30c7 	:	val_out <= 16'hf723;
         16'h30c8, 16'h30c9, 16'h30ca, 16'h30cb, 16'h30cc, 16'h30cd, 16'h30ce, 16'h30cf 	:	val_out <= 16'hf72c;
         16'h30d0, 16'h30d1, 16'h30d2, 16'h30d3, 16'h30d4, 16'h30d5, 16'h30d6, 16'h30d7 	:	val_out <= 16'hf735;
         16'h30d8, 16'h30d9, 16'h30da, 16'h30db, 16'h30dc, 16'h30dd, 16'h30de, 16'h30df 	:	val_out <= 16'hf73e;
         16'h30e0, 16'h30e1, 16'h30e2, 16'h30e3, 16'h30e4, 16'h30e5, 16'h30e6, 16'h30e7 	:	val_out <= 16'hf747;
         16'h30e8, 16'h30e9, 16'h30ea, 16'h30eb, 16'h30ec, 16'h30ed, 16'h30ee, 16'h30ef 	:	val_out <= 16'hf751;
         16'h30f0, 16'h30f1, 16'h30f2, 16'h30f3, 16'h30f4, 16'h30f5, 16'h30f6, 16'h30f7 	:	val_out <= 16'hf75a;
         16'h30f8, 16'h30f9, 16'h30fa, 16'h30fb, 16'h30fc, 16'h30fd, 16'h30fe, 16'h30ff 	:	val_out <= 16'hf763;
         16'h3100, 16'h3101, 16'h3102, 16'h3103, 16'h3104, 16'h3105, 16'h3106, 16'h3107 	:	val_out <= 16'hf76c;
         16'h3108, 16'h3109, 16'h310a, 16'h310b, 16'h310c, 16'h310d, 16'h310e, 16'h310f 	:	val_out <= 16'hf775;
         16'h3110, 16'h3111, 16'h3112, 16'h3113, 16'h3114, 16'h3115, 16'h3116, 16'h3117 	:	val_out <= 16'hf77e;
         16'h3118, 16'h3119, 16'h311a, 16'h311b, 16'h311c, 16'h311d, 16'h311e, 16'h311f 	:	val_out <= 16'hf787;
         16'h3120, 16'h3121, 16'h3122, 16'h3123, 16'h3124, 16'h3125, 16'h3126, 16'h3127 	:	val_out <= 16'hf790;
         16'h3128, 16'h3129, 16'h312a, 16'h312b, 16'h312c, 16'h312d, 16'h312e, 16'h312f 	:	val_out <= 16'hf799;
         16'h3130, 16'h3131, 16'h3132, 16'h3133, 16'h3134, 16'h3135, 16'h3136, 16'h3137 	:	val_out <= 16'hf7a2;
         16'h3138, 16'h3139, 16'h313a, 16'h313b, 16'h313c, 16'h313d, 16'h313e, 16'h313f 	:	val_out <= 16'hf7ab;
         16'h3140, 16'h3141, 16'h3142, 16'h3143, 16'h3144, 16'h3145, 16'h3146, 16'h3147 	:	val_out <= 16'hf7b4;
         16'h3148, 16'h3149, 16'h314a, 16'h314b, 16'h314c, 16'h314d, 16'h314e, 16'h314f 	:	val_out <= 16'hf7bc;
         16'h3150, 16'h3151, 16'h3152, 16'h3153, 16'h3154, 16'h3155, 16'h3156, 16'h3157 	:	val_out <= 16'hf7c5;
         16'h3158, 16'h3159, 16'h315a, 16'h315b, 16'h315c, 16'h315d, 16'h315e, 16'h315f 	:	val_out <= 16'hf7ce;
         16'h3160, 16'h3161, 16'h3162, 16'h3163, 16'h3164, 16'h3165, 16'h3166, 16'h3167 	:	val_out <= 16'hf7d7;
         16'h3168, 16'h3169, 16'h316a, 16'h316b, 16'h316c, 16'h316d, 16'h316e, 16'h316f 	:	val_out <= 16'hf7e0;
         16'h3170, 16'h3171, 16'h3172, 16'h3173, 16'h3174, 16'h3175, 16'h3176, 16'h3177 	:	val_out <= 16'hf7e9;
         16'h3178, 16'h3179, 16'h317a, 16'h317b, 16'h317c, 16'h317d, 16'h317e, 16'h317f 	:	val_out <= 16'hf7f1;
         16'h3180, 16'h3181, 16'h3182, 16'h3183, 16'h3184, 16'h3185, 16'h3186, 16'h3187 	:	val_out <= 16'hf7fa;
         16'h3188, 16'h3189, 16'h318a, 16'h318b, 16'h318c, 16'h318d, 16'h318e, 16'h318f 	:	val_out <= 16'hf803;
         16'h3190, 16'h3191, 16'h3192, 16'h3193, 16'h3194, 16'h3195, 16'h3196, 16'h3197 	:	val_out <= 16'hf80c;
         16'h3198, 16'h3199, 16'h319a, 16'h319b, 16'h319c, 16'h319d, 16'h319e, 16'h319f 	:	val_out <= 16'hf814;
         16'h31a0, 16'h31a1, 16'h31a2, 16'h31a3, 16'h31a4, 16'h31a5, 16'h31a6, 16'h31a7 	:	val_out <= 16'hf81d;
         16'h31a8, 16'h31a9, 16'h31aa, 16'h31ab, 16'h31ac, 16'h31ad, 16'h31ae, 16'h31af 	:	val_out <= 16'hf826;
         16'h31b0, 16'h31b1, 16'h31b2, 16'h31b3, 16'h31b4, 16'h31b5, 16'h31b6, 16'h31b7 	:	val_out <= 16'hf82e;
         16'h31b8, 16'h31b9, 16'h31ba, 16'h31bb, 16'h31bc, 16'h31bd, 16'h31be, 16'h31bf 	:	val_out <= 16'hf837;
         16'h31c0, 16'h31c1, 16'h31c2, 16'h31c3, 16'h31c4, 16'h31c5, 16'h31c6, 16'h31c7 	:	val_out <= 16'hf840;
         16'h31c8, 16'h31c9, 16'h31ca, 16'h31cb, 16'h31cc, 16'h31cd, 16'h31ce, 16'h31cf 	:	val_out <= 16'hf848;
         16'h31d0, 16'h31d1, 16'h31d2, 16'h31d3, 16'h31d4, 16'h31d5, 16'h31d6, 16'h31d7 	:	val_out <= 16'hf851;
         16'h31d8, 16'h31d9, 16'h31da, 16'h31db, 16'h31dc, 16'h31dd, 16'h31de, 16'h31df 	:	val_out <= 16'hf859;
         16'h31e0, 16'h31e1, 16'h31e2, 16'h31e3, 16'h31e4, 16'h31e5, 16'h31e6, 16'h31e7 	:	val_out <= 16'hf862;
         16'h31e8, 16'h31e9, 16'h31ea, 16'h31eb, 16'h31ec, 16'h31ed, 16'h31ee, 16'h31ef 	:	val_out <= 16'hf86b;
         16'h31f0, 16'h31f1, 16'h31f2, 16'h31f3, 16'h31f4, 16'h31f5, 16'h31f6, 16'h31f7 	:	val_out <= 16'hf873;
         16'h31f8, 16'h31f9, 16'h31fa, 16'h31fb, 16'h31fc, 16'h31fd, 16'h31fe, 16'h31ff 	:	val_out <= 16'hf87c;
         16'h3200, 16'h3201, 16'h3202, 16'h3203, 16'h3204, 16'h3205, 16'h3206, 16'h3207 	:	val_out <= 16'hf884;
         16'h3208, 16'h3209, 16'h320a, 16'h320b, 16'h320c, 16'h320d, 16'h320e, 16'h320f 	:	val_out <= 16'hf88c;
         16'h3210, 16'h3211, 16'h3212, 16'h3213, 16'h3214, 16'h3215, 16'h3216, 16'h3217 	:	val_out <= 16'hf895;
         16'h3218, 16'h3219, 16'h321a, 16'h321b, 16'h321c, 16'h321d, 16'h321e, 16'h321f 	:	val_out <= 16'hf89d;
         16'h3220, 16'h3221, 16'h3222, 16'h3223, 16'h3224, 16'h3225, 16'h3226, 16'h3227 	:	val_out <= 16'hf8a6;
         16'h3228, 16'h3229, 16'h322a, 16'h322b, 16'h322c, 16'h322d, 16'h322e, 16'h322f 	:	val_out <= 16'hf8ae;
         16'h3230, 16'h3231, 16'h3232, 16'h3233, 16'h3234, 16'h3235, 16'h3236, 16'h3237 	:	val_out <= 16'hf8b6;
         16'h3238, 16'h3239, 16'h323a, 16'h323b, 16'h323c, 16'h323d, 16'h323e, 16'h323f 	:	val_out <= 16'hf8bf;
         16'h3240, 16'h3241, 16'h3242, 16'h3243, 16'h3244, 16'h3245, 16'h3246, 16'h3247 	:	val_out <= 16'hf8c7;
         16'h3248, 16'h3249, 16'h324a, 16'h324b, 16'h324c, 16'h324d, 16'h324e, 16'h324f 	:	val_out <= 16'hf8cf;
         16'h3250, 16'h3251, 16'h3252, 16'h3253, 16'h3254, 16'h3255, 16'h3256, 16'h3257 	:	val_out <= 16'hf8d8;
         16'h3258, 16'h3259, 16'h325a, 16'h325b, 16'h325c, 16'h325d, 16'h325e, 16'h325f 	:	val_out <= 16'hf8e0;
         16'h3260, 16'h3261, 16'h3262, 16'h3263, 16'h3264, 16'h3265, 16'h3266, 16'h3267 	:	val_out <= 16'hf8e8;
         16'h3268, 16'h3269, 16'h326a, 16'h326b, 16'h326c, 16'h326d, 16'h326e, 16'h326f 	:	val_out <= 16'hf8f1;
         16'h3270, 16'h3271, 16'h3272, 16'h3273, 16'h3274, 16'h3275, 16'h3276, 16'h3277 	:	val_out <= 16'hf8f9;
         16'h3278, 16'h3279, 16'h327a, 16'h327b, 16'h327c, 16'h327d, 16'h327e, 16'h327f 	:	val_out <= 16'hf901;
         16'h3280, 16'h3281, 16'h3282, 16'h3283, 16'h3284, 16'h3285, 16'h3286, 16'h3287 	:	val_out <= 16'hf909;
         16'h3288, 16'h3289, 16'h328a, 16'h328b, 16'h328c, 16'h328d, 16'h328e, 16'h328f 	:	val_out <= 16'hf911;
         16'h3290, 16'h3291, 16'h3292, 16'h3293, 16'h3294, 16'h3295, 16'h3296, 16'h3297 	:	val_out <= 16'hf919;
         16'h3298, 16'h3299, 16'h329a, 16'h329b, 16'h329c, 16'h329d, 16'h329e, 16'h329f 	:	val_out <= 16'hf922;
         16'h32a0, 16'h32a1, 16'h32a2, 16'h32a3, 16'h32a4, 16'h32a5, 16'h32a6, 16'h32a7 	:	val_out <= 16'hf92a;
         16'h32a8, 16'h32a9, 16'h32aa, 16'h32ab, 16'h32ac, 16'h32ad, 16'h32ae, 16'h32af 	:	val_out <= 16'hf932;
         16'h32b0, 16'h32b1, 16'h32b2, 16'h32b3, 16'h32b4, 16'h32b5, 16'h32b6, 16'h32b7 	:	val_out <= 16'hf93a;
         16'h32b8, 16'h32b9, 16'h32ba, 16'h32bb, 16'h32bc, 16'h32bd, 16'h32be, 16'h32bf 	:	val_out <= 16'hf942;
         16'h32c0, 16'h32c1, 16'h32c2, 16'h32c3, 16'h32c4, 16'h32c5, 16'h32c6, 16'h32c7 	:	val_out <= 16'hf94a;
         16'h32c8, 16'h32c9, 16'h32ca, 16'h32cb, 16'h32cc, 16'h32cd, 16'h32ce, 16'h32cf 	:	val_out <= 16'hf952;
         16'h32d0, 16'h32d1, 16'h32d2, 16'h32d3, 16'h32d4, 16'h32d5, 16'h32d6, 16'h32d7 	:	val_out <= 16'hf95a;
         16'h32d8, 16'h32d9, 16'h32da, 16'h32db, 16'h32dc, 16'h32dd, 16'h32de, 16'h32df 	:	val_out <= 16'hf962;
         16'h32e0, 16'h32e1, 16'h32e2, 16'h32e3, 16'h32e4, 16'h32e5, 16'h32e6, 16'h32e7 	:	val_out <= 16'hf96a;
         16'h32e8, 16'h32e9, 16'h32ea, 16'h32eb, 16'h32ec, 16'h32ed, 16'h32ee, 16'h32ef 	:	val_out <= 16'hf972;
         16'h32f0, 16'h32f1, 16'h32f2, 16'h32f3, 16'h32f4, 16'h32f5, 16'h32f6, 16'h32f7 	:	val_out <= 16'hf97a;
         16'h32f8, 16'h32f9, 16'h32fa, 16'h32fb, 16'h32fc, 16'h32fd, 16'h32fe, 16'h32ff 	:	val_out <= 16'hf982;
         16'h3300, 16'h3301, 16'h3302, 16'h3303, 16'h3304, 16'h3305, 16'h3306, 16'h3307 	:	val_out <= 16'hf98a;
         16'h3308, 16'h3309, 16'h330a, 16'h330b, 16'h330c, 16'h330d, 16'h330e, 16'h330f 	:	val_out <= 16'hf992;
         16'h3310, 16'h3311, 16'h3312, 16'h3313, 16'h3314, 16'h3315, 16'h3316, 16'h3317 	:	val_out <= 16'hf999;
         16'h3318, 16'h3319, 16'h331a, 16'h331b, 16'h331c, 16'h331d, 16'h331e, 16'h331f 	:	val_out <= 16'hf9a1;
         16'h3320, 16'h3321, 16'h3322, 16'h3323, 16'h3324, 16'h3325, 16'h3326, 16'h3327 	:	val_out <= 16'hf9a9;
         16'h3328, 16'h3329, 16'h332a, 16'h332b, 16'h332c, 16'h332d, 16'h332e, 16'h332f 	:	val_out <= 16'hf9b1;
         16'h3330, 16'h3331, 16'h3332, 16'h3333, 16'h3334, 16'h3335, 16'h3336, 16'h3337 	:	val_out <= 16'hf9b9;
         16'h3338, 16'h3339, 16'h333a, 16'h333b, 16'h333c, 16'h333d, 16'h333e, 16'h333f 	:	val_out <= 16'hf9c0;
         16'h3340, 16'h3341, 16'h3342, 16'h3343, 16'h3344, 16'h3345, 16'h3346, 16'h3347 	:	val_out <= 16'hf9c8;
         16'h3348, 16'h3349, 16'h334a, 16'h334b, 16'h334c, 16'h334d, 16'h334e, 16'h334f 	:	val_out <= 16'hf9d0;
         16'h3350, 16'h3351, 16'h3352, 16'h3353, 16'h3354, 16'h3355, 16'h3356, 16'h3357 	:	val_out <= 16'hf9d8;
         16'h3358, 16'h3359, 16'h335a, 16'h335b, 16'h335c, 16'h335d, 16'h335e, 16'h335f 	:	val_out <= 16'hf9df;
         16'h3360, 16'h3361, 16'h3362, 16'h3363, 16'h3364, 16'h3365, 16'h3366, 16'h3367 	:	val_out <= 16'hf9e7;
         16'h3368, 16'h3369, 16'h336a, 16'h336b, 16'h336c, 16'h336d, 16'h336e, 16'h336f 	:	val_out <= 16'hf9ef;
         16'h3370, 16'h3371, 16'h3372, 16'h3373, 16'h3374, 16'h3375, 16'h3376, 16'h3377 	:	val_out <= 16'hf9f6;
         16'h3378, 16'h3379, 16'h337a, 16'h337b, 16'h337c, 16'h337d, 16'h337e, 16'h337f 	:	val_out <= 16'hf9fe;
         16'h3380, 16'h3381, 16'h3382, 16'h3383, 16'h3384, 16'h3385, 16'h3386, 16'h3387 	:	val_out <= 16'hfa05;
         16'h3388, 16'h3389, 16'h338a, 16'h338b, 16'h338c, 16'h338d, 16'h338e, 16'h338f 	:	val_out <= 16'hfa0d;
         16'h3390, 16'h3391, 16'h3392, 16'h3393, 16'h3394, 16'h3395, 16'h3396, 16'h3397 	:	val_out <= 16'hfa15;
         16'h3398, 16'h3399, 16'h339a, 16'h339b, 16'h339c, 16'h339d, 16'h339e, 16'h339f 	:	val_out <= 16'hfa1c;
         16'h33a0, 16'h33a1, 16'h33a2, 16'h33a3, 16'h33a4, 16'h33a5, 16'h33a6, 16'h33a7 	:	val_out <= 16'hfa24;
         16'h33a8, 16'h33a9, 16'h33aa, 16'h33ab, 16'h33ac, 16'h33ad, 16'h33ae, 16'h33af 	:	val_out <= 16'hfa2b;
         16'h33b0, 16'h33b1, 16'h33b2, 16'h33b3, 16'h33b4, 16'h33b5, 16'h33b6, 16'h33b7 	:	val_out <= 16'hfa33;
         16'h33b8, 16'h33b9, 16'h33ba, 16'h33bb, 16'h33bc, 16'h33bd, 16'h33be, 16'h33bf 	:	val_out <= 16'hfa3a;
         16'h33c0, 16'h33c1, 16'h33c2, 16'h33c3, 16'h33c4, 16'h33c5, 16'h33c6, 16'h33c7 	:	val_out <= 16'hfa42;
         16'h33c8, 16'h33c9, 16'h33ca, 16'h33cb, 16'h33cc, 16'h33cd, 16'h33ce, 16'h33cf 	:	val_out <= 16'hfa49;
         16'h33d0, 16'h33d1, 16'h33d2, 16'h33d3, 16'h33d4, 16'h33d5, 16'h33d6, 16'h33d7 	:	val_out <= 16'hfa50;
         16'h33d8, 16'h33d9, 16'h33da, 16'h33db, 16'h33dc, 16'h33dd, 16'h33de, 16'h33df 	:	val_out <= 16'hfa58;
         16'h33e0, 16'h33e1, 16'h33e2, 16'h33e3, 16'h33e4, 16'h33e5, 16'h33e6, 16'h33e7 	:	val_out <= 16'hfa5f;
         16'h33e8, 16'h33e9, 16'h33ea, 16'h33eb, 16'h33ec, 16'h33ed, 16'h33ee, 16'h33ef 	:	val_out <= 16'hfa67;
         16'h33f0, 16'h33f1, 16'h33f2, 16'h33f3, 16'h33f4, 16'h33f5, 16'h33f6, 16'h33f7 	:	val_out <= 16'hfa6e;
         16'h33f8, 16'h33f9, 16'h33fa, 16'h33fb, 16'h33fc, 16'h33fd, 16'h33fe, 16'h33ff 	:	val_out <= 16'hfa75;
         16'h3400, 16'h3401, 16'h3402, 16'h3403, 16'h3404, 16'h3405, 16'h3406, 16'h3407 	:	val_out <= 16'hfa7d;
         16'h3408, 16'h3409, 16'h340a, 16'h340b, 16'h340c, 16'h340d, 16'h340e, 16'h340f 	:	val_out <= 16'hfa84;
         16'h3410, 16'h3411, 16'h3412, 16'h3413, 16'h3414, 16'h3415, 16'h3416, 16'h3417 	:	val_out <= 16'hfa8b;
         16'h3418, 16'h3419, 16'h341a, 16'h341b, 16'h341c, 16'h341d, 16'h341e, 16'h341f 	:	val_out <= 16'hfa92;
         16'h3420, 16'h3421, 16'h3422, 16'h3423, 16'h3424, 16'h3425, 16'h3426, 16'h3427 	:	val_out <= 16'hfa9a;
         16'h3428, 16'h3429, 16'h342a, 16'h342b, 16'h342c, 16'h342d, 16'h342e, 16'h342f 	:	val_out <= 16'hfaa1;
         16'h3430, 16'h3431, 16'h3432, 16'h3433, 16'h3434, 16'h3435, 16'h3436, 16'h3437 	:	val_out <= 16'hfaa8;
         16'h3438, 16'h3439, 16'h343a, 16'h343b, 16'h343c, 16'h343d, 16'h343e, 16'h343f 	:	val_out <= 16'hfaaf;
         16'h3440, 16'h3441, 16'h3442, 16'h3443, 16'h3444, 16'h3445, 16'h3446, 16'h3447 	:	val_out <= 16'hfab6;
         16'h3448, 16'h3449, 16'h344a, 16'h344b, 16'h344c, 16'h344d, 16'h344e, 16'h344f 	:	val_out <= 16'hfabd;
         16'h3450, 16'h3451, 16'h3452, 16'h3453, 16'h3454, 16'h3455, 16'h3456, 16'h3457 	:	val_out <= 16'hfac5;
         16'h3458, 16'h3459, 16'h345a, 16'h345b, 16'h345c, 16'h345d, 16'h345e, 16'h345f 	:	val_out <= 16'hfacc;
         16'h3460, 16'h3461, 16'h3462, 16'h3463, 16'h3464, 16'h3465, 16'h3466, 16'h3467 	:	val_out <= 16'hfad3;
         16'h3468, 16'h3469, 16'h346a, 16'h346b, 16'h346c, 16'h346d, 16'h346e, 16'h346f 	:	val_out <= 16'hfada;
         16'h3470, 16'h3471, 16'h3472, 16'h3473, 16'h3474, 16'h3475, 16'h3476, 16'h3477 	:	val_out <= 16'hfae1;
         16'h3478, 16'h3479, 16'h347a, 16'h347b, 16'h347c, 16'h347d, 16'h347e, 16'h347f 	:	val_out <= 16'hfae8;
         16'h3480, 16'h3481, 16'h3482, 16'h3483, 16'h3484, 16'h3485, 16'h3486, 16'h3487 	:	val_out <= 16'hfaef;
         16'h3488, 16'h3489, 16'h348a, 16'h348b, 16'h348c, 16'h348d, 16'h348e, 16'h348f 	:	val_out <= 16'hfaf6;
         16'h3490, 16'h3491, 16'h3492, 16'h3493, 16'h3494, 16'h3495, 16'h3496, 16'h3497 	:	val_out <= 16'hfafd;
         16'h3498, 16'h3499, 16'h349a, 16'h349b, 16'h349c, 16'h349d, 16'h349e, 16'h349f 	:	val_out <= 16'hfb04;
         16'h34a0, 16'h34a1, 16'h34a2, 16'h34a3, 16'h34a4, 16'h34a5, 16'h34a6, 16'h34a7 	:	val_out <= 16'hfb0b;
         16'h34a8, 16'h34a9, 16'h34aa, 16'h34ab, 16'h34ac, 16'h34ad, 16'h34ae, 16'h34af 	:	val_out <= 16'hfb12;
         16'h34b0, 16'h34b1, 16'h34b2, 16'h34b3, 16'h34b4, 16'h34b5, 16'h34b6, 16'h34b7 	:	val_out <= 16'hfb19;
         16'h34b8, 16'h34b9, 16'h34ba, 16'h34bb, 16'h34bc, 16'h34bd, 16'h34be, 16'h34bf 	:	val_out <= 16'hfb1f;
         16'h34c0, 16'h34c1, 16'h34c2, 16'h34c3, 16'h34c4, 16'h34c5, 16'h34c6, 16'h34c7 	:	val_out <= 16'hfb26;
         16'h34c8, 16'h34c9, 16'h34ca, 16'h34cb, 16'h34cc, 16'h34cd, 16'h34ce, 16'h34cf 	:	val_out <= 16'hfb2d;
         16'h34d0, 16'h34d1, 16'h34d2, 16'h34d3, 16'h34d4, 16'h34d5, 16'h34d6, 16'h34d7 	:	val_out <= 16'hfb34;
         16'h34d8, 16'h34d9, 16'h34da, 16'h34db, 16'h34dc, 16'h34dd, 16'h34de, 16'h34df 	:	val_out <= 16'hfb3b;
         16'h34e0, 16'h34e1, 16'h34e2, 16'h34e3, 16'h34e4, 16'h34e5, 16'h34e6, 16'h34e7 	:	val_out <= 16'hfb42;
         16'h34e8, 16'h34e9, 16'h34ea, 16'h34eb, 16'h34ec, 16'h34ed, 16'h34ee, 16'h34ef 	:	val_out <= 16'hfb48;
         16'h34f0, 16'h34f1, 16'h34f2, 16'h34f3, 16'h34f4, 16'h34f5, 16'h34f6, 16'h34f7 	:	val_out <= 16'hfb4f;
         16'h34f8, 16'h34f9, 16'h34fa, 16'h34fb, 16'h34fc, 16'h34fd, 16'h34fe, 16'h34ff 	:	val_out <= 16'hfb56;
         16'h3500, 16'h3501, 16'h3502, 16'h3503, 16'h3504, 16'h3505, 16'h3506, 16'h3507 	:	val_out <= 16'hfb5d;
         16'h3508, 16'h3509, 16'h350a, 16'h350b, 16'h350c, 16'h350d, 16'h350e, 16'h350f 	:	val_out <= 16'hfb63;
         16'h3510, 16'h3511, 16'h3512, 16'h3513, 16'h3514, 16'h3515, 16'h3516, 16'h3517 	:	val_out <= 16'hfb6a;
         16'h3518, 16'h3519, 16'h351a, 16'h351b, 16'h351c, 16'h351d, 16'h351e, 16'h351f 	:	val_out <= 16'hfb71;
         16'h3520, 16'h3521, 16'h3522, 16'h3523, 16'h3524, 16'h3525, 16'h3526, 16'h3527 	:	val_out <= 16'hfb77;
         16'h3528, 16'h3529, 16'h352a, 16'h352b, 16'h352c, 16'h352d, 16'h352e, 16'h352f 	:	val_out <= 16'hfb7e;
         16'h3530, 16'h3531, 16'h3532, 16'h3533, 16'h3534, 16'h3535, 16'h3536, 16'h3537 	:	val_out <= 16'hfb84;
         16'h3538, 16'h3539, 16'h353a, 16'h353b, 16'h353c, 16'h353d, 16'h353e, 16'h353f 	:	val_out <= 16'hfb8b;
         16'h3540, 16'h3541, 16'h3542, 16'h3543, 16'h3544, 16'h3545, 16'h3546, 16'h3547 	:	val_out <= 16'hfb92;
         16'h3548, 16'h3549, 16'h354a, 16'h354b, 16'h354c, 16'h354d, 16'h354e, 16'h354f 	:	val_out <= 16'hfb98;
         16'h3550, 16'h3551, 16'h3552, 16'h3553, 16'h3554, 16'h3555, 16'h3556, 16'h3557 	:	val_out <= 16'hfb9f;
         16'h3558, 16'h3559, 16'h355a, 16'h355b, 16'h355c, 16'h355d, 16'h355e, 16'h355f 	:	val_out <= 16'hfba5;
         16'h3560, 16'h3561, 16'h3562, 16'h3563, 16'h3564, 16'h3565, 16'h3566, 16'h3567 	:	val_out <= 16'hfbac;
         16'h3568, 16'h3569, 16'h356a, 16'h356b, 16'h356c, 16'h356d, 16'h356e, 16'h356f 	:	val_out <= 16'hfbb2;
         16'h3570, 16'h3571, 16'h3572, 16'h3573, 16'h3574, 16'h3575, 16'h3576, 16'h3577 	:	val_out <= 16'hfbb9;
         16'h3578, 16'h3579, 16'h357a, 16'h357b, 16'h357c, 16'h357d, 16'h357e, 16'h357f 	:	val_out <= 16'hfbbf;
         16'h3580, 16'h3581, 16'h3582, 16'h3583, 16'h3584, 16'h3585, 16'h3586, 16'h3587 	:	val_out <= 16'hfbc5;
         16'h3588, 16'h3589, 16'h358a, 16'h358b, 16'h358c, 16'h358d, 16'h358e, 16'h358f 	:	val_out <= 16'hfbcc;
         16'h3590, 16'h3591, 16'h3592, 16'h3593, 16'h3594, 16'h3595, 16'h3596, 16'h3597 	:	val_out <= 16'hfbd2;
         16'h3598, 16'h3599, 16'h359a, 16'h359b, 16'h359c, 16'h359d, 16'h359e, 16'h359f 	:	val_out <= 16'hfbd9;
         16'h35a0, 16'h35a1, 16'h35a2, 16'h35a3, 16'h35a4, 16'h35a5, 16'h35a6, 16'h35a7 	:	val_out <= 16'hfbdf;
         16'h35a8, 16'h35a9, 16'h35aa, 16'h35ab, 16'h35ac, 16'h35ad, 16'h35ae, 16'h35af 	:	val_out <= 16'hfbe5;
         16'h35b0, 16'h35b1, 16'h35b2, 16'h35b3, 16'h35b4, 16'h35b5, 16'h35b6, 16'h35b7 	:	val_out <= 16'hfbeb;
         16'h35b8, 16'h35b9, 16'h35ba, 16'h35bb, 16'h35bc, 16'h35bd, 16'h35be, 16'h35bf 	:	val_out <= 16'hfbf2;
         16'h35c0, 16'h35c1, 16'h35c2, 16'h35c3, 16'h35c4, 16'h35c5, 16'h35c6, 16'h35c7 	:	val_out <= 16'hfbf8;
         16'h35c8, 16'h35c9, 16'h35ca, 16'h35cb, 16'h35cc, 16'h35cd, 16'h35ce, 16'h35cf 	:	val_out <= 16'hfbfe;
         16'h35d0, 16'h35d1, 16'h35d2, 16'h35d3, 16'h35d4, 16'h35d5, 16'h35d6, 16'h35d7 	:	val_out <= 16'hfc05;
         16'h35d8, 16'h35d9, 16'h35da, 16'h35db, 16'h35dc, 16'h35dd, 16'h35de, 16'h35df 	:	val_out <= 16'hfc0b;
         16'h35e0, 16'h35e1, 16'h35e2, 16'h35e3, 16'h35e4, 16'h35e5, 16'h35e6, 16'h35e7 	:	val_out <= 16'hfc11;
         16'h35e8, 16'h35e9, 16'h35ea, 16'h35eb, 16'h35ec, 16'h35ed, 16'h35ee, 16'h35ef 	:	val_out <= 16'hfc17;
         16'h35f0, 16'h35f1, 16'h35f2, 16'h35f3, 16'h35f4, 16'h35f5, 16'h35f6, 16'h35f7 	:	val_out <= 16'hfc1d;
         16'h35f8, 16'h35f9, 16'h35fa, 16'h35fb, 16'h35fc, 16'h35fd, 16'h35fe, 16'h35ff 	:	val_out <= 16'hfc23;
         16'h3600, 16'h3601, 16'h3602, 16'h3603, 16'h3604, 16'h3605, 16'h3606, 16'h3607 	:	val_out <= 16'hfc29;
         16'h3608, 16'h3609, 16'h360a, 16'h360b, 16'h360c, 16'h360d, 16'h360e, 16'h360f 	:	val_out <= 16'hfc30;
         16'h3610, 16'h3611, 16'h3612, 16'h3613, 16'h3614, 16'h3615, 16'h3616, 16'h3617 	:	val_out <= 16'hfc36;
         16'h3618, 16'h3619, 16'h361a, 16'h361b, 16'h361c, 16'h361d, 16'h361e, 16'h361f 	:	val_out <= 16'hfc3c;
         16'h3620, 16'h3621, 16'h3622, 16'h3623, 16'h3624, 16'h3625, 16'h3626, 16'h3627 	:	val_out <= 16'hfc42;
         16'h3628, 16'h3629, 16'h362a, 16'h362b, 16'h362c, 16'h362d, 16'h362e, 16'h362f 	:	val_out <= 16'hfc48;
         16'h3630, 16'h3631, 16'h3632, 16'h3633, 16'h3634, 16'h3635, 16'h3636, 16'h3637 	:	val_out <= 16'hfc4e;
         16'h3638, 16'h3639, 16'h363a, 16'h363b, 16'h363c, 16'h363d, 16'h363e, 16'h363f 	:	val_out <= 16'hfc54;
         16'h3640, 16'h3641, 16'h3642, 16'h3643, 16'h3644, 16'h3645, 16'h3646, 16'h3647 	:	val_out <= 16'hfc5a;
         16'h3648, 16'h3649, 16'h364a, 16'h364b, 16'h364c, 16'h364d, 16'h364e, 16'h364f 	:	val_out <= 16'hfc60;
         16'h3650, 16'h3651, 16'h3652, 16'h3653, 16'h3654, 16'h3655, 16'h3656, 16'h3657 	:	val_out <= 16'hfc66;
         16'h3658, 16'h3659, 16'h365a, 16'h365b, 16'h365c, 16'h365d, 16'h365e, 16'h365f 	:	val_out <= 16'hfc6c;
         16'h3660, 16'h3661, 16'h3662, 16'h3663, 16'h3664, 16'h3665, 16'h3666, 16'h3667 	:	val_out <= 16'hfc71;
         16'h3668, 16'h3669, 16'h366a, 16'h366b, 16'h366c, 16'h366d, 16'h366e, 16'h366f 	:	val_out <= 16'hfc77;
         16'h3670, 16'h3671, 16'h3672, 16'h3673, 16'h3674, 16'h3675, 16'h3676, 16'h3677 	:	val_out <= 16'hfc7d;
         16'h3678, 16'h3679, 16'h367a, 16'h367b, 16'h367c, 16'h367d, 16'h367e, 16'h367f 	:	val_out <= 16'hfc83;
         16'h3680, 16'h3681, 16'h3682, 16'h3683, 16'h3684, 16'h3685, 16'h3686, 16'h3687 	:	val_out <= 16'hfc89;
         16'h3688, 16'h3689, 16'h368a, 16'h368b, 16'h368c, 16'h368d, 16'h368e, 16'h368f 	:	val_out <= 16'hfc8f;
         16'h3690, 16'h3691, 16'h3692, 16'h3693, 16'h3694, 16'h3695, 16'h3696, 16'h3697 	:	val_out <= 16'hfc94;
         16'h3698, 16'h3699, 16'h369a, 16'h369b, 16'h369c, 16'h369d, 16'h369e, 16'h369f 	:	val_out <= 16'hfc9a;
         16'h36a0, 16'h36a1, 16'h36a2, 16'h36a3, 16'h36a4, 16'h36a5, 16'h36a6, 16'h36a7 	:	val_out <= 16'hfca0;
         16'h36a8, 16'h36a9, 16'h36aa, 16'h36ab, 16'h36ac, 16'h36ad, 16'h36ae, 16'h36af 	:	val_out <= 16'hfca6;
         16'h36b0, 16'h36b1, 16'h36b2, 16'h36b3, 16'h36b4, 16'h36b5, 16'h36b6, 16'h36b7 	:	val_out <= 16'hfcab;
         16'h36b8, 16'h36b9, 16'h36ba, 16'h36bb, 16'h36bc, 16'h36bd, 16'h36be, 16'h36bf 	:	val_out <= 16'hfcb1;
         16'h36c0, 16'h36c1, 16'h36c2, 16'h36c3, 16'h36c4, 16'h36c5, 16'h36c6, 16'h36c7 	:	val_out <= 16'hfcb7;
         16'h36c8, 16'h36c9, 16'h36ca, 16'h36cb, 16'h36cc, 16'h36cd, 16'h36ce, 16'h36cf 	:	val_out <= 16'hfcbc;
         16'h36d0, 16'h36d1, 16'h36d2, 16'h36d3, 16'h36d4, 16'h36d5, 16'h36d6, 16'h36d7 	:	val_out <= 16'hfcc2;
         16'h36d8, 16'h36d9, 16'h36da, 16'h36db, 16'h36dc, 16'h36dd, 16'h36de, 16'h36df 	:	val_out <= 16'hfcc8;
         16'h36e0, 16'h36e1, 16'h36e2, 16'h36e3, 16'h36e4, 16'h36e5, 16'h36e6, 16'h36e7 	:	val_out <= 16'hfccd;
         16'h36e8, 16'h36e9, 16'h36ea, 16'h36eb, 16'h36ec, 16'h36ed, 16'h36ee, 16'h36ef 	:	val_out <= 16'hfcd3;
         16'h36f0, 16'h36f1, 16'h36f2, 16'h36f3, 16'h36f4, 16'h36f5, 16'h36f6, 16'h36f7 	:	val_out <= 16'hfcd8;
         16'h36f8, 16'h36f9, 16'h36fa, 16'h36fb, 16'h36fc, 16'h36fd, 16'h36fe, 16'h36ff 	:	val_out <= 16'hfcde;
         16'h3700, 16'h3701, 16'h3702, 16'h3703, 16'h3704, 16'h3705, 16'h3706, 16'h3707 	:	val_out <= 16'hfce3;
         16'h3708, 16'h3709, 16'h370a, 16'h370b, 16'h370c, 16'h370d, 16'h370e, 16'h370f 	:	val_out <= 16'hfce9;
         16'h3710, 16'h3711, 16'h3712, 16'h3713, 16'h3714, 16'h3715, 16'h3716, 16'h3717 	:	val_out <= 16'hfcee;
         16'h3718, 16'h3719, 16'h371a, 16'h371b, 16'h371c, 16'h371d, 16'h371e, 16'h371f 	:	val_out <= 16'hfcf4;
         16'h3720, 16'h3721, 16'h3722, 16'h3723, 16'h3724, 16'h3725, 16'h3726, 16'h3727 	:	val_out <= 16'hfcf9;
         16'h3728, 16'h3729, 16'h372a, 16'h372b, 16'h372c, 16'h372d, 16'h372e, 16'h372f 	:	val_out <= 16'hfcff;
         16'h3730, 16'h3731, 16'h3732, 16'h3733, 16'h3734, 16'h3735, 16'h3736, 16'h3737 	:	val_out <= 16'hfd04;
         16'h3738, 16'h3739, 16'h373a, 16'h373b, 16'h373c, 16'h373d, 16'h373e, 16'h373f 	:	val_out <= 16'hfd09;
         16'h3740, 16'h3741, 16'h3742, 16'h3743, 16'h3744, 16'h3745, 16'h3746, 16'h3747 	:	val_out <= 16'hfd0f;
         16'h3748, 16'h3749, 16'h374a, 16'h374b, 16'h374c, 16'h374d, 16'h374e, 16'h374f 	:	val_out <= 16'hfd14;
         16'h3750, 16'h3751, 16'h3752, 16'h3753, 16'h3754, 16'h3755, 16'h3756, 16'h3757 	:	val_out <= 16'hfd19;
         16'h3758, 16'h3759, 16'h375a, 16'h375b, 16'h375c, 16'h375d, 16'h375e, 16'h375f 	:	val_out <= 16'hfd1f;
         16'h3760, 16'h3761, 16'h3762, 16'h3763, 16'h3764, 16'h3765, 16'h3766, 16'h3767 	:	val_out <= 16'hfd24;
         16'h3768, 16'h3769, 16'h376a, 16'h376b, 16'h376c, 16'h376d, 16'h376e, 16'h376f 	:	val_out <= 16'hfd29;
         16'h3770, 16'h3771, 16'h3772, 16'h3773, 16'h3774, 16'h3775, 16'h3776, 16'h3777 	:	val_out <= 16'hfd2f;
         16'h3778, 16'h3779, 16'h377a, 16'h377b, 16'h377c, 16'h377d, 16'h377e, 16'h377f 	:	val_out <= 16'hfd34;
         16'h3780, 16'h3781, 16'h3782, 16'h3783, 16'h3784, 16'h3785, 16'h3786, 16'h3787 	:	val_out <= 16'hfd39;
         16'h3788, 16'h3789, 16'h378a, 16'h378b, 16'h378c, 16'h378d, 16'h378e, 16'h378f 	:	val_out <= 16'hfd3e;
         16'h3790, 16'h3791, 16'h3792, 16'h3793, 16'h3794, 16'h3795, 16'h3796, 16'h3797 	:	val_out <= 16'hfd43;
         16'h3798, 16'h3799, 16'h379a, 16'h379b, 16'h379c, 16'h379d, 16'h379e, 16'h379f 	:	val_out <= 16'hfd49;
         16'h37a0, 16'h37a1, 16'h37a2, 16'h37a3, 16'h37a4, 16'h37a5, 16'h37a6, 16'h37a7 	:	val_out <= 16'hfd4e;
         16'h37a8, 16'h37a9, 16'h37aa, 16'h37ab, 16'h37ac, 16'h37ad, 16'h37ae, 16'h37af 	:	val_out <= 16'hfd53;
         16'h37b0, 16'h37b1, 16'h37b2, 16'h37b3, 16'h37b4, 16'h37b5, 16'h37b6, 16'h37b7 	:	val_out <= 16'hfd58;
         16'h37b8, 16'h37b9, 16'h37ba, 16'h37bb, 16'h37bc, 16'h37bd, 16'h37be, 16'h37bf 	:	val_out <= 16'hfd5d;
         16'h37c0, 16'h37c1, 16'h37c2, 16'h37c3, 16'h37c4, 16'h37c5, 16'h37c6, 16'h37c7 	:	val_out <= 16'hfd62;
         16'h37c8, 16'h37c9, 16'h37ca, 16'h37cb, 16'h37cc, 16'h37cd, 16'h37ce, 16'h37cf 	:	val_out <= 16'hfd67;
         16'h37d0, 16'h37d1, 16'h37d2, 16'h37d3, 16'h37d4, 16'h37d5, 16'h37d6, 16'h37d7 	:	val_out <= 16'hfd6c;
         16'h37d8, 16'h37d9, 16'h37da, 16'h37db, 16'h37dc, 16'h37dd, 16'h37de, 16'h37df 	:	val_out <= 16'hfd71;
         16'h37e0, 16'h37e1, 16'h37e2, 16'h37e3, 16'h37e4, 16'h37e5, 16'h37e6, 16'h37e7 	:	val_out <= 16'hfd76;
         16'h37e8, 16'h37e9, 16'h37ea, 16'h37eb, 16'h37ec, 16'h37ed, 16'h37ee, 16'h37ef 	:	val_out <= 16'hfd7b;
         16'h37f0, 16'h37f1, 16'h37f2, 16'h37f3, 16'h37f4, 16'h37f5, 16'h37f6, 16'h37f7 	:	val_out <= 16'hfd80;
         16'h37f8, 16'h37f9, 16'h37fa, 16'h37fb, 16'h37fc, 16'h37fd, 16'h37fe, 16'h37ff 	:	val_out <= 16'hfd85;
         16'h3800, 16'h3801, 16'h3802, 16'h3803, 16'h3804, 16'h3805, 16'h3806, 16'h3807 	:	val_out <= 16'hfd8a;
         16'h3808, 16'h3809, 16'h380a, 16'h380b, 16'h380c, 16'h380d, 16'h380e, 16'h380f 	:	val_out <= 16'hfd8f;
         16'h3810, 16'h3811, 16'h3812, 16'h3813, 16'h3814, 16'h3815, 16'h3816, 16'h3817 	:	val_out <= 16'hfd94;
         16'h3818, 16'h3819, 16'h381a, 16'h381b, 16'h381c, 16'h381d, 16'h381e, 16'h381f 	:	val_out <= 16'hfd98;
         16'h3820, 16'h3821, 16'h3822, 16'h3823, 16'h3824, 16'h3825, 16'h3826, 16'h3827 	:	val_out <= 16'hfd9d;
         16'h3828, 16'h3829, 16'h382a, 16'h382b, 16'h382c, 16'h382d, 16'h382e, 16'h382f 	:	val_out <= 16'hfda2;
         16'h3830, 16'h3831, 16'h3832, 16'h3833, 16'h3834, 16'h3835, 16'h3836, 16'h3837 	:	val_out <= 16'hfda7;
         16'h3838, 16'h3839, 16'h383a, 16'h383b, 16'h383c, 16'h383d, 16'h383e, 16'h383f 	:	val_out <= 16'hfdac;
         16'h3840, 16'h3841, 16'h3842, 16'h3843, 16'h3844, 16'h3845, 16'h3846, 16'h3847 	:	val_out <= 16'hfdb0;
         16'h3848, 16'h3849, 16'h384a, 16'h384b, 16'h384c, 16'h384d, 16'h384e, 16'h384f 	:	val_out <= 16'hfdb5;
         16'h3850, 16'h3851, 16'h3852, 16'h3853, 16'h3854, 16'h3855, 16'h3856, 16'h3857 	:	val_out <= 16'hfdba;
         16'h3858, 16'h3859, 16'h385a, 16'h385b, 16'h385c, 16'h385d, 16'h385e, 16'h385f 	:	val_out <= 16'hfdbf;
         16'h3860, 16'h3861, 16'h3862, 16'h3863, 16'h3864, 16'h3865, 16'h3866, 16'h3867 	:	val_out <= 16'hfdc3;
         16'h3868, 16'h3869, 16'h386a, 16'h386b, 16'h386c, 16'h386d, 16'h386e, 16'h386f 	:	val_out <= 16'hfdc8;
         16'h3870, 16'h3871, 16'h3872, 16'h3873, 16'h3874, 16'h3875, 16'h3876, 16'h3877 	:	val_out <= 16'hfdcd;
         16'h3878, 16'h3879, 16'h387a, 16'h387b, 16'h387c, 16'h387d, 16'h387e, 16'h387f 	:	val_out <= 16'hfdd1;
         16'h3880, 16'h3881, 16'h3882, 16'h3883, 16'h3884, 16'h3885, 16'h3886, 16'h3887 	:	val_out <= 16'hfdd6;
         16'h3888, 16'h3889, 16'h388a, 16'h388b, 16'h388c, 16'h388d, 16'h388e, 16'h388f 	:	val_out <= 16'hfdda;
         16'h3890, 16'h3891, 16'h3892, 16'h3893, 16'h3894, 16'h3895, 16'h3896, 16'h3897 	:	val_out <= 16'hfddf;
         16'h3898, 16'h3899, 16'h389a, 16'h389b, 16'h389c, 16'h389d, 16'h389e, 16'h389f 	:	val_out <= 16'hfde4;
         16'h38a0, 16'h38a1, 16'h38a2, 16'h38a3, 16'h38a4, 16'h38a5, 16'h38a6, 16'h38a7 	:	val_out <= 16'hfde8;
         16'h38a8, 16'h38a9, 16'h38aa, 16'h38ab, 16'h38ac, 16'h38ad, 16'h38ae, 16'h38af 	:	val_out <= 16'hfded;
         16'h38b0, 16'h38b1, 16'h38b2, 16'h38b3, 16'h38b4, 16'h38b5, 16'h38b6, 16'h38b7 	:	val_out <= 16'hfdf1;
         16'h38b8, 16'h38b9, 16'h38ba, 16'h38bb, 16'h38bc, 16'h38bd, 16'h38be, 16'h38bf 	:	val_out <= 16'hfdf6;
         16'h38c0, 16'h38c1, 16'h38c2, 16'h38c3, 16'h38c4, 16'h38c5, 16'h38c6, 16'h38c7 	:	val_out <= 16'hfdfa;
         16'h38c8, 16'h38c9, 16'h38ca, 16'h38cb, 16'h38cc, 16'h38cd, 16'h38ce, 16'h38cf 	:	val_out <= 16'hfdff;
         16'h38d0, 16'h38d1, 16'h38d2, 16'h38d3, 16'h38d4, 16'h38d5, 16'h38d6, 16'h38d7 	:	val_out <= 16'hfe03;
         16'h38d8, 16'h38d9, 16'h38da, 16'h38db, 16'h38dc, 16'h38dd, 16'h38de, 16'h38df 	:	val_out <= 16'hfe07;
         16'h38e0, 16'h38e1, 16'h38e2, 16'h38e3, 16'h38e4, 16'h38e5, 16'h38e6, 16'h38e7 	:	val_out <= 16'hfe0c;
         16'h38e8, 16'h38e9, 16'h38ea, 16'h38eb, 16'h38ec, 16'h38ed, 16'h38ee, 16'h38ef 	:	val_out <= 16'hfe10;
         16'h38f0, 16'h38f1, 16'h38f2, 16'h38f3, 16'h38f4, 16'h38f5, 16'h38f6, 16'h38f7 	:	val_out <= 16'hfe14;
         16'h38f8, 16'h38f9, 16'h38fa, 16'h38fb, 16'h38fc, 16'h38fd, 16'h38fe, 16'h38ff 	:	val_out <= 16'hfe19;
         16'h3900, 16'h3901, 16'h3902, 16'h3903, 16'h3904, 16'h3905, 16'h3906, 16'h3907 	:	val_out <= 16'hfe1d;
         16'h3908, 16'h3909, 16'h390a, 16'h390b, 16'h390c, 16'h390d, 16'h390e, 16'h390f 	:	val_out <= 16'hfe21;
         16'h3910, 16'h3911, 16'h3912, 16'h3913, 16'h3914, 16'h3915, 16'h3916, 16'h3917 	:	val_out <= 16'hfe26;
         16'h3918, 16'h3919, 16'h391a, 16'h391b, 16'h391c, 16'h391d, 16'h391e, 16'h391f 	:	val_out <= 16'hfe2a;
         16'h3920, 16'h3921, 16'h3922, 16'h3923, 16'h3924, 16'h3925, 16'h3926, 16'h3927 	:	val_out <= 16'hfe2e;
         16'h3928, 16'h3929, 16'h392a, 16'h392b, 16'h392c, 16'h392d, 16'h392e, 16'h392f 	:	val_out <= 16'hfe32;
         16'h3930, 16'h3931, 16'h3932, 16'h3933, 16'h3934, 16'h3935, 16'h3936, 16'h3937 	:	val_out <= 16'hfe37;
         16'h3938, 16'h3939, 16'h393a, 16'h393b, 16'h393c, 16'h393d, 16'h393e, 16'h393f 	:	val_out <= 16'hfe3b;
         16'h3940, 16'h3941, 16'h3942, 16'h3943, 16'h3944, 16'h3945, 16'h3946, 16'h3947 	:	val_out <= 16'hfe3f;
         16'h3948, 16'h3949, 16'h394a, 16'h394b, 16'h394c, 16'h394d, 16'h394e, 16'h394f 	:	val_out <= 16'hfe43;
         16'h3950, 16'h3951, 16'h3952, 16'h3953, 16'h3954, 16'h3955, 16'h3956, 16'h3957 	:	val_out <= 16'hfe47;
         16'h3958, 16'h3959, 16'h395a, 16'h395b, 16'h395c, 16'h395d, 16'h395e, 16'h395f 	:	val_out <= 16'hfe4b;
         16'h3960, 16'h3961, 16'h3962, 16'h3963, 16'h3964, 16'h3965, 16'h3966, 16'h3967 	:	val_out <= 16'hfe4f;
         16'h3968, 16'h3969, 16'h396a, 16'h396b, 16'h396c, 16'h396d, 16'h396e, 16'h396f 	:	val_out <= 16'hfe53;
         16'h3970, 16'h3971, 16'h3972, 16'h3973, 16'h3974, 16'h3975, 16'h3976, 16'h3977 	:	val_out <= 16'hfe57;
         16'h3978, 16'h3979, 16'h397a, 16'h397b, 16'h397c, 16'h397d, 16'h397e, 16'h397f 	:	val_out <= 16'hfe5b;
         16'h3980, 16'h3981, 16'h3982, 16'h3983, 16'h3984, 16'h3985, 16'h3986, 16'h3987 	:	val_out <= 16'hfe5f;
         16'h3988, 16'h3989, 16'h398a, 16'h398b, 16'h398c, 16'h398d, 16'h398e, 16'h398f 	:	val_out <= 16'hfe63;
         16'h3990, 16'h3991, 16'h3992, 16'h3993, 16'h3994, 16'h3995, 16'h3996, 16'h3997 	:	val_out <= 16'hfe67;
         16'h3998, 16'h3999, 16'h399a, 16'h399b, 16'h399c, 16'h399d, 16'h399e, 16'h399f 	:	val_out <= 16'hfe6b;
         16'h39a0, 16'h39a1, 16'h39a2, 16'h39a3, 16'h39a4, 16'h39a5, 16'h39a6, 16'h39a7 	:	val_out <= 16'hfe6f;
         16'h39a8, 16'h39a9, 16'h39aa, 16'h39ab, 16'h39ac, 16'h39ad, 16'h39ae, 16'h39af 	:	val_out <= 16'hfe73;
         16'h39b0, 16'h39b1, 16'h39b2, 16'h39b3, 16'h39b4, 16'h39b5, 16'h39b6, 16'h39b7 	:	val_out <= 16'hfe77;
         16'h39b8, 16'h39b9, 16'h39ba, 16'h39bb, 16'h39bc, 16'h39bd, 16'h39be, 16'h39bf 	:	val_out <= 16'hfe7b;
         16'h39c0, 16'h39c1, 16'h39c2, 16'h39c3, 16'h39c4, 16'h39c5, 16'h39c6, 16'h39c7 	:	val_out <= 16'hfe7f;
         16'h39c8, 16'h39c9, 16'h39ca, 16'h39cb, 16'h39cc, 16'h39cd, 16'h39ce, 16'h39cf 	:	val_out <= 16'hfe83;
         16'h39d0, 16'h39d1, 16'h39d2, 16'h39d3, 16'h39d4, 16'h39d5, 16'h39d6, 16'h39d7 	:	val_out <= 16'hfe86;
         16'h39d8, 16'h39d9, 16'h39da, 16'h39db, 16'h39dc, 16'h39dd, 16'h39de, 16'h39df 	:	val_out <= 16'hfe8a;
         16'h39e0, 16'h39e1, 16'h39e2, 16'h39e3, 16'h39e4, 16'h39e5, 16'h39e6, 16'h39e7 	:	val_out <= 16'hfe8e;
         16'h39e8, 16'h39e9, 16'h39ea, 16'h39eb, 16'h39ec, 16'h39ed, 16'h39ee, 16'h39ef 	:	val_out <= 16'hfe92;
         16'h39f0, 16'h39f1, 16'h39f2, 16'h39f3, 16'h39f4, 16'h39f5, 16'h39f6, 16'h39f7 	:	val_out <= 16'hfe95;
         16'h39f8, 16'h39f9, 16'h39fa, 16'h39fb, 16'h39fc, 16'h39fd, 16'h39fe, 16'h39ff 	:	val_out <= 16'hfe99;
         16'h3a00, 16'h3a01, 16'h3a02, 16'h3a03, 16'h3a04, 16'h3a05, 16'h3a06, 16'h3a07 	:	val_out <= 16'hfe9d;
         16'h3a08, 16'h3a09, 16'h3a0a, 16'h3a0b, 16'h3a0c, 16'h3a0d, 16'h3a0e, 16'h3a0f 	:	val_out <= 16'hfea1;
         16'h3a10, 16'h3a11, 16'h3a12, 16'h3a13, 16'h3a14, 16'h3a15, 16'h3a16, 16'h3a17 	:	val_out <= 16'hfea4;
         16'h3a18, 16'h3a19, 16'h3a1a, 16'h3a1b, 16'h3a1c, 16'h3a1d, 16'h3a1e, 16'h3a1f 	:	val_out <= 16'hfea8;
         16'h3a20, 16'h3a21, 16'h3a22, 16'h3a23, 16'h3a24, 16'h3a25, 16'h3a26, 16'h3a27 	:	val_out <= 16'hfeab;
         16'h3a28, 16'h3a29, 16'h3a2a, 16'h3a2b, 16'h3a2c, 16'h3a2d, 16'h3a2e, 16'h3a2f 	:	val_out <= 16'hfeaf;
         16'h3a30, 16'h3a31, 16'h3a32, 16'h3a33, 16'h3a34, 16'h3a35, 16'h3a36, 16'h3a37 	:	val_out <= 16'hfeb3;
         16'h3a38, 16'h3a39, 16'h3a3a, 16'h3a3b, 16'h3a3c, 16'h3a3d, 16'h3a3e, 16'h3a3f 	:	val_out <= 16'hfeb6;
         16'h3a40, 16'h3a41, 16'h3a42, 16'h3a43, 16'h3a44, 16'h3a45, 16'h3a46, 16'h3a47 	:	val_out <= 16'hfeba;
         16'h3a48, 16'h3a49, 16'h3a4a, 16'h3a4b, 16'h3a4c, 16'h3a4d, 16'h3a4e, 16'h3a4f 	:	val_out <= 16'hfebd;
         16'h3a50, 16'h3a51, 16'h3a52, 16'h3a53, 16'h3a54, 16'h3a55, 16'h3a56, 16'h3a57 	:	val_out <= 16'hfec1;
         16'h3a58, 16'h3a59, 16'h3a5a, 16'h3a5b, 16'h3a5c, 16'h3a5d, 16'h3a5e, 16'h3a5f 	:	val_out <= 16'hfec4;
         16'h3a60, 16'h3a61, 16'h3a62, 16'h3a63, 16'h3a64, 16'h3a65, 16'h3a66, 16'h3a67 	:	val_out <= 16'hfec8;
         16'h3a68, 16'h3a69, 16'h3a6a, 16'h3a6b, 16'h3a6c, 16'h3a6d, 16'h3a6e, 16'h3a6f 	:	val_out <= 16'hfecb;
         16'h3a70, 16'h3a71, 16'h3a72, 16'h3a73, 16'h3a74, 16'h3a75, 16'h3a76, 16'h3a77 	:	val_out <= 16'hfecf;
         16'h3a78, 16'h3a79, 16'h3a7a, 16'h3a7b, 16'h3a7c, 16'h3a7d, 16'h3a7e, 16'h3a7f 	:	val_out <= 16'hfed2;
         16'h3a80, 16'h3a81, 16'h3a82, 16'h3a83, 16'h3a84, 16'h3a85, 16'h3a86, 16'h3a87 	:	val_out <= 16'hfed5;
         16'h3a88, 16'h3a89, 16'h3a8a, 16'h3a8b, 16'h3a8c, 16'h3a8d, 16'h3a8e, 16'h3a8f 	:	val_out <= 16'hfed9;
         16'h3a90, 16'h3a91, 16'h3a92, 16'h3a93, 16'h3a94, 16'h3a95, 16'h3a96, 16'h3a97 	:	val_out <= 16'hfedc;
         16'h3a98, 16'h3a99, 16'h3a9a, 16'h3a9b, 16'h3a9c, 16'h3a9d, 16'h3a9e, 16'h3a9f 	:	val_out <= 16'hfedf;
         16'h3aa0, 16'h3aa1, 16'h3aa2, 16'h3aa3, 16'h3aa4, 16'h3aa5, 16'h3aa6, 16'h3aa7 	:	val_out <= 16'hfee3;
         16'h3aa8, 16'h3aa9, 16'h3aaa, 16'h3aab, 16'h3aac, 16'h3aad, 16'h3aae, 16'h3aaf 	:	val_out <= 16'hfee6;
         16'h3ab0, 16'h3ab1, 16'h3ab2, 16'h3ab3, 16'h3ab4, 16'h3ab5, 16'h3ab6, 16'h3ab7 	:	val_out <= 16'hfee9;
         16'h3ab8, 16'h3ab9, 16'h3aba, 16'h3abb, 16'h3abc, 16'h3abd, 16'h3abe, 16'h3abf 	:	val_out <= 16'hfeed;
         16'h3ac0, 16'h3ac1, 16'h3ac2, 16'h3ac3, 16'h3ac4, 16'h3ac5, 16'h3ac6, 16'h3ac7 	:	val_out <= 16'hfef0;
         16'h3ac8, 16'h3ac9, 16'h3aca, 16'h3acb, 16'h3acc, 16'h3acd, 16'h3ace, 16'h3acf 	:	val_out <= 16'hfef3;
         16'h3ad0, 16'h3ad1, 16'h3ad2, 16'h3ad3, 16'h3ad4, 16'h3ad5, 16'h3ad6, 16'h3ad7 	:	val_out <= 16'hfef6;
         16'h3ad8, 16'h3ad9, 16'h3ada, 16'h3adb, 16'h3adc, 16'h3add, 16'h3ade, 16'h3adf 	:	val_out <= 16'hfef9;
         16'h3ae0, 16'h3ae1, 16'h3ae2, 16'h3ae3, 16'h3ae4, 16'h3ae5, 16'h3ae6, 16'h3ae7 	:	val_out <= 16'hfefd;
         16'h3ae8, 16'h3ae9, 16'h3aea, 16'h3aeb, 16'h3aec, 16'h3aed, 16'h3aee, 16'h3aef 	:	val_out <= 16'hff00;
         16'h3af0, 16'h3af1, 16'h3af2, 16'h3af3, 16'h3af4, 16'h3af5, 16'h3af6, 16'h3af7 	:	val_out <= 16'hff03;
         16'h3af8, 16'h3af9, 16'h3afa, 16'h3afb, 16'h3afc, 16'h3afd, 16'h3afe, 16'h3aff 	:	val_out <= 16'hff06;
         16'h3b00, 16'h3b01, 16'h3b02, 16'h3b03, 16'h3b04, 16'h3b05, 16'h3b06, 16'h3b07 	:	val_out <= 16'hff09;
         16'h3b08, 16'h3b09, 16'h3b0a, 16'h3b0b, 16'h3b0c, 16'h3b0d, 16'h3b0e, 16'h3b0f 	:	val_out <= 16'hff0c;
         16'h3b10, 16'h3b11, 16'h3b12, 16'h3b13, 16'h3b14, 16'h3b15, 16'h3b16, 16'h3b17 	:	val_out <= 16'hff0f;
         16'h3b18, 16'h3b19, 16'h3b1a, 16'h3b1b, 16'h3b1c, 16'h3b1d, 16'h3b1e, 16'h3b1f 	:	val_out <= 16'hff12;
         16'h3b20, 16'h3b21, 16'h3b22, 16'h3b23, 16'h3b24, 16'h3b25, 16'h3b26, 16'h3b27 	:	val_out <= 16'hff15;
         16'h3b28, 16'h3b29, 16'h3b2a, 16'h3b2b, 16'h3b2c, 16'h3b2d, 16'h3b2e, 16'h3b2f 	:	val_out <= 16'hff18;
         16'h3b30, 16'h3b31, 16'h3b32, 16'h3b33, 16'h3b34, 16'h3b35, 16'h3b36, 16'h3b37 	:	val_out <= 16'hff1b;
         16'h3b38, 16'h3b39, 16'h3b3a, 16'h3b3b, 16'h3b3c, 16'h3b3d, 16'h3b3e, 16'h3b3f 	:	val_out <= 16'hff1e;
         16'h3b40, 16'h3b41, 16'h3b42, 16'h3b43, 16'h3b44, 16'h3b45, 16'h3b46, 16'h3b47 	:	val_out <= 16'hff21;
         16'h3b48, 16'h3b49, 16'h3b4a, 16'h3b4b, 16'h3b4c, 16'h3b4d, 16'h3b4e, 16'h3b4f 	:	val_out <= 16'hff24;
         16'h3b50, 16'h3b51, 16'h3b52, 16'h3b53, 16'h3b54, 16'h3b55, 16'h3b56, 16'h3b57 	:	val_out <= 16'hff27;
         16'h3b58, 16'h3b59, 16'h3b5a, 16'h3b5b, 16'h3b5c, 16'h3b5d, 16'h3b5e, 16'h3b5f 	:	val_out <= 16'hff2a;
         16'h3b60, 16'h3b61, 16'h3b62, 16'h3b63, 16'h3b64, 16'h3b65, 16'h3b66, 16'h3b67 	:	val_out <= 16'hff2d;
         16'h3b68, 16'h3b69, 16'h3b6a, 16'h3b6b, 16'h3b6c, 16'h3b6d, 16'h3b6e, 16'h3b6f 	:	val_out <= 16'hff2f;
         16'h3b70, 16'h3b71, 16'h3b72, 16'h3b73, 16'h3b74, 16'h3b75, 16'h3b76, 16'h3b77 	:	val_out <= 16'hff32;
         16'h3b78, 16'h3b79, 16'h3b7a, 16'h3b7b, 16'h3b7c, 16'h3b7d, 16'h3b7e, 16'h3b7f 	:	val_out <= 16'hff35;
         16'h3b80, 16'h3b81, 16'h3b82, 16'h3b83, 16'h3b84, 16'h3b85, 16'h3b86, 16'h3b87 	:	val_out <= 16'hff38;
         16'h3b88, 16'h3b89, 16'h3b8a, 16'h3b8b, 16'h3b8c, 16'h3b8d, 16'h3b8e, 16'h3b8f 	:	val_out <= 16'hff3b;
         16'h3b90, 16'h3b91, 16'h3b92, 16'h3b93, 16'h3b94, 16'h3b95, 16'h3b96, 16'h3b97 	:	val_out <= 16'hff3d;
         16'h3b98, 16'h3b99, 16'h3b9a, 16'h3b9b, 16'h3b9c, 16'h3b9d, 16'h3b9e, 16'h3b9f 	:	val_out <= 16'hff40;
         16'h3ba0, 16'h3ba1, 16'h3ba2, 16'h3ba3, 16'h3ba4, 16'h3ba5, 16'h3ba6, 16'h3ba7 	:	val_out <= 16'hff43;
         16'h3ba8, 16'h3ba9, 16'h3baa, 16'h3bab, 16'h3bac, 16'h3bad, 16'h3bae, 16'h3baf 	:	val_out <= 16'hff45;
         16'h3bb0, 16'h3bb1, 16'h3bb2, 16'h3bb3, 16'h3bb4, 16'h3bb5, 16'h3bb6, 16'h3bb7 	:	val_out <= 16'hff48;
         16'h3bb8, 16'h3bb9, 16'h3bba, 16'h3bbb, 16'h3bbc, 16'h3bbd, 16'h3bbe, 16'h3bbf 	:	val_out <= 16'hff4b;
         16'h3bc0, 16'h3bc1, 16'h3bc2, 16'h3bc3, 16'h3bc4, 16'h3bc5, 16'h3bc6, 16'h3bc7 	:	val_out <= 16'hff4d;
         16'h3bc8, 16'h3bc9, 16'h3bca, 16'h3bcb, 16'h3bcc, 16'h3bcd, 16'h3bce, 16'h3bcf 	:	val_out <= 16'hff50;
         16'h3bd0, 16'h3bd1, 16'h3bd2, 16'h3bd3, 16'h3bd4, 16'h3bd5, 16'h3bd6, 16'h3bd7 	:	val_out <= 16'hff53;
         16'h3bd8, 16'h3bd9, 16'h3bda, 16'h3bdb, 16'h3bdc, 16'h3bdd, 16'h3bde, 16'h3bdf 	:	val_out <= 16'hff55;
         16'h3be0, 16'h3be1, 16'h3be2, 16'h3be3, 16'h3be4, 16'h3be5, 16'h3be6, 16'h3be7 	:	val_out <= 16'hff58;
         16'h3be8, 16'h3be9, 16'h3bea, 16'h3beb, 16'h3bec, 16'h3bed, 16'h3bee, 16'h3bef 	:	val_out <= 16'hff5a;
         16'h3bf0, 16'h3bf1, 16'h3bf2, 16'h3bf3, 16'h3bf4, 16'h3bf5, 16'h3bf6, 16'h3bf7 	:	val_out <= 16'hff5d;
         16'h3bf8, 16'h3bf9, 16'h3bfa, 16'h3bfb, 16'h3bfc, 16'h3bfd, 16'h3bfe, 16'h3bff 	:	val_out <= 16'hff5f;
         16'h3c00, 16'h3c01, 16'h3c02, 16'h3c03, 16'h3c04, 16'h3c05, 16'h3c06, 16'h3c07 	:	val_out <= 16'hff62;
         16'h3c08, 16'h3c09, 16'h3c0a, 16'h3c0b, 16'h3c0c, 16'h3c0d, 16'h3c0e, 16'h3c0f 	:	val_out <= 16'hff64;
         16'h3c10, 16'h3c11, 16'h3c12, 16'h3c13, 16'h3c14, 16'h3c15, 16'h3c16, 16'h3c17 	:	val_out <= 16'hff67;
         16'h3c18, 16'h3c19, 16'h3c1a, 16'h3c1b, 16'h3c1c, 16'h3c1d, 16'h3c1e, 16'h3c1f 	:	val_out <= 16'hff69;
         16'h3c20, 16'h3c21, 16'h3c22, 16'h3c23, 16'h3c24, 16'h3c25, 16'h3c26, 16'h3c27 	:	val_out <= 16'hff6b;
         16'h3c28, 16'h3c29, 16'h3c2a, 16'h3c2b, 16'h3c2c, 16'h3c2d, 16'h3c2e, 16'h3c2f 	:	val_out <= 16'hff6e;
         16'h3c30, 16'h3c31, 16'h3c32, 16'h3c33, 16'h3c34, 16'h3c35, 16'h3c36, 16'h3c37 	:	val_out <= 16'hff70;
         16'h3c38, 16'h3c39, 16'h3c3a, 16'h3c3b, 16'h3c3c, 16'h3c3d, 16'h3c3e, 16'h3c3f 	:	val_out <= 16'hff72;
         16'h3c40, 16'h3c41, 16'h3c42, 16'h3c43, 16'h3c44, 16'h3c45, 16'h3c46, 16'h3c47 	:	val_out <= 16'hff75;
         16'h3c48, 16'h3c49, 16'h3c4a, 16'h3c4b, 16'h3c4c, 16'h3c4d, 16'h3c4e, 16'h3c4f 	:	val_out <= 16'hff77;
         16'h3c50, 16'h3c51, 16'h3c52, 16'h3c53, 16'h3c54, 16'h3c55, 16'h3c56, 16'h3c57 	:	val_out <= 16'hff79;
         16'h3c58, 16'h3c59, 16'h3c5a, 16'h3c5b, 16'h3c5c, 16'h3c5d, 16'h3c5e, 16'h3c5f 	:	val_out <= 16'hff7c;
         16'h3c60, 16'h3c61, 16'h3c62, 16'h3c63, 16'h3c64, 16'h3c65, 16'h3c66, 16'h3c67 	:	val_out <= 16'hff7e;
         16'h3c68, 16'h3c69, 16'h3c6a, 16'h3c6b, 16'h3c6c, 16'h3c6d, 16'h3c6e, 16'h3c6f 	:	val_out <= 16'hff80;
         16'h3c70, 16'h3c71, 16'h3c72, 16'h3c73, 16'h3c74, 16'h3c75, 16'h3c76, 16'h3c77 	:	val_out <= 16'hff82;
         16'h3c78, 16'h3c79, 16'h3c7a, 16'h3c7b, 16'h3c7c, 16'h3c7d, 16'h3c7e, 16'h3c7f 	:	val_out <= 16'hff85;
         16'h3c80, 16'h3c81, 16'h3c82, 16'h3c83, 16'h3c84, 16'h3c85, 16'h3c86, 16'h3c87 	:	val_out <= 16'hff87;
         16'h3c88, 16'h3c89, 16'h3c8a, 16'h3c8b, 16'h3c8c, 16'h3c8d, 16'h3c8e, 16'h3c8f 	:	val_out <= 16'hff89;
         16'h3c90, 16'h3c91, 16'h3c92, 16'h3c93, 16'h3c94, 16'h3c95, 16'h3c96, 16'h3c97 	:	val_out <= 16'hff8b;
         16'h3c98, 16'h3c99, 16'h3c9a, 16'h3c9b, 16'h3c9c, 16'h3c9d, 16'h3c9e, 16'h3c9f 	:	val_out <= 16'hff8d;
         16'h3ca0, 16'h3ca1, 16'h3ca2, 16'h3ca3, 16'h3ca4, 16'h3ca5, 16'h3ca6, 16'h3ca7 	:	val_out <= 16'hff8f;
         16'h3ca8, 16'h3ca9, 16'h3caa, 16'h3cab, 16'h3cac, 16'h3cad, 16'h3cae, 16'h3caf 	:	val_out <= 16'hff91;
         16'h3cb0, 16'h3cb1, 16'h3cb2, 16'h3cb3, 16'h3cb4, 16'h3cb5, 16'h3cb6, 16'h3cb7 	:	val_out <= 16'hff93;
         16'h3cb8, 16'h3cb9, 16'h3cba, 16'h3cbb, 16'h3cbc, 16'h3cbd, 16'h3cbe, 16'h3cbf 	:	val_out <= 16'hff95;
         16'h3cc0, 16'h3cc1, 16'h3cc2, 16'h3cc3, 16'h3cc4, 16'h3cc5, 16'h3cc6, 16'h3cc7 	:	val_out <= 16'hff97;
         16'h3cc8, 16'h3cc9, 16'h3cca, 16'h3ccb, 16'h3ccc, 16'h3ccd, 16'h3cce, 16'h3ccf 	:	val_out <= 16'hff99;
         16'h3cd0, 16'h3cd1, 16'h3cd2, 16'h3cd3, 16'h3cd4, 16'h3cd5, 16'h3cd6, 16'h3cd7 	:	val_out <= 16'hff9b;
         16'h3cd8, 16'h3cd9, 16'h3cda, 16'h3cdb, 16'h3cdc, 16'h3cdd, 16'h3cde, 16'h3cdf 	:	val_out <= 16'hff9d;
         16'h3ce0, 16'h3ce1, 16'h3ce2, 16'h3ce3, 16'h3ce4, 16'h3ce5, 16'h3ce6, 16'h3ce7 	:	val_out <= 16'hff9f;
         16'h3ce8, 16'h3ce9, 16'h3cea, 16'h3ceb, 16'h3cec, 16'h3ced, 16'h3cee, 16'h3cef 	:	val_out <= 16'hffa1;
         16'h3cf0, 16'h3cf1, 16'h3cf2, 16'h3cf3, 16'h3cf4, 16'h3cf5, 16'h3cf6, 16'h3cf7 	:	val_out <= 16'hffa3;
         16'h3cf8, 16'h3cf9, 16'h3cfa, 16'h3cfb, 16'h3cfc, 16'h3cfd, 16'h3cfe, 16'h3cff 	:	val_out <= 16'hffa5;
         16'h3d00, 16'h3d01, 16'h3d02, 16'h3d03, 16'h3d04, 16'h3d05, 16'h3d06, 16'h3d07 	:	val_out <= 16'hffa7;
         16'h3d08, 16'h3d09, 16'h3d0a, 16'h3d0b, 16'h3d0c, 16'h3d0d, 16'h3d0e, 16'h3d0f 	:	val_out <= 16'hffa9;
         16'h3d10, 16'h3d11, 16'h3d12, 16'h3d13, 16'h3d14, 16'h3d15, 16'h3d16, 16'h3d17 	:	val_out <= 16'hffaa;
         16'h3d18, 16'h3d19, 16'h3d1a, 16'h3d1b, 16'h3d1c, 16'h3d1d, 16'h3d1e, 16'h3d1f 	:	val_out <= 16'hffac;
         16'h3d20, 16'h3d21, 16'h3d22, 16'h3d23, 16'h3d24, 16'h3d25, 16'h3d26, 16'h3d27 	:	val_out <= 16'hffae;
         16'h3d28, 16'h3d29, 16'h3d2a, 16'h3d2b, 16'h3d2c, 16'h3d2d, 16'h3d2e, 16'h3d2f 	:	val_out <= 16'hffb0;
         16'h3d30, 16'h3d31, 16'h3d32, 16'h3d33, 16'h3d34, 16'h3d35, 16'h3d36, 16'h3d37 	:	val_out <= 16'hffb1;
         16'h3d38, 16'h3d39, 16'h3d3a, 16'h3d3b, 16'h3d3c, 16'h3d3d, 16'h3d3e, 16'h3d3f 	:	val_out <= 16'hffb3;
         16'h3d40, 16'h3d41, 16'h3d42, 16'h3d43, 16'h3d44, 16'h3d45, 16'h3d46, 16'h3d47 	:	val_out <= 16'hffb5;
         16'h3d48, 16'h3d49, 16'h3d4a, 16'h3d4b, 16'h3d4c, 16'h3d4d, 16'h3d4e, 16'h3d4f 	:	val_out <= 16'hffb7;
         16'h3d50, 16'h3d51, 16'h3d52, 16'h3d53, 16'h3d54, 16'h3d55, 16'h3d56, 16'h3d57 	:	val_out <= 16'hffb8;
         16'h3d58, 16'h3d59, 16'h3d5a, 16'h3d5b, 16'h3d5c, 16'h3d5d, 16'h3d5e, 16'h3d5f 	:	val_out <= 16'hffba;
         16'h3d60, 16'h3d61, 16'h3d62, 16'h3d63, 16'h3d64, 16'h3d65, 16'h3d66, 16'h3d67 	:	val_out <= 16'hffbc;
         16'h3d68, 16'h3d69, 16'h3d6a, 16'h3d6b, 16'h3d6c, 16'h3d6d, 16'h3d6e, 16'h3d6f 	:	val_out <= 16'hffbd;
         16'h3d70, 16'h3d71, 16'h3d72, 16'h3d73, 16'h3d74, 16'h3d75, 16'h3d76, 16'h3d77 	:	val_out <= 16'hffbf;
         16'h3d78, 16'h3d79, 16'h3d7a, 16'h3d7b, 16'h3d7c, 16'h3d7d, 16'h3d7e, 16'h3d7f 	:	val_out <= 16'hffc0;
         16'h3d80, 16'h3d81, 16'h3d82, 16'h3d83, 16'h3d84, 16'h3d85, 16'h3d86, 16'h3d87 	:	val_out <= 16'hffc2;
         16'h3d88, 16'h3d89, 16'h3d8a, 16'h3d8b, 16'h3d8c, 16'h3d8d, 16'h3d8e, 16'h3d8f 	:	val_out <= 16'hffc3;
         16'h3d90, 16'h3d91, 16'h3d92, 16'h3d93, 16'h3d94, 16'h3d95, 16'h3d96, 16'h3d97 	:	val_out <= 16'hffc5;
         16'h3d98, 16'h3d99, 16'h3d9a, 16'h3d9b, 16'h3d9c, 16'h3d9d, 16'h3d9e, 16'h3d9f 	:	val_out <= 16'hffc6;
         16'h3da0, 16'h3da1, 16'h3da2, 16'h3da3, 16'h3da4, 16'h3da5, 16'h3da6, 16'h3da7 	:	val_out <= 16'hffc8;
         16'h3da8, 16'h3da9, 16'h3daa, 16'h3dab, 16'h3dac, 16'h3dad, 16'h3dae, 16'h3daf 	:	val_out <= 16'hffc9;
         16'h3db0, 16'h3db1, 16'h3db2, 16'h3db3, 16'h3db4, 16'h3db5, 16'h3db6, 16'h3db7 	:	val_out <= 16'hffcb;
         16'h3db8, 16'h3db9, 16'h3dba, 16'h3dbb, 16'h3dbc, 16'h3dbd, 16'h3dbe, 16'h3dbf 	:	val_out <= 16'hffcc;
         16'h3dc0, 16'h3dc1, 16'h3dc2, 16'h3dc3, 16'h3dc4, 16'h3dc5, 16'h3dc6, 16'h3dc7 	:	val_out <= 16'hffce;
         16'h3dc8, 16'h3dc9, 16'h3dca, 16'h3dcb, 16'h3dcc, 16'h3dcd, 16'h3dce, 16'h3dcf 	:	val_out <= 16'hffcf;
         16'h3dd0, 16'h3dd1, 16'h3dd2, 16'h3dd3, 16'h3dd4, 16'h3dd5, 16'h3dd6, 16'h3dd7 	:	val_out <= 16'hffd0;
         16'h3dd8, 16'h3dd9, 16'h3dda, 16'h3ddb, 16'h3ddc, 16'h3ddd, 16'h3dde, 16'h3ddf 	:	val_out <= 16'hffd2;
         16'h3de0, 16'h3de1, 16'h3de2, 16'h3de3, 16'h3de4, 16'h3de5, 16'h3de6, 16'h3de7 	:	val_out <= 16'hffd3;
         16'h3de8, 16'h3de9, 16'h3dea, 16'h3deb, 16'h3dec, 16'h3ded, 16'h3dee, 16'h3def 	:	val_out <= 16'hffd4;
         16'h3df0, 16'h3df1, 16'h3df2, 16'h3df3, 16'h3df4, 16'h3df5, 16'h3df6, 16'h3df7 	:	val_out <= 16'hffd6;
         16'h3df8, 16'h3df9, 16'h3dfa, 16'h3dfb, 16'h3dfc, 16'h3dfd, 16'h3dfe, 16'h3dff 	:	val_out <= 16'hffd7;
         16'h3e00, 16'h3e01, 16'h3e02, 16'h3e03, 16'h3e04, 16'h3e05, 16'h3e06, 16'h3e07 	:	val_out <= 16'hffd8;
         16'h3e08, 16'h3e09, 16'h3e0a, 16'h3e0b, 16'h3e0c, 16'h3e0d, 16'h3e0e, 16'h3e0f 	:	val_out <= 16'hffd9;
         16'h3e10, 16'h3e11, 16'h3e12, 16'h3e13, 16'h3e14, 16'h3e15, 16'h3e16, 16'h3e17 	:	val_out <= 16'hffda;
         16'h3e18, 16'h3e19, 16'h3e1a, 16'h3e1b, 16'h3e1c, 16'h3e1d, 16'h3e1e, 16'h3e1f 	:	val_out <= 16'hffdc;
         16'h3e20, 16'h3e21, 16'h3e22, 16'h3e23, 16'h3e24, 16'h3e25, 16'h3e26, 16'h3e27 	:	val_out <= 16'hffdd;
         16'h3e28, 16'h3e29, 16'h3e2a, 16'h3e2b, 16'h3e2c, 16'h3e2d, 16'h3e2e, 16'h3e2f 	:	val_out <= 16'hffde;
         16'h3e30, 16'h3e31, 16'h3e32, 16'h3e33, 16'h3e34, 16'h3e35, 16'h3e36, 16'h3e37 	:	val_out <= 16'hffdf;
         16'h3e38, 16'h3e39, 16'h3e3a, 16'h3e3b, 16'h3e3c, 16'h3e3d, 16'h3e3e, 16'h3e3f 	:	val_out <= 16'hffe0;
         16'h3e40, 16'h3e41, 16'h3e42, 16'h3e43, 16'h3e44, 16'h3e45, 16'h3e46, 16'h3e47 	:	val_out <= 16'hffe1;
         16'h3e48, 16'h3e49, 16'h3e4a, 16'h3e4b, 16'h3e4c, 16'h3e4d, 16'h3e4e, 16'h3e4f 	:	val_out <= 16'hffe2;
         16'h3e50, 16'h3e51, 16'h3e52, 16'h3e53, 16'h3e54, 16'h3e55, 16'h3e56, 16'h3e57 	:	val_out <= 16'hffe3;
         16'h3e58, 16'h3e59, 16'h3e5a, 16'h3e5b, 16'h3e5c, 16'h3e5d, 16'h3e5e, 16'h3e5f 	:	val_out <= 16'hffe4;
         16'h3e60, 16'h3e61, 16'h3e62, 16'h3e63, 16'h3e64, 16'h3e65, 16'h3e66, 16'h3e67 	:	val_out <= 16'hffe5;
         16'h3e68, 16'h3e69, 16'h3e6a, 16'h3e6b, 16'h3e6c, 16'h3e6d, 16'h3e6e, 16'h3e6f 	:	val_out <= 16'hffe6;
         16'h3e70, 16'h3e71, 16'h3e72, 16'h3e73, 16'h3e74, 16'h3e75, 16'h3e76, 16'h3e77 	:	val_out <= 16'hffe7;
         16'h3e78, 16'h3e79, 16'h3e7a, 16'h3e7b, 16'h3e7c, 16'h3e7d, 16'h3e7e, 16'h3e7f 	:	val_out <= 16'hffe8;
         16'h3e80, 16'h3e81, 16'h3e82, 16'h3e83, 16'h3e84, 16'h3e85, 16'h3e86, 16'h3e87 	:	val_out <= 16'hffe9;
         16'h3e88, 16'h3e89, 16'h3e8a, 16'h3e8b, 16'h3e8c, 16'h3e8d, 16'h3e8e, 16'h3e8f 	:	val_out <= 16'hffea;
         16'h3e90, 16'h3e91, 16'h3e92, 16'h3e93, 16'h3e94, 16'h3e95, 16'h3e96, 16'h3e97 	:	val_out <= 16'hffeb;
         16'h3e98, 16'h3e99, 16'h3e9a, 16'h3e9b, 16'h3e9c, 16'h3e9d, 16'h3e9e, 16'h3e9f 	:	val_out <= 16'hffec;
         16'h3ea0, 16'h3ea1, 16'h3ea2, 16'h3ea3, 16'h3ea4, 16'h3ea5, 16'h3ea6, 16'h3ea7 	:	val_out <= 16'hffed;
         16'h3ea8, 16'h3ea9, 16'h3eaa, 16'h3eab, 16'h3eac, 16'h3ead, 16'h3eae, 16'h3eaf 	:	val_out <= 16'hffee;
         16'h3eb0, 16'h3eb1, 16'h3eb2, 16'h3eb3, 16'h3eb4, 16'h3eb5, 16'h3eb6, 16'h3eb7 	:	val_out <= 16'hffee;
         16'h3eb8, 16'h3eb9, 16'h3eba, 16'h3ebb, 16'h3ebc, 16'h3ebd, 16'h3ebe, 16'h3ebf 	:	val_out <= 16'hffef;
         16'h3ec0, 16'h3ec1, 16'h3ec2, 16'h3ec3, 16'h3ec4, 16'h3ec5, 16'h3ec6, 16'h3ec7 	:	val_out <= 16'hfff0;
         16'h3ec8, 16'h3ec9, 16'h3eca, 16'h3ecb, 16'h3ecc, 16'h3ecd, 16'h3ece, 16'h3ecf 	:	val_out <= 16'hfff1;
         16'h3ed0, 16'h3ed1, 16'h3ed2, 16'h3ed3, 16'h3ed4, 16'h3ed5, 16'h3ed6, 16'h3ed7 	:	val_out <= 16'hfff2;
         16'h3ed8, 16'h3ed9, 16'h3eda, 16'h3edb, 16'h3edc, 16'h3edd, 16'h3ede, 16'h3edf 	:	val_out <= 16'hfff2;
         16'h3ee0, 16'h3ee1, 16'h3ee2, 16'h3ee3, 16'h3ee4, 16'h3ee5, 16'h3ee6, 16'h3ee7 	:	val_out <= 16'hfff3;
         16'h3ee8, 16'h3ee9, 16'h3eea, 16'h3eeb, 16'h3eec, 16'h3eed, 16'h3eee, 16'h3eef 	:	val_out <= 16'hfff4;
         16'h3ef0, 16'h3ef1, 16'h3ef2, 16'h3ef3, 16'h3ef4, 16'h3ef5, 16'h3ef6, 16'h3ef7 	:	val_out <= 16'hfff4;
         16'h3ef8, 16'h3ef9, 16'h3efa, 16'h3efb, 16'h3efc, 16'h3efd, 16'h3efe, 16'h3eff 	:	val_out <= 16'hfff5;
         16'h3f00, 16'h3f01, 16'h3f02, 16'h3f03, 16'h3f04, 16'h3f05, 16'h3f06, 16'h3f07 	:	val_out <= 16'hfff6;
         16'h3f08, 16'h3f09, 16'h3f0a, 16'h3f0b, 16'h3f0c, 16'h3f0d, 16'h3f0e, 16'h3f0f 	:	val_out <= 16'hfff6;
         16'h3f10, 16'h3f11, 16'h3f12, 16'h3f13, 16'h3f14, 16'h3f15, 16'h3f16, 16'h3f17 	:	val_out <= 16'hfff7;
         16'h3f18, 16'h3f19, 16'h3f1a, 16'h3f1b, 16'h3f1c, 16'h3f1d, 16'h3f1e, 16'h3f1f 	:	val_out <= 16'hfff7;
         16'h3f20, 16'h3f21, 16'h3f22, 16'h3f23, 16'h3f24, 16'h3f25, 16'h3f26, 16'h3f27 	:	val_out <= 16'hfff8;
         16'h3f28, 16'h3f29, 16'h3f2a, 16'h3f2b, 16'h3f2c, 16'h3f2d, 16'h3f2e, 16'h3f2f 	:	val_out <= 16'hfff8;
         16'h3f30, 16'h3f31, 16'h3f32, 16'h3f33, 16'h3f34, 16'h3f35, 16'h3f36, 16'h3f37 	:	val_out <= 16'hfff9;
         16'h3f38, 16'h3f39, 16'h3f3a, 16'h3f3b, 16'h3f3c, 16'h3f3d, 16'h3f3e, 16'h3f3f 	:	val_out <= 16'hfff9;
         16'h3f40, 16'h3f41, 16'h3f42, 16'h3f43, 16'h3f44, 16'h3f45, 16'h3f46, 16'h3f47 	:	val_out <= 16'hfffa;
         16'h3f48, 16'h3f49, 16'h3f4a, 16'h3f4b, 16'h3f4c, 16'h3f4d, 16'h3f4e, 16'h3f4f 	:	val_out <= 16'hfffa;
         16'h3f50, 16'h3f51, 16'h3f52, 16'h3f53, 16'h3f54, 16'h3f55, 16'h3f56, 16'h3f57 	:	val_out <= 16'hfffb;
         16'h3f58, 16'h3f59, 16'h3f5a, 16'h3f5b, 16'h3f5c, 16'h3f5d, 16'h3f5e, 16'h3f5f 	:	val_out <= 16'hfffb;
         16'h3f60, 16'h3f61, 16'h3f62, 16'h3f63, 16'h3f64, 16'h3f65, 16'h3f66, 16'h3f67 	:	val_out <= 16'hfffc;
         16'h3f68, 16'h3f69, 16'h3f6a, 16'h3f6b, 16'h3f6c, 16'h3f6d, 16'h3f6e, 16'h3f6f 	:	val_out <= 16'hfffc;
         16'h3f70, 16'h3f71, 16'h3f72, 16'h3f73, 16'h3f74, 16'h3f75, 16'h3f76, 16'h3f77 	:	val_out <= 16'hfffc;
         16'h3f78, 16'h3f79, 16'h3f7a, 16'h3f7b, 16'h3f7c, 16'h3f7d, 16'h3f7e, 16'h3f7f 	:	val_out <= 16'hfffd;
         16'h3f80, 16'h3f81, 16'h3f82, 16'h3f83, 16'h3f84, 16'h3f85, 16'h3f86, 16'h3f87 	:	val_out <= 16'hfffd;
         16'h3f88, 16'h3f89, 16'h3f8a, 16'h3f8b, 16'h3f8c, 16'h3f8d, 16'h3f8e, 16'h3f8f 	:	val_out <= 16'hfffd;
         16'h3f90, 16'h3f91, 16'h3f92, 16'h3f93, 16'h3f94, 16'h3f95, 16'h3f96, 16'h3f97 	:	val_out <= 16'hfffe;
         16'h3f98, 16'h3f99, 16'h3f9a, 16'h3f9b, 16'h3f9c, 16'h3f9d, 16'h3f9e, 16'h3f9f 	:	val_out <= 16'hfffe;
         16'h3fa0, 16'h3fa1, 16'h3fa2, 16'h3fa3, 16'h3fa4, 16'h3fa5, 16'h3fa6, 16'h3fa7 	:	val_out <= 16'hfffe;
         16'h3fa8, 16'h3fa9, 16'h3faa, 16'h3fab, 16'h3fac, 16'h3fad, 16'h3fae, 16'h3faf 	:	val_out <= 16'hfffe;
         16'h3fb0, 16'h3fb1, 16'h3fb2, 16'h3fb3, 16'h3fb4, 16'h3fb5, 16'h3fb6, 16'h3fb7 	:	val_out <= 16'hffff;
         16'h3fb8, 16'h3fb9, 16'h3fba, 16'h3fbb, 16'h3fbc, 16'h3fbd, 16'h3fbe, 16'h3fbf 	:	val_out <= 16'hffff;
         16'h3fc0, 16'h3fc1, 16'h3fc2, 16'h3fc3, 16'h3fc4, 16'h3fc5, 16'h3fc6, 16'h3fc7 	:	val_out <= 16'hffff;
         16'h3fc8, 16'h3fc9, 16'h3fca, 16'h3fcb, 16'h3fcc, 16'h3fcd, 16'h3fce, 16'h3fcf 	:	val_out <= 16'hffff;
         16'h3fd0, 16'h3fd1, 16'h3fd2, 16'h3fd3, 16'h3fd4, 16'h3fd5, 16'h3fd6, 16'h3fd7 	:	val_out <= 16'hffff;
         16'h3fd8, 16'h3fd9, 16'h3fda, 16'h3fdb, 16'h3fdc, 16'h3fdd, 16'h3fde, 16'h3fdf 	:	val_out <= 16'hffff;
         16'h3fe0, 16'h3fe1, 16'h3fe2, 16'h3fe3, 16'h3fe4, 16'h3fe5, 16'h3fe6, 16'h3fe7 	:	val_out <= 16'hffff;
         16'h3fe8, 16'h3fe9, 16'h3fea, 16'h3feb, 16'h3fec, 16'h3fed, 16'h3fee, 16'h3fef 	:	val_out <= 16'hffff;
         16'h3ff0, 16'h3ff1, 16'h3ff2, 16'h3ff3, 16'h3ff4, 16'h3ff5, 16'h3ff6, 16'h3ff7 	:	val_out <= 16'hffff;
         16'h3ff8, 16'h3ff9, 16'h3ffa, 16'h3ffb, 16'h3ffc, 16'h3ffd, 16'h3ffe, 16'h3fff 	:	val_out <= 16'hffff;
         16'h4000, 16'h4001, 16'h4002, 16'h4003, 16'h4004, 16'h4005, 16'h4006, 16'h4007 	:	val_out <= 16'h10000;
         16'h4008, 16'h4009, 16'h400a, 16'h400b, 16'h400c, 16'h400d, 16'h400e, 16'h400f 	:	val_out <= 16'hffff;
         16'h4010, 16'h4011, 16'h4012, 16'h4013, 16'h4014, 16'h4015, 16'h4016, 16'h4017 	:	val_out <= 16'hffff;
         16'h4018, 16'h4019, 16'h401a, 16'h401b, 16'h401c, 16'h401d, 16'h401e, 16'h401f 	:	val_out <= 16'hffff;
         16'h4020, 16'h4021, 16'h4022, 16'h4023, 16'h4024, 16'h4025, 16'h4026, 16'h4027 	:	val_out <= 16'hffff;
         16'h4028, 16'h4029, 16'h402a, 16'h402b, 16'h402c, 16'h402d, 16'h402e, 16'h402f 	:	val_out <= 16'hffff;
         16'h4030, 16'h4031, 16'h4032, 16'h4033, 16'h4034, 16'h4035, 16'h4036, 16'h4037 	:	val_out <= 16'hffff;
         16'h4038, 16'h4039, 16'h403a, 16'h403b, 16'h403c, 16'h403d, 16'h403e, 16'h403f 	:	val_out <= 16'hffff;
         16'h4040, 16'h4041, 16'h4042, 16'h4043, 16'h4044, 16'h4045, 16'h4046, 16'h4047 	:	val_out <= 16'hffff;
         16'h4048, 16'h4049, 16'h404a, 16'h404b, 16'h404c, 16'h404d, 16'h404e, 16'h404f 	:	val_out <= 16'hffff;
         16'h4050, 16'h4051, 16'h4052, 16'h4053, 16'h4054, 16'h4055, 16'h4056, 16'h4057 	:	val_out <= 16'hffff;
         16'h4058, 16'h4059, 16'h405a, 16'h405b, 16'h405c, 16'h405d, 16'h405e, 16'h405f 	:	val_out <= 16'hfffe;
         16'h4060, 16'h4061, 16'h4062, 16'h4063, 16'h4064, 16'h4065, 16'h4066, 16'h4067 	:	val_out <= 16'hfffe;
         16'h4068, 16'h4069, 16'h406a, 16'h406b, 16'h406c, 16'h406d, 16'h406e, 16'h406f 	:	val_out <= 16'hfffe;
         16'h4070, 16'h4071, 16'h4072, 16'h4073, 16'h4074, 16'h4075, 16'h4076, 16'h4077 	:	val_out <= 16'hfffe;
         16'h4078, 16'h4079, 16'h407a, 16'h407b, 16'h407c, 16'h407d, 16'h407e, 16'h407f 	:	val_out <= 16'hfffd;
         16'h4080, 16'h4081, 16'h4082, 16'h4083, 16'h4084, 16'h4085, 16'h4086, 16'h4087 	:	val_out <= 16'hfffd;
         16'h4088, 16'h4089, 16'h408a, 16'h408b, 16'h408c, 16'h408d, 16'h408e, 16'h408f 	:	val_out <= 16'hfffd;
         16'h4090, 16'h4091, 16'h4092, 16'h4093, 16'h4094, 16'h4095, 16'h4096, 16'h4097 	:	val_out <= 16'hfffc;
         16'h4098, 16'h4099, 16'h409a, 16'h409b, 16'h409c, 16'h409d, 16'h409e, 16'h409f 	:	val_out <= 16'hfffc;
         16'h40a0, 16'h40a1, 16'h40a2, 16'h40a3, 16'h40a4, 16'h40a5, 16'h40a6, 16'h40a7 	:	val_out <= 16'hfffc;
         16'h40a8, 16'h40a9, 16'h40aa, 16'h40ab, 16'h40ac, 16'h40ad, 16'h40ae, 16'h40af 	:	val_out <= 16'hfffb;
         16'h40b0, 16'h40b1, 16'h40b2, 16'h40b3, 16'h40b4, 16'h40b5, 16'h40b6, 16'h40b7 	:	val_out <= 16'hfffb;
         16'h40b8, 16'h40b9, 16'h40ba, 16'h40bb, 16'h40bc, 16'h40bd, 16'h40be, 16'h40bf 	:	val_out <= 16'hfffa;
         16'h40c0, 16'h40c1, 16'h40c2, 16'h40c3, 16'h40c4, 16'h40c5, 16'h40c6, 16'h40c7 	:	val_out <= 16'hfffa;
         16'h40c8, 16'h40c9, 16'h40ca, 16'h40cb, 16'h40cc, 16'h40cd, 16'h40ce, 16'h40cf 	:	val_out <= 16'hfff9;
         16'h40d0, 16'h40d1, 16'h40d2, 16'h40d3, 16'h40d4, 16'h40d5, 16'h40d6, 16'h40d7 	:	val_out <= 16'hfff9;
         16'h40d8, 16'h40d9, 16'h40da, 16'h40db, 16'h40dc, 16'h40dd, 16'h40de, 16'h40df 	:	val_out <= 16'hfff8;
         16'h40e0, 16'h40e1, 16'h40e2, 16'h40e3, 16'h40e4, 16'h40e5, 16'h40e6, 16'h40e7 	:	val_out <= 16'hfff8;
         16'h40e8, 16'h40e9, 16'h40ea, 16'h40eb, 16'h40ec, 16'h40ed, 16'h40ee, 16'h40ef 	:	val_out <= 16'hfff7;
         16'h40f0, 16'h40f1, 16'h40f2, 16'h40f3, 16'h40f4, 16'h40f5, 16'h40f6, 16'h40f7 	:	val_out <= 16'hfff7;
         16'h40f8, 16'h40f9, 16'h40fa, 16'h40fb, 16'h40fc, 16'h40fd, 16'h40fe, 16'h40ff 	:	val_out <= 16'hfff6;
         16'h4100, 16'h4101, 16'h4102, 16'h4103, 16'h4104, 16'h4105, 16'h4106, 16'h4107 	:	val_out <= 16'hfff6;
         16'h4108, 16'h4109, 16'h410a, 16'h410b, 16'h410c, 16'h410d, 16'h410e, 16'h410f 	:	val_out <= 16'hfff5;
         16'h4110, 16'h4111, 16'h4112, 16'h4113, 16'h4114, 16'h4115, 16'h4116, 16'h4117 	:	val_out <= 16'hfff4;
         16'h4118, 16'h4119, 16'h411a, 16'h411b, 16'h411c, 16'h411d, 16'h411e, 16'h411f 	:	val_out <= 16'hfff4;
         16'h4120, 16'h4121, 16'h4122, 16'h4123, 16'h4124, 16'h4125, 16'h4126, 16'h4127 	:	val_out <= 16'hfff3;
         16'h4128, 16'h4129, 16'h412a, 16'h412b, 16'h412c, 16'h412d, 16'h412e, 16'h412f 	:	val_out <= 16'hfff2;
         16'h4130, 16'h4131, 16'h4132, 16'h4133, 16'h4134, 16'h4135, 16'h4136, 16'h4137 	:	val_out <= 16'hfff2;
         16'h4138, 16'h4139, 16'h413a, 16'h413b, 16'h413c, 16'h413d, 16'h413e, 16'h413f 	:	val_out <= 16'hfff1;
         16'h4140, 16'h4141, 16'h4142, 16'h4143, 16'h4144, 16'h4145, 16'h4146, 16'h4147 	:	val_out <= 16'hfff0;
         16'h4148, 16'h4149, 16'h414a, 16'h414b, 16'h414c, 16'h414d, 16'h414e, 16'h414f 	:	val_out <= 16'hffef;
         16'h4150, 16'h4151, 16'h4152, 16'h4153, 16'h4154, 16'h4155, 16'h4156, 16'h4157 	:	val_out <= 16'hffee;
         16'h4158, 16'h4159, 16'h415a, 16'h415b, 16'h415c, 16'h415d, 16'h415e, 16'h415f 	:	val_out <= 16'hffee;
         16'h4160, 16'h4161, 16'h4162, 16'h4163, 16'h4164, 16'h4165, 16'h4166, 16'h4167 	:	val_out <= 16'hffed;
         16'h4168, 16'h4169, 16'h416a, 16'h416b, 16'h416c, 16'h416d, 16'h416e, 16'h416f 	:	val_out <= 16'hffec;
         16'h4170, 16'h4171, 16'h4172, 16'h4173, 16'h4174, 16'h4175, 16'h4176, 16'h4177 	:	val_out <= 16'hffeb;
         16'h4178, 16'h4179, 16'h417a, 16'h417b, 16'h417c, 16'h417d, 16'h417e, 16'h417f 	:	val_out <= 16'hffea;
         16'h4180, 16'h4181, 16'h4182, 16'h4183, 16'h4184, 16'h4185, 16'h4186, 16'h4187 	:	val_out <= 16'hffe9;
         16'h4188, 16'h4189, 16'h418a, 16'h418b, 16'h418c, 16'h418d, 16'h418e, 16'h418f 	:	val_out <= 16'hffe8;
         16'h4190, 16'h4191, 16'h4192, 16'h4193, 16'h4194, 16'h4195, 16'h4196, 16'h4197 	:	val_out <= 16'hffe7;
         16'h4198, 16'h4199, 16'h419a, 16'h419b, 16'h419c, 16'h419d, 16'h419e, 16'h419f 	:	val_out <= 16'hffe6;
         16'h41a0, 16'h41a1, 16'h41a2, 16'h41a3, 16'h41a4, 16'h41a5, 16'h41a6, 16'h41a7 	:	val_out <= 16'hffe5;
         16'h41a8, 16'h41a9, 16'h41aa, 16'h41ab, 16'h41ac, 16'h41ad, 16'h41ae, 16'h41af 	:	val_out <= 16'hffe4;
         16'h41b0, 16'h41b1, 16'h41b2, 16'h41b3, 16'h41b4, 16'h41b5, 16'h41b6, 16'h41b7 	:	val_out <= 16'hffe3;
         16'h41b8, 16'h41b9, 16'h41ba, 16'h41bb, 16'h41bc, 16'h41bd, 16'h41be, 16'h41bf 	:	val_out <= 16'hffe2;
         16'h41c0, 16'h41c1, 16'h41c2, 16'h41c3, 16'h41c4, 16'h41c5, 16'h41c6, 16'h41c7 	:	val_out <= 16'hffe1;
         16'h41c8, 16'h41c9, 16'h41ca, 16'h41cb, 16'h41cc, 16'h41cd, 16'h41ce, 16'h41cf 	:	val_out <= 16'hffe0;
         16'h41d0, 16'h41d1, 16'h41d2, 16'h41d3, 16'h41d4, 16'h41d5, 16'h41d6, 16'h41d7 	:	val_out <= 16'hffdf;
         16'h41d8, 16'h41d9, 16'h41da, 16'h41db, 16'h41dc, 16'h41dd, 16'h41de, 16'h41df 	:	val_out <= 16'hffde;
         16'h41e0, 16'h41e1, 16'h41e2, 16'h41e3, 16'h41e4, 16'h41e5, 16'h41e6, 16'h41e7 	:	val_out <= 16'hffdd;
         16'h41e8, 16'h41e9, 16'h41ea, 16'h41eb, 16'h41ec, 16'h41ed, 16'h41ee, 16'h41ef 	:	val_out <= 16'hffdc;
         16'h41f0, 16'h41f1, 16'h41f2, 16'h41f3, 16'h41f4, 16'h41f5, 16'h41f6, 16'h41f7 	:	val_out <= 16'hffda;
         16'h41f8, 16'h41f9, 16'h41fa, 16'h41fb, 16'h41fc, 16'h41fd, 16'h41fe, 16'h41ff 	:	val_out <= 16'hffd9;
         16'h4200, 16'h4201, 16'h4202, 16'h4203, 16'h4204, 16'h4205, 16'h4206, 16'h4207 	:	val_out <= 16'hffd8;
         16'h4208, 16'h4209, 16'h420a, 16'h420b, 16'h420c, 16'h420d, 16'h420e, 16'h420f 	:	val_out <= 16'hffd7;
         16'h4210, 16'h4211, 16'h4212, 16'h4213, 16'h4214, 16'h4215, 16'h4216, 16'h4217 	:	val_out <= 16'hffd6;
         16'h4218, 16'h4219, 16'h421a, 16'h421b, 16'h421c, 16'h421d, 16'h421e, 16'h421f 	:	val_out <= 16'hffd4;
         16'h4220, 16'h4221, 16'h4222, 16'h4223, 16'h4224, 16'h4225, 16'h4226, 16'h4227 	:	val_out <= 16'hffd3;
         16'h4228, 16'h4229, 16'h422a, 16'h422b, 16'h422c, 16'h422d, 16'h422e, 16'h422f 	:	val_out <= 16'hffd2;
         16'h4230, 16'h4231, 16'h4232, 16'h4233, 16'h4234, 16'h4235, 16'h4236, 16'h4237 	:	val_out <= 16'hffd0;
         16'h4238, 16'h4239, 16'h423a, 16'h423b, 16'h423c, 16'h423d, 16'h423e, 16'h423f 	:	val_out <= 16'hffcf;
         16'h4240, 16'h4241, 16'h4242, 16'h4243, 16'h4244, 16'h4245, 16'h4246, 16'h4247 	:	val_out <= 16'hffce;
         16'h4248, 16'h4249, 16'h424a, 16'h424b, 16'h424c, 16'h424d, 16'h424e, 16'h424f 	:	val_out <= 16'hffcc;
         16'h4250, 16'h4251, 16'h4252, 16'h4253, 16'h4254, 16'h4255, 16'h4256, 16'h4257 	:	val_out <= 16'hffcb;
         16'h4258, 16'h4259, 16'h425a, 16'h425b, 16'h425c, 16'h425d, 16'h425e, 16'h425f 	:	val_out <= 16'hffc9;
         16'h4260, 16'h4261, 16'h4262, 16'h4263, 16'h4264, 16'h4265, 16'h4266, 16'h4267 	:	val_out <= 16'hffc8;
         16'h4268, 16'h4269, 16'h426a, 16'h426b, 16'h426c, 16'h426d, 16'h426e, 16'h426f 	:	val_out <= 16'hffc6;
         16'h4270, 16'h4271, 16'h4272, 16'h4273, 16'h4274, 16'h4275, 16'h4276, 16'h4277 	:	val_out <= 16'hffc5;
         16'h4278, 16'h4279, 16'h427a, 16'h427b, 16'h427c, 16'h427d, 16'h427e, 16'h427f 	:	val_out <= 16'hffc3;
         16'h4280, 16'h4281, 16'h4282, 16'h4283, 16'h4284, 16'h4285, 16'h4286, 16'h4287 	:	val_out <= 16'hffc2;
         16'h4288, 16'h4289, 16'h428a, 16'h428b, 16'h428c, 16'h428d, 16'h428e, 16'h428f 	:	val_out <= 16'hffc0;
         16'h4290, 16'h4291, 16'h4292, 16'h4293, 16'h4294, 16'h4295, 16'h4296, 16'h4297 	:	val_out <= 16'hffbf;
         16'h4298, 16'h4299, 16'h429a, 16'h429b, 16'h429c, 16'h429d, 16'h429e, 16'h429f 	:	val_out <= 16'hffbd;
         16'h42a0, 16'h42a1, 16'h42a2, 16'h42a3, 16'h42a4, 16'h42a5, 16'h42a6, 16'h42a7 	:	val_out <= 16'hffbc;
         16'h42a8, 16'h42a9, 16'h42aa, 16'h42ab, 16'h42ac, 16'h42ad, 16'h42ae, 16'h42af 	:	val_out <= 16'hffba;
         16'h42b0, 16'h42b1, 16'h42b2, 16'h42b3, 16'h42b4, 16'h42b5, 16'h42b6, 16'h42b7 	:	val_out <= 16'hffb8;
         16'h42b8, 16'h42b9, 16'h42ba, 16'h42bb, 16'h42bc, 16'h42bd, 16'h42be, 16'h42bf 	:	val_out <= 16'hffb7;
         16'h42c0, 16'h42c1, 16'h42c2, 16'h42c3, 16'h42c4, 16'h42c5, 16'h42c6, 16'h42c7 	:	val_out <= 16'hffb5;
         16'h42c8, 16'h42c9, 16'h42ca, 16'h42cb, 16'h42cc, 16'h42cd, 16'h42ce, 16'h42cf 	:	val_out <= 16'hffb3;
         16'h42d0, 16'h42d1, 16'h42d2, 16'h42d3, 16'h42d4, 16'h42d5, 16'h42d6, 16'h42d7 	:	val_out <= 16'hffb1;
         16'h42d8, 16'h42d9, 16'h42da, 16'h42db, 16'h42dc, 16'h42dd, 16'h42de, 16'h42df 	:	val_out <= 16'hffb0;
         16'h42e0, 16'h42e1, 16'h42e2, 16'h42e3, 16'h42e4, 16'h42e5, 16'h42e6, 16'h42e7 	:	val_out <= 16'hffae;
         16'h42e8, 16'h42e9, 16'h42ea, 16'h42eb, 16'h42ec, 16'h42ed, 16'h42ee, 16'h42ef 	:	val_out <= 16'hffac;
         16'h42f0, 16'h42f1, 16'h42f2, 16'h42f3, 16'h42f4, 16'h42f5, 16'h42f6, 16'h42f7 	:	val_out <= 16'hffaa;
         16'h42f8, 16'h42f9, 16'h42fa, 16'h42fb, 16'h42fc, 16'h42fd, 16'h42fe, 16'h42ff 	:	val_out <= 16'hffa9;
         16'h4300, 16'h4301, 16'h4302, 16'h4303, 16'h4304, 16'h4305, 16'h4306, 16'h4307 	:	val_out <= 16'hffa7;
         16'h4308, 16'h4309, 16'h430a, 16'h430b, 16'h430c, 16'h430d, 16'h430e, 16'h430f 	:	val_out <= 16'hffa5;
         16'h4310, 16'h4311, 16'h4312, 16'h4313, 16'h4314, 16'h4315, 16'h4316, 16'h4317 	:	val_out <= 16'hffa3;
         16'h4318, 16'h4319, 16'h431a, 16'h431b, 16'h431c, 16'h431d, 16'h431e, 16'h431f 	:	val_out <= 16'hffa1;
         16'h4320, 16'h4321, 16'h4322, 16'h4323, 16'h4324, 16'h4325, 16'h4326, 16'h4327 	:	val_out <= 16'hff9f;
         16'h4328, 16'h4329, 16'h432a, 16'h432b, 16'h432c, 16'h432d, 16'h432e, 16'h432f 	:	val_out <= 16'hff9d;
         16'h4330, 16'h4331, 16'h4332, 16'h4333, 16'h4334, 16'h4335, 16'h4336, 16'h4337 	:	val_out <= 16'hff9b;
         16'h4338, 16'h4339, 16'h433a, 16'h433b, 16'h433c, 16'h433d, 16'h433e, 16'h433f 	:	val_out <= 16'hff99;
         16'h4340, 16'h4341, 16'h4342, 16'h4343, 16'h4344, 16'h4345, 16'h4346, 16'h4347 	:	val_out <= 16'hff97;
         16'h4348, 16'h4349, 16'h434a, 16'h434b, 16'h434c, 16'h434d, 16'h434e, 16'h434f 	:	val_out <= 16'hff95;
         16'h4350, 16'h4351, 16'h4352, 16'h4353, 16'h4354, 16'h4355, 16'h4356, 16'h4357 	:	val_out <= 16'hff93;
         16'h4358, 16'h4359, 16'h435a, 16'h435b, 16'h435c, 16'h435d, 16'h435e, 16'h435f 	:	val_out <= 16'hff91;
         16'h4360, 16'h4361, 16'h4362, 16'h4363, 16'h4364, 16'h4365, 16'h4366, 16'h4367 	:	val_out <= 16'hff8f;
         16'h4368, 16'h4369, 16'h436a, 16'h436b, 16'h436c, 16'h436d, 16'h436e, 16'h436f 	:	val_out <= 16'hff8d;
         16'h4370, 16'h4371, 16'h4372, 16'h4373, 16'h4374, 16'h4375, 16'h4376, 16'h4377 	:	val_out <= 16'hff8b;
         16'h4378, 16'h4379, 16'h437a, 16'h437b, 16'h437c, 16'h437d, 16'h437e, 16'h437f 	:	val_out <= 16'hff89;
         16'h4380, 16'h4381, 16'h4382, 16'h4383, 16'h4384, 16'h4385, 16'h4386, 16'h4387 	:	val_out <= 16'hff87;
         16'h4388, 16'h4389, 16'h438a, 16'h438b, 16'h438c, 16'h438d, 16'h438e, 16'h438f 	:	val_out <= 16'hff85;
         16'h4390, 16'h4391, 16'h4392, 16'h4393, 16'h4394, 16'h4395, 16'h4396, 16'h4397 	:	val_out <= 16'hff82;
         16'h4398, 16'h4399, 16'h439a, 16'h439b, 16'h439c, 16'h439d, 16'h439e, 16'h439f 	:	val_out <= 16'hff80;
         16'h43a0, 16'h43a1, 16'h43a2, 16'h43a3, 16'h43a4, 16'h43a5, 16'h43a6, 16'h43a7 	:	val_out <= 16'hff7e;
         16'h43a8, 16'h43a9, 16'h43aa, 16'h43ab, 16'h43ac, 16'h43ad, 16'h43ae, 16'h43af 	:	val_out <= 16'hff7c;
         16'h43b0, 16'h43b1, 16'h43b2, 16'h43b3, 16'h43b4, 16'h43b5, 16'h43b6, 16'h43b7 	:	val_out <= 16'hff79;
         16'h43b8, 16'h43b9, 16'h43ba, 16'h43bb, 16'h43bc, 16'h43bd, 16'h43be, 16'h43bf 	:	val_out <= 16'hff77;
         16'h43c0, 16'h43c1, 16'h43c2, 16'h43c3, 16'h43c4, 16'h43c5, 16'h43c6, 16'h43c7 	:	val_out <= 16'hff75;
         16'h43c8, 16'h43c9, 16'h43ca, 16'h43cb, 16'h43cc, 16'h43cd, 16'h43ce, 16'h43cf 	:	val_out <= 16'hff72;
         16'h43d0, 16'h43d1, 16'h43d2, 16'h43d3, 16'h43d4, 16'h43d5, 16'h43d6, 16'h43d7 	:	val_out <= 16'hff70;
         16'h43d8, 16'h43d9, 16'h43da, 16'h43db, 16'h43dc, 16'h43dd, 16'h43de, 16'h43df 	:	val_out <= 16'hff6e;
         16'h43e0, 16'h43e1, 16'h43e2, 16'h43e3, 16'h43e4, 16'h43e5, 16'h43e6, 16'h43e7 	:	val_out <= 16'hff6b;
         16'h43e8, 16'h43e9, 16'h43ea, 16'h43eb, 16'h43ec, 16'h43ed, 16'h43ee, 16'h43ef 	:	val_out <= 16'hff69;
         16'h43f0, 16'h43f1, 16'h43f2, 16'h43f3, 16'h43f4, 16'h43f5, 16'h43f6, 16'h43f7 	:	val_out <= 16'hff67;
         16'h43f8, 16'h43f9, 16'h43fa, 16'h43fb, 16'h43fc, 16'h43fd, 16'h43fe, 16'h43ff 	:	val_out <= 16'hff64;
         16'h4400, 16'h4401, 16'h4402, 16'h4403, 16'h4404, 16'h4405, 16'h4406, 16'h4407 	:	val_out <= 16'hff62;
         16'h4408, 16'h4409, 16'h440a, 16'h440b, 16'h440c, 16'h440d, 16'h440e, 16'h440f 	:	val_out <= 16'hff5f;
         16'h4410, 16'h4411, 16'h4412, 16'h4413, 16'h4414, 16'h4415, 16'h4416, 16'h4417 	:	val_out <= 16'hff5d;
         16'h4418, 16'h4419, 16'h441a, 16'h441b, 16'h441c, 16'h441d, 16'h441e, 16'h441f 	:	val_out <= 16'hff5a;
         16'h4420, 16'h4421, 16'h4422, 16'h4423, 16'h4424, 16'h4425, 16'h4426, 16'h4427 	:	val_out <= 16'hff58;
         16'h4428, 16'h4429, 16'h442a, 16'h442b, 16'h442c, 16'h442d, 16'h442e, 16'h442f 	:	val_out <= 16'hff55;
         16'h4430, 16'h4431, 16'h4432, 16'h4433, 16'h4434, 16'h4435, 16'h4436, 16'h4437 	:	val_out <= 16'hff53;
         16'h4438, 16'h4439, 16'h443a, 16'h443b, 16'h443c, 16'h443d, 16'h443e, 16'h443f 	:	val_out <= 16'hff50;
         16'h4440, 16'h4441, 16'h4442, 16'h4443, 16'h4444, 16'h4445, 16'h4446, 16'h4447 	:	val_out <= 16'hff4d;
         16'h4448, 16'h4449, 16'h444a, 16'h444b, 16'h444c, 16'h444d, 16'h444e, 16'h444f 	:	val_out <= 16'hff4b;
         16'h4450, 16'h4451, 16'h4452, 16'h4453, 16'h4454, 16'h4455, 16'h4456, 16'h4457 	:	val_out <= 16'hff48;
         16'h4458, 16'h4459, 16'h445a, 16'h445b, 16'h445c, 16'h445d, 16'h445e, 16'h445f 	:	val_out <= 16'hff45;
         16'h4460, 16'h4461, 16'h4462, 16'h4463, 16'h4464, 16'h4465, 16'h4466, 16'h4467 	:	val_out <= 16'hff43;
         16'h4468, 16'h4469, 16'h446a, 16'h446b, 16'h446c, 16'h446d, 16'h446e, 16'h446f 	:	val_out <= 16'hff40;
         16'h4470, 16'h4471, 16'h4472, 16'h4473, 16'h4474, 16'h4475, 16'h4476, 16'h4477 	:	val_out <= 16'hff3d;
         16'h4478, 16'h4479, 16'h447a, 16'h447b, 16'h447c, 16'h447d, 16'h447e, 16'h447f 	:	val_out <= 16'hff3b;
         16'h4480, 16'h4481, 16'h4482, 16'h4483, 16'h4484, 16'h4485, 16'h4486, 16'h4487 	:	val_out <= 16'hff38;
         16'h4488, 16'h4489, 16'h448a, 16'h448b, 16'h448c, 16'h448d, 16'h448e, 16'h448f 	:	val_out <= 16'hff35;
         16'h4490, 16'h4491, 16'h4492, 16'h4493, 16'h4494, 16'h4495, 16'h4496, 16'h4497 	:	val_out <= 16'hff32;
         16'h4498, 16'h4499, 16'h449a, 16'h449b, 16'h449c, 16'h449d, 16'h449e, 16'h449f 	:	val_out <= 16'hff2f;
         16'h44a0, 16'h44a1, 16'h44a2, 16'h44a3, 16'h44a4, 16'h44a5, 16'h44a6, 16'h44a7 	:	val_out <= 16'hff2d;
         16'h44a8, 16'h44a9, 16'h44aa, 16'h44ab, 16'h44ac, 16'h44ad, 16'h44ae, 16'h44af 	:	val_out <= 16'hff2a;
         16'h44b0, 16'h44b1, 16'h44b2, 16'h44b3, 16'h44b4, 16'h44b5, 16'h44b6, 16'h44b7 	:	val_out <= 16'hff27;
         16'h44b8, 16'h44b9, 16'h44ba, 16'h44bb, 16'h44bc, 16'h44bd, 16'h44be, 16'h44bf 	:	val_out <= 16'hff24;
         16'h44c0, 16'h44c1, 16'h44c2, 16'h44c3, 16'h44c4, 16'h44c5, 16'h44c6, 16'h44c7 	:	val_out <= 16'hff21;
         16'h44c8, 16'h44c9, 16'h44ca, 16'h44cb, 16'h44cc, 16'h44cd, 16'h44ce, 16'h44cf 	:	val_out <= 16'hff1e;
         16'h44d0, 16'h44d1, 16'h44d2, 16'h44d3, 16'h44d4, 16'h44d5, 16'h44d6, 16'h44d7 	:	val_out <= 16'hff1b;
         16'h44d8, 16'h44d9, 16'h44da, 16'h44db, 16'h44dc, 16'h44dd, 16'h44de, 16'h44df 	:	val_out <= 16'hff18;
         16'h44e0, 16'h44e1, 16'h44e2, 16'h44e3, 16'h44e4, 16'h44e5, 16'h44e6, 16'h44e7 	:	val_out <= 16'hff15;
         16'h44e8, 16'h44e9, 16'h44ea, 16'h44eb, 16'h44ec, 16'h44ed, 16'h44ee, 16'h44ef 	:	val_out <= 16'hff12;
         16'h44f0, 16'h44f1, 16'h44f2, 16'h44f3, 16'h44f4, 16'h44f5, 16'h44f6, 16'h44f7 	:	val_out <= 16'hff0f;
         16'h44f8, 16'h44f9, 16'h44fa, 16'h44fb, 16'h44fc, 16'h44fd, 16'h44fe, 16'h44ff 	:	val_out <= 16'hff0c;
         16'h4500, 16'h4501, 16'h4502, 16'h4503, 16'h4504, 16'h4505, 16'h4506, 16'h4507 	:	val_out <= 16'hff09;
         16'h4508, 16'h4509, 16'h450a, 16'h450b, 16'h450c, 16'h450d, 16'h450e, 16'h450f 	:	val_out <= 16'hff06;
         16'h4510, 16'h4511, 16'h4512, 16'h4513, 16'h4514, 16'h4515, 16'h4516, 16'h4517 	:	val_out <= 16'hff03;
         16'h4518, 16'h4519, 16'h451a, 16'h451b, 16'h451c, 16'h451d, 16'h451e, 16'h451f 	:	val_out <= 16'hff00;
         16'h4520, 16'h4521, 16'h4522, 16'h4523, 16'h4524, 16'h4525, 16'h4526, 16'h4527 	:	val_out <= 16'hfefd;
         16'h4528, 16'h4529, 16'h452a, 16'h452b, 16'h452c, 16'h452d, 16'h452e, 16'h452f 	:	val_out <= 16'hfef9;
         16'h4530, 16'h4531, 16'h4532, 16'h4533, 16'h4534, 16'h4535, 16'h4536, 16'h4537 	:	val_out <= 16'hfef6;
         16'h4538, 16'h4539, 16'h453a, 16'h453b, 16'h453c, 16'h453d, 16'h453e, 16'h453f 	:	val_out <= 16'hfef3;
         16'h4540, 16'h4541, 16'h4542, 16'h4543, 16'h4544, 16'h4545, 16'h4546, 16'h4547 	:	val_out <= 16'hfef0;
         16'h4548, 16'h4549, 16'h454a, 16'h454b, 16'h454c, 16'h454d, 16'h454e, 16'h454f 	:	val_out <= 16'hfeed;
         16'h4550, 16'h4551, 16'h4552, 16'h4553, 16'h4554, 16'h4555, 16'h4556, 16'h4557 	:	val_out <= 16'hfee9;
         16'h4558, 16'h4559, 16'h455a, 16'h455b, 16'h455c, 16'h455d, 16'h455e, 16'h455f 	:	val_out <= 16'hfee6;
         16'h4560, 16'h4561, 16'h4562, 16'h4563, 16'h4564, 16'h4565, 16'h4566, 16'h4567 	:	val_out <= 16'hfee3;
         16'h4568, 16'h4569, 16'h456a, 16'h456b, 16'h456c, 16'h456d, 16'h456e, 16'h456f 	:	val_out <= 16'hfedf;
         16'h4570, 16'h4571, 16'h4572, 16'h4573, 16'h4574, 16'h4575, 16'h4576, 16'h4577 	:	val_out <= 16'hfedc;
         16'h4578, 16'h4579, 16'h457a, 16'h457b, 16'h457c, 16'h457d, 16'h457e, 16'h457f 	:	val_out <= 16'hfed9;
         16'h4580, 16'h4581, 16'h4582, 16'h4583, 16'h4584, 16'h4585, 16'h4586, 16'h4587 	:	val_out <= 16'hfed5;
         16'h4588, 16'h4589, 16'h458a, 16'h458b, 16'h458c, 16'h458d, 16'h458e, 16'h458f 	:	val_out <= 16'hfed2;
         16'h4590, 16'h4591, 16'h4592, 16'h4593, 16'h4594, 16'h4595, 16'h4596, 16'h4597 	:	val_out <= 16'hfecf;
         16'h4598, 16'h4599, 16'h459a, 16'h459b, 16'h459c, 16'h459d, 16'h459e, 16'h459f 	:	val_out <= 16'hfecb;
         16'h45a0, 16'h45a1, 16'h45a2, 16'h45a3, 16'h45a4, 16'h45a5, 16'h45a6, 16'h45a7 	:	val_out <= 16'hfec8;
         16'h45a8, 16'h45a9, 16'h45aa, 16'h45ab, 16'h45ac, 16'h45ad, 16'h45ae, 16'h45af 	:	val_out <= 16'hfec4;
         16'h45b0, 16'h45b1, 16'h45b2, 16'h45b3, 16'h45b4, 16'h45b5, 16'h45b6, 16'h45b7 	:	val_out <= 16'hfec1;
         16'h45b8, 16'h45b9, 16'h45ba, 16'h45bb, 16'h45bc, 16'h45bd, 16'h45be, 16'h45bf 	:	val_out <= 16'hfebd;
         16'h45c0, 16'h45c1, 16'h45c2, 16'h45c3, 16'h45c4, 16'h45c5, 16'h45c6, 16'h45c7 	:	val_out <= 16'hfeba;
         16'h45c8, 16'h45c9, 16'h45ca, 16'h45cb, 16'h45cc, 16'h45cd, 16'h45ce, 16'h45cf 	:	val_out <= 16'hfeb6;
         16'h45d0, 16'h45d1, 16'h45d2, 16'h45d3, 16'h45d4, 16'h45d5, 16'h45d6, 16'h45d7 	:	val_out <= 16'hfeb3;
         16'h45d8, 16'h45d9, 16'h45da, 16'h45db, 16'h45dc, 16'h45dd, 16'h45de, 16'h45df 	:	val_out <= 16'hfeaf;
         16'h45e0, 16'h45e1, 16'h45e2, 16'h45e3, 16'h45e4, 16'h45e5, 16'h45e6, 16'h45e7 	:	val_out <= 16'hfeab;
         16'h45e8, 16'h45e9, 16'h45ea, 16'h45eb, 16'h45ec, 16'h45ed, 16'h45ee, 16'h45ef 	:	val_out <= 16'hfea8;
         16'h45f0, 16'h45f1, 16'h45f2, 16'h45f3, 16'h45f4, 16'h45f5, 16'h45f6, 16'h45f7 	:	val_out <= 16'hfea4;
         16'h45f8, 16'h45f9, 16'h45fa, 16'h45fb, 16'h45fc, 16'h45fd, 16'h45fe, 16'h45ff 	:	val_out <= 16'hfea1;
         16'h4600, 16'h4601, 16'h4602, 16'h4603, 16'h4604, 16'h4605, 16'h4606, 16'h4607 	:	val_out <= 16'hfe9d;
         16'h4608, 16'h4609, 16'h460a, 16'h460b, 16'h460c, 16'h460d, 16'h460e, 16'h460f 	:	val_out <= 16'hfe99;
         16'h4610, 16'h4611, 16'h4612, 16'h4613, 16'h4614, 16'h4615, 16'h4616, 16'h4617 	:	val_out <= 16'hfe95;
         16'h4618, 16'h4619, 16'h461a, 16'h461b, 16'h461c, 16'h461d, 16'h461e, 16'h461f 	:	val_out <= 16'hfe92;
         16'h4620, 16'h4621, 16'h4622, 16'h4623, 16'h4624, 16'h4625, 16'h4626, 16'h4627 	:	val_out <= 16'hfe8e;
         16'h4628, 16'h4629, 16'h462a, 16'h462b, 16'h462c, 16'h462d, 16'h462e, 16'h462f 	:	val_out <= 16'hfe8a;
         16'h4630, 16'h4631, 16'h4632, 16'h4633, 16'h4634, 16'h4635, 16'h4636, 16'h4637 	:	val_out <= 16'hfe86;
         16'h4638, 16'h4639, 16'h463a, 16'h463b, 16'h463c, 16'h463d, 16'h463e, 16'h463f 	:	val_out <= 16'hfe83;
         16'h4640, 16'h4641, 16'h4642, 16'h4643, 16'h4644, 16'h4645, 16'h4646, 16'h4647 	:	val_out <= 16'hfe7f;
         16'h4648, 16'h4649, 16'h464a, 16'h464b, 16'h464c, 16'h464d, 16'h464e, 16'h464f 	:	val_out <= 16'hfe7b;
         16'h4650, 16'h4651, 16'h4652, 16'h4653, 16'h4654, 16'h4655, 16'h4656, 16'h4657 	:	val_out <= 16'hfe77;
         16'h4658, 16'h4659, 16'h465a, 16'h465b, 16'h465c, 16'h465d, 16'h465e, 16'h465f 	:	val_out <= 16'hfe73;
         16'h4660, 16'h4661, 16'h4662, 16'h4663, 16'h4664, 16'h4665, 16'h4666, 16'h4667 	:	val_out <= 16'hfe6f;
         16'h4668, 16'h4669, 16'h466a, 16'h466b, 16'h466c, 16'h466d, 16'h466e, 16'h466f 	:	val_out <= 16'hfe6b;
         16'h4670, 16'h4671, 16'h4672, 16'h4673, 16'h4674, 16'h4675, 16'h4676, 16'h4677 	:	val_out <= 16'hfe67;
         16'h4678, 16'h4679, 16'h467a, 16'h467b, 16'h467c, 16'h467d, 16'h467e, 16'h467f 	:	val_out <= 16'hfe63;
         16'h4680, 16'h4681, 16'h4682, 16'h4683, 16'h4684, 16'h4685, 16'h4686, 16'h4687 	:	val_out <= 16'hfe5f;
         16'h4688, 16'h4689, 16'h468a, 16'h468b, 16'h468c, 16'h468d, 16'h468e, 16'h468f 	:	val_out <= 16'hfe5b;
         16'h4690, 16'h4691, 16'h4692, 16'h4693, 16'h4694, 16'h4695, 16'h4696, 16'h4697 	:	val_out <= 16'hfe57;
         16'h4698, 16'h4699, 16'h469a, 16'h469b, 16'h469c, 16'h469d, 16'h469e, 16'h469f 	:	val_out <= 16'hfe53;
         16'h46a0, 16'h46a1, 16'h46a2, 16'h46a3, 16'h46a4, 16'h46a5, 16'h46a6, 16'h46a7 	:	val_out <= 16'hfe4f;
         16'h46a8, 16'h46a9, 16'h46aa, 16'h46ab, 16'h46ac, 16'h46ad, 16'h46ae, 16'h46af 	:	val_out <= 16'hfe4b;
         16'h46b0, 16'h46b1, 16'h46b2, 16'h46b3, 16'h46b4, 16'h46b5, 16'h46b6, 16'h46b7 	:	val_out <= 16'hfe47;
         16'h46b8, 16'h46b9, 16'h46ba, 16'h46bb, 16'h46bc, 16'h46bd, 16'h46be, 16'h46bf 	:	val_out <= 16'hfe43;
         16'h46c0, 16'h46c1, 16'h46c2, 16'h46c3, 16'h46c4, 16'h46c5, 16'h46c6, 16'h46c7 	:	val_out <= 16'hfe3f;
         16'h46c8, 16'h46c9, 16'h46ca, 16'h46cb, 16'h46cc, 16'h46cd, 16'h46ce, 16'h46cf 	:	val_out <= 16'hfe3b;
         16'h46d0, 16'h46d1, 16'h46d2, 16'h46d3, 16'h46d4, 16'h46d5, 16'h46d6, 16'h46d7 	:	val_out <= 16'hfe37;
         16'h46d8, 16'h46d9, 16'h46da, 16'h46db, 16'h46dc, 16'h46dd, 16'h46de, 16'h46df 	:	val_out <= 16'hfe32;
         16'h46e0, 16'h46e1, 16'h46e2, 16'h46e3, 16'h46e4, 16'h46e5, 16'h46e6, 16'h46e7 	:	val_out <= 16'hfe2e;
         16'h46e8, 16'h46e9, 16'h46ea, 16'h46eb, 16'h46ec, 16'h46ed, 16'h46ee, 16'h46ef 	:	val_out <= 16'hfe2a;
         16'h46f0, 16'h46f1, 16'h46f2, 16'h46f3, 16'h46f4, 16'h46f5, 16'h46f6, 16'h46f7 	:	val_out <= 16'hfe26;
         16'h46f8, 16'h46f9, 16'h46fa, 16'h46fb, 16'h46fc, 16'h46fd, 16'h46fe, 16'h46ff 	:	val_out <= 16'hfe21;
         16'h4700, 16'h4701, 16'h4702, 16'h4703, 16'h4704, 16'h4705, 16'h4706, 16'h4707 	:	val_out <= 16'hfe1d;
         16'h4708, 16'h4709, 16'h470a, 16'h470b, 16'h470c, 16'h470d, 16'h470e, 16'h470f 	:	val_out <= 16'hfe19;
         16'h4710, 16'h4711, 16'h4712, 16'h4713, 16'h4714, 16'h4715, 16'h4716, 16'h4717 	:	val_out <= 16'hfe14;
         16'h4718, 16'h4719, 16'h471a, 16'h471b, 16'h471c, 16'h471d, 16'h471e, 16'h471f 	:	val_out <= 16'hfe10;
         16'h4720, 16'h4721, 16'h4722, 16'h4723, 16'h4724, 16'h4725, 16'h4726, 16'h4727 	:	val_out <= 16'hfe0c;
         16'h4728, 16'h4729, 16'h472a, 16'h472b, 16'h472c, 16'h472d, 16'h472e, 16'h472f 	:	val_out <= 16'hfe07;
         16'h4730, 16'h4731, 16'h4732, 16'h4733, 16'h4734, 16'h4735, 16'h4736, 16'h4737 	:	val_out <= 16'hfe03;
         16'h4738, 16'h4739, 16'h473a, 16'h473b, 16'h473c, 16'h473d, 16'h473e, 16'h473f 	:	val_out <= 16'hfdff;
         16'h4740, 16'h4741, 16'h4742, 16'h4743, 16'h4744, 16'h4745, 16'h4746, 16'h4747 	:	val_out <= 16'hfdfa;
         16'h4748, 16'h4749, 16'h474a, 16'h474b, 16'h474c, 16'h474d, 16'h474e, 16'h474f 	:	val_out <= 16'hfdf6;
         16'h4750, 16'h4751, 16'h4752, 16'h4753, 16'h4754, 16'h4755, 16'h4756, 16'h4757 	:	val_out <= 16'hfdf1;
         16'h4758, 16'h4759, 16'h475a, 16'h475b, 16'h475c, 16'h475d, 16'h475e, 16'h475f 	:	val_out <= 16'hfded;
         16'h4760, 16'h4761, 16'h4762, 16'h4763, 16'h4764, 16'h4765, 16'h4766, 16'h4767 	:	val_out <= 16'hfde8;
         16'h4768, 16'h4769, 16'h476a, 16'h476b, 16'h476c, 16'h476d, 16'h476e, 16'h476f 	:	val_out <= 16'hfde4;
         16'h4770, 16'h4771, 16'h4772, 16'h4773, 16'h4774, 16'h4775, 16'h4776, 16'h4777 	:	val_out <= 16'hfddf;
         16'h4778, 16'h4779, 16'h477a, 16'h477b, 16'h477c, 16'h477d, 16'h477e, 16'h477f 	:	val_out <= 16'hfdda;
         16'h4780, 16'h4781, 16'h4782, 16'h4783, 16'h4784, 16'h4785, 16'h4786, 16'h4787 	:	val_out <= 16'hfdd6;
         16'h4788, 16'h4789, 16'h478a, 16'h478b, 16'h478c, 16'h478d, 16'h478e, 16'h478f 	:	val_out <= 16'hfdd1;
         16'h4790, 16'h4791, 16'h4792, 16'h4793, 16'h4794, 16'h4795, 16'h4796, 16'h4797 	:	val_out <= 16'hfdcd;
         16'h4798, 16'h4799, 16'h479a, 16'h479b, 16'h479c, 16'h479d, 16'h479e, 16'h479f 	:	val_out <= 16'hfdc8;
         16'h47a0, 16'h47a1, 16'h47a2, 16'h47a3, 16'h47a4, 16'h47a5, 16'h47a6, 16'h47a7 	:	val_out <= 16'hfdc3;
         16'h47a8, 16'h47a9, 16'h47aa, 16'h47ab, 16'h47ac, 16'h47ad, 16'h47ae, 16'h47af 	:	val_out <= 16'hfdbf;
         16'h47b0, 16'h47b1, 16'h47b2, 16'h47b3, 16'h47b4, 16'h47b5, 16'h47b6, 16'h47b7 	:	val_out <= 16'hfdba;
         16'h47b8, 16'h47b9, 16'h47ba, 16'h47bb, 16'h47bc, 16'h47bd, 16'h47be, 16'h47bf 	:	val_out <= 16'hfdb5;
         16'h47c0, 16'h47c1, 16'h47c2, 16'h47c3, 16'h47c4, 16'h47c5, 16'h47c6, 16'h47c7 	:	val_out <= 16'hfdb0;
         16'h47c8, 16'h47c9, 16'h47ca, 16'h47cb, 16'h47cc, 16'h47cd, 16'h47ce, 16'h47cf 	:	val_out <= 16'hfdac;
         16'h47d0, 16'h47d1, 16'h47d2, 16'h47d3, 16'h47d4, 16'h47d5, 16'h47d6, 16'h47d7 	:	val_out <= 16'hfda7;
         16'h47d8, 16'h47d9, 16'h47da, 16'h47db, 16'h47dc, 16'h47dd, 16'h47de, 16'h47df 	:	val_out <= 16'hfda2;
         16'h47e0, 16'h47e1, 16'h47e2, 16'h47e3, 16'h47e4, 16'h47e5, 16'h47e6, 16'h47e7 	:	val_out <= 16'hfd9d;
         16'h47e8, 16'h47e9, 16'h47ea, 16'h47eb, 16'h47ec, 16'h47ed, 16'h47ee, 16'h47ef 	:	val_out <= 16'hfd98;
         16'h47f0, 16'h47f1, 16'h47f2, 16'h47f3, 16'h47f4, 16'h47f5, 16'h47f6, 16'h47f7 	:	val_out <= 16'hfd94;
         16'h47f8, 16'h47f9, 16'h47fa, 16'h47fb, 16'h47fc, 16'h47fd, 16'h47fe, 16'h47ff 	:	val_out <= 16'hfd8f;
         16'h4800, 16'h4801, 16'h4802, 16'h4803, 16'h4804, 16'h4805, 16'h4806, 16'h4807 	:	val_out <= 16'hfd8a;
         16'h4808, 16'h4809, 16'h480a, 16'h480b, 16'h480c, 16'h480d, 16'h480e, 16'h480f 	:	val_out <= 16'hfd85;
         16'h4810, 16'h4811, 16'h4812, 16'h4813, 16'h4814, 16'h4815, 16'h4816, 16'h4817 	:	val_out <= 16'hfd80;
         16'h4818, 16'h4819, 16'h481a, 16'h481b, 16'h481c, 16'h481d, 16'h481e, 16'h481f 	:	val_out <= 16'hfd7b;
         16'h4820, 16'h4821, 16'h4822, 16'h4823, 16'h4824, 16'h4825, 16'h4826, 16'h4827 	:	val_out <= 16'hfd76;
         16'h4828, 16'h4829, 16'h482a, 16'h482b, 16'h482c, 16'h482d, 16'h482e, 16'h482f 	:	val_out <= 16'hfd71;
         16'h4830, 16'h4831, 16'h4832, 16'h4833, 16'h4834, 16'h4835, 16'h4836, 16'h4837 	:	val_out <= 16'hfd6c;
         16'h4838, 16'h4839, 16'h483a, 16'h483b, 16'h483c, 16'h483d, 16'h483e, 16'h483f 	:	val_out <= 16'hfd67;
         16'h4840, 16'h4841, 16'h4842, 16'h4843, 16'h4844, 16'h4845, 16'h4846, 16'h4847 	:	val_out <= 16'hfd62;
         16'h4848, 16'h4849, 16'h484a, 16'h484b, 16'h484c, 16'h484d, 16'h484e, 16'h484f 	:	val_out <= 16'hfd5d;
         16'h4850, 16'h4851, 16'h4852, 16'h4853, 16'h4854, 16'h4855, 16'h4856, 16'h4857 	:	val_out <= 16'hfd58;
         16'h4858, 16'h4859, 16'h485a, 16'h485b, 16'h485c, 16'h485d, 16'h485e, 16'h485f 	:	val_out <= 16'hfd53;
         16'h4860, 16'h4861, 16'h4862, 16'h4863, 16'h4864, 16'h4865, 16'h4866, 16'h4867 	:	val_out <= 16'hfd4e;
         16'h4868, 16'h4869, 16'h486a, 16'h486b, 16'h486c, 16'h486d, 16'h486e, 16'h486f 	:	val_out <= 16'hfd49;
         16'h4870, 16'h4871, 16'h4872, 16'h4873, 16'h4874, 16'h4875, 16'h4876, 16'h4877 	:	val_out <= 16'hfd43;
         16'h4878, 16'h4879, 16'h487a, 16'h487b, 16'h487c, 16'h487d, 16'h487e, 16'h487f 	:	val_out <= 16'hfd3e;
         16'h4880, 16'h4881, 16'h4882, 16'h4883, 16'h4884, 16'h4885, 16'h4886, 16'h4887 	:	val_out <= 16'hfd39;
         16'h4888, 16'h4889, 16'h488a, 16'h488b, 16'h488c, 16'h488d, 16'h488e, 16'h488f 	:	val_out <= 16'hfd34;
         16'h4890, 16'h4891, 16'h4892, 16'h4893, 16'h4894, 16'h4895, 16'h4896, 16'h4897 	:	val_out <= 16'hfd2f;
         16'h4898, 16'h4899, 16'h489a, 16'h489b, 16'h489c, 16'h489d, 16'h489e, 16'h489f 	:	val_out <= 16'hfd29;
         16'h48a0, 16'h48a1, 16'h48a2, 16'h48a3, 16'h48a4, 16'h48a5, 16'h48a6, 16'h48a7 	:	val_out <= 16'hfd24;
         16'h48a8, 16'h48a9, 16'h48aa, 16'h48ab, 16'h48ac, 16'h48ad, 16'h48ae, 16'h48af 	:	val_out <= 16'hfd1f;
         16'h48b0, 16'h48b1, 16'h48b2, 16'h48b3, 16'h48b4, 16'h48b5, 16'h48b6, 16'h48b7 	:	val_out <= 16'hfd19;
         16'h48b8, 16'h48b9, 16'h48ba, 16'h48bb, 16'h48bc, 16'h48bd, 16'h48be, 16'h48bf 	:	val_out <= 16'hfd14;
         16'h48c0, 16'h48c1, 16'h48c2, 16'h48c3, 16'h48c4, 16'h48c5, 16'h48c6, 16'h48c7 	:	val_out <= 16'hfd0f;
         16'h48c8, 16'h48c9, 16'h48ca, 16'h48cb, 16'h48cc, 16'h48cd, 16'h48ce, 16'h48cf 	:	val_out <= 16'hfd09;
         16'h48d0, 16'h48d1, 16'h48d2, 16'h48d3, 16'h48d4, 16'h48d5, 16'h48d6, 16'h48d7 	:	val_out <= 16'hfd04;
         16'h48d8, 16'h48d9, 16'h48da, 16'h48db, 16'h48dc, 16'h48dd, 16'h48de, 16'h48df 	:	val_out <= 16'hfcff;
         16'h48e0, 16'h48e1, 16'h48e2, 16'h48e3, 16'h48e4, 16'h48e5, 16'h48e6, 16'h48e7 	:	val_out <= 16'hfcf9;
         16'h48e8, 16'h48e9, 16'h48ea, 16'h48eb, 16'h48ec, 16'h48ed, 16'h48ee, 16'h48ef 	:	val_out <= 16'hfcf4;
         16'h48f0, 16'h48f1, 16'h48f2, 16'h48f3, 16'h48f4, 16'h48f5, 16'h48f6, 16'h48f7 	:	val_out <= 16'hfcee;
         16'h48f8, 16'h48f9, 16'h48fa, 16'h48fb, 16'h48fc, 16'h48fd, 16'h48fe, 16'h48ff 	:	val_out <= 16'hfce9;
         16'h4900, 16'h4901, 16'h4902, 16'h4903, 16'h4904, 16'h4905, 16'h4906, 16'h4907 	:	val_out <= 16'hfce3;
         16'h4908, 16'h4909, 16'h490a, 16'h490b, 16'h490c, 16'h490d, 16'h490e, 16'h490f 	:	val_out <= 16'hfcde;
         16'h4910, 16'h4911, 16'h4912, 16'h4913, 16'h4914, 16'h4915, 16'h4916, 16'h4917 	:	val_out <= 16'hfcd8;
         16'h4918, 16'h4919, 16'h491a, 16'h491b, 16'h491c, 16'h491d, 16'h491e, 16'h491f 	:	val_out <= 16'hfcd3;
         16'h4920, 16'h4921, 16'h4922, 16'h4923, 16'h4924, 16'h4925, 16'h4926, 16'h4927 	:	val_out <= 16'hfccd;
         16'h4928, 16'h4929, 16'h492a, 16'h492b, 16'h492c, 16'h492d, 16'h492e, 16'h492f 	:	val_out <= 16'hfcc8;
         16'h4930, 16'h4931, 16'h4932, 16'h4933, 16'h4934, 16'h4935, 16'h4936, 16'h4937 	:	val_out <= 16'hfcc2;
         16'h4938, 16'h4939, 16'h493a, 16'h493b, 16'h493c, 16'h493d, 16'h493e, 16'h493f 	:	val_out <= 16'hfcbc;
         16'h4940, 16'h4941, 16'h4942, 16'h4943, 16'h4944, 16'h4945, 16'h4946, 16'h4947 	:	val_out <= 16'hfcb7;
         16'h4948, 16'h4949, 16'h494a, 16'h494b, 16'h494c, 16'h494d, 16'h494e, 16'h494f 	:	val_out <= 16'hfcb1;
         16'h4950, 16'h4951, 16'h4952, 16'h4953, 16'h4954, 16'h4955, 16'h4956, 16'h4957 	:	val_out <= 16'hfcab;
         16'h4958, 16'h4959, 16'h495a, 16'h495b, 16'h495c, 16'h495d, 16'h495e, 16'h495f 	:	val_out <= 16'hfca6;
         16'h4960, 16'h4961, 16'h4962, 16'h4963, 16'h4964, 16'h4965, 16'h4966, 16'h4967 	:	val_out <= 16'hfca0;
         16'h4968, 16'h4969, 16'h496a, 16'h496b, 16'h496c, 16'h496d, 16'h496e, 16'h496f 	:	val_out <= 16'hfc9a;
         16'h4970, 16'h4971, 16'h4972, 16'h4973, 16'h4974, 16'h4975, 16'h4976, 16'h4977 	:	val_out <= 16'hfc94;
         16'h4978, 16'h4979, 16'h497a, 16'h497b, 16'h497c, 16'h497d, 16'h497e, 16'h497f 	:	val_out <= 16'hfc8f;
         16'h4980, 16'h4981, 16'h4982, 16'h4983, 16'h4984, 16'h4985, 16'h4986, 16'h4987 	:	val_out <= 16'hfc89;
         16'h4988, 16'h4989, 16'h498a, 16'h498b, 16'h498c, 16'h498d, 16'h498e, 16'h498f 	:	val_out <= 16'hfc83;
         16'h4990, 16'h4991, 16'h4992, 16'h4993, 16'h4994, 16'h4995, 16'h4996, 16'h4997 	:	val_out <= 16'hfc7d;
         16'h4998, 16'h4999, 16'h499a, 16'h499b, 16'h499c, 16'h499d, 16'h499e, 16'h499f 	:	val_out <= 16'hfc77;
         16'h49a0, 16'h49a1, 16'h49a2, 16'h49a3, 16'h49a4, 16'h49a5, 16'h49a6, 16'h49a7 	:	val_out <= 16'hfc71;
         16'h49a8, 16'h49a9, 16'h49aa, 16'h49ab, 16'h49ac, 16'h49ad, 16'h49ae, 16'h49af 	:	val_out <= 16'hfc6c;
         16'h49b0, 16'h49b1, 16'h49b2, 16'h49b3, 16'h49b4, 16'h49b5, 16'h49b6, 16'h49b7 	:	val_out <= 16'hfc66;
         16'h49b8, 16'h49b9, 16'h49ba, 16'h49bb, 16'h49bc, 16'h49bd, 16'h49be, 16'h49bf 	:	val_out <= 16'hfc60;
         16'h49c0, 16'h49c1, 16'h49c2, 16'h49c3, 16'h49c4, 16'h49c5, 16'h49c6, 16'h49c7 	:	val_out <= 16'hfc5a;
         16'h49c8, 16'h49c9, 16'h49ca, 16'h49cb, 16'h49cc, 16'h49cd, 16'h49ce, 16'h49cf 	:	val_out <= 16'hfc54;
         16'h49d0, 16'h49d1, 16'h49d2, 16'h49d3, 16'h49d4, 16'h49d5, 16'h49d6, 16'h49d7 	:	val_out <= 16'hfc4e;
         16'h49d8, 16'h49d9, 16'h49da, 16'h49db, 16'h49dc, 16'h49dd, 16'h49de, 16'h49df 	:	val_out <= 16'hfc48;
         16'h49e0, 16'h49e1, 16'h49e2, 16'h49e3, 16'h49e4, 16'h49e5, 16'h49e6, 16'h49e7 	:	val_out <= 16'hfc42;
         16'h49e8, 16'h49e9, 16'h49ea, 16'h49eb, 16'h49ec, 16'h49ed, 16'h49ee, 16'h49ef 	:	val_out <= 16'hfc3c;
         16'h49f0, 16'h49f1, 16'h49f2, 16'h49f3, 16'h49f4, 16'h49f5, 16'h49f6, 16'h49f7 	:	val_out <= 16'hfc36;
         16'h49f8, 16'h49f9, 16'h49fa, 16'h49fb, 16'h49fc, 16'h49fd, 16'h49fe, 16'h49ff 	:	val_out <= 16'hfc30;
         16'h4a00, 16'h4a01, 16'h4a02, 16'h4a03, 16'h4a04, 16'h4a05, 16'h4a06, 16'h4a07 	:	val_out <= 16'hfc29;
         16'h4a08, 16'h4a09, 16'h4a0a, 16'h4a0b, 16'h4a0c, 16'h4a0d, 16'h4a0e, 16'h4a0f 	:	val_out <= 16'hfc23;
         16'h4a10, 16'h4a11, 16'h4a12, 16'h4a13, 16'h4a14, 16'h4a15, 16'h4a16, 16'h4a17 	:	val_out <= 16'hfc1d;
         16'h4a18, 16'h4a19, 16'h4a1a, 16'h4a1b, 16'h4a1c, 16'h4a1d, 16'h4a1e, 16'h4a1f 	:	val_out <= 16'hfc17;
         16'h4a20, 16'h4a21, 16'h4a22, 16'h4a23, 16'h4a24, 16'h4a25, 16'h4a26, 16'h4a27 	:	val_out <= 16'hfc11;
         16'h4a28, 16'h4a29, 16'h4a2a, 16'h4a2b, 16'h4a2c, 16'h4a2d, 16'h4a2e, 16'h4a2f 	:	val_out <= 16'hfc0b;
         16'h4a30, 16'h4a31, 16'h4a32, 16'h4a33, 16'h4a34, 16'h4a35, 16'h4a36, 16'h4a37 	:	val_out <= 16'hfc05;
         16'h4a38, 16'h4a39, 16'h4a3a, 16'h4a3b, 16'h4a3c, 16'h4a3d, 16'h4a3e, 16'h4a3f 	:	val_out <= 16'hfbfe;
         16'h4a40, 16'h4a41, 16'h4a42, 16'h4a43, 16'h4a44, 16'h4a45, 16'h4a46, 16'h4a47 	:	val_out <= 16'hfbf8;
         16'h4a48, 16'h4a49, 16'h4a4a, 16'h4a4b, 16'h4a4c, 16'h4a4d, 16'h4a4e, 16'h4a4f 	:	val_out <= 16'hfbf2;
         16'h4a50, 16'h4a51, 16'h4a52, 16'h4a53, 16'h4a54, 16'h4a55, 16'h4a56, 16'h4a57 	:	val_out <= 16'hfbeb;
         16'h4a58, 16'h4a59, 16'h4a5a, 16'h4a5b, 16'h4a5c, 16'h4a5d, 16'h4a5e, 16'h4a5f 	:	val_out <= 16'hfbe5;
         16'h4a60, 16'h4a61, 16'h4a62, 16'h4a63, 16'h4a64, 16'h4a65, 16'h4a66, 16'h4a67 	:	val_out <= 16'hfbdf;
         16'h4a68, 16'h4a69, 16'h4a6a, 16'h4a6b, 16'h4a6c, 16'h4a6d, 16'h4a6e, 16'h4a6f 	:	val_out <= 16'hfbd9;
         16'h4a70, 16'h4a71, 16'h4a72, 16'h4a73, 16'h4a74, 16'h4a75, 16'h4a76, 16'h4a77 	:	val_out <= 16'hfbd2;
         16'h4a78, 16'h4a79, 16'h4a7a, 16'h4a7b, 16'h4a7c, 16'h4a7d, 16'h4a7e, 16'h4a7f 	:	val_out <= 16'hfbcc;
         16'h4a80, 16'h4a81, 16'h4a82, 16'h4a83, 16'h4a84, 16'h4a85, 16'h4a86, 16'h4a87 	:	val_out <= 16'hfbc5;
         16'h4a88, 16'h4a89, 16'h4a8a, 16'h4a8b, 16'h4a8c, 16'h4a8d, 16'h4a8e, 16'h4a8f 	:	val_out <= 16'hfbbf;
         16'h4a90, 16'h4a91, 16'h4a92, 16'h4a93, 16'h4a94, 16'h4a95, 16'h4a96, 16'h4a97 	:	val_out <= 16'hfbb9;
         16'h4a98, 16'h4a99, 16'h4a9a, 16'h4a9b, 16'h4a9c, 16'h4a9d, 16'h4a9e, 16'h4a9f 	:	val_out <= 16'hfbb2;
         16'h4aa0, 16'h4aa1, 16'h4aa2, 16'h4aa3, 16'h4aa4, 16'h4aa5, 16'h4aa6, 16'h4aa7 	:	val_out <= 16'hfbac;
         16'h4aa8, 16'h4aa9, 16'h4aaa, 16'h4aab, 16'h4aac, 16'h4aad, 16'h4aae, 16'h4aaf 	:	val_out <= 16'hfba5;
         16'h4ab0, 16'h4ab1, 16'h4ab2, 16'h4ab3, 16'h4ab4, 16'h4ab5, 16'h4ab6, 16'h4ab7 	:	val_out <= 16'hfb9f;
         16'h4ab8, 16'h4ab9, 16'h4aba, 16'h4abb, 16'h4abc, 16'h4abd, 16'h4abe, 16'h4abf 	:	val_out <= 16'hfb98;
         16'h4ac0, 16'h4ac1, 16'h4ac2, 16'h4ac3, 16'h4ac4, 16'h4ac5, 16'h4ac6, 16'h4ac7 	:	val_out <= 16'hfb92;
         16'h4ac8, 16'h4ac9, 16'h4aca, 16'h4acb, 16'h4acc, 16'h4acd, 16'h4ace, 16'h4acf 	:	val_out <= 16'hfb8b;
         16'h4ad0, 16'h4ad1, 16'h4ad2, 16'h4ad3, 16'h4ad4, 16'h4ad5, 16'h4ad6, 16'h4ad7 	:	val_out <= 16'hfb84;
         16'h4ad8, 16'h4ad9, 16'h4ada, 16'h4adb, 16'h4adc, 16'h4add, 16'h4ade, 16'h4adf 	:	val_out <= 16'hfb7e;
         16'h4ae0, 16'h4ae1, 16'h4ae2, 16'h4ae3, 16'h4ae4, 16'h4ae5, 16'h4ae6, 16'h4ae7 	:	val_out <= 16'hfb77;
         16'h4ae8, 16'h4ae9, 16'h4aea, 16'h4aeb, 16'h4aec, 16'h4aed, 16'h4aee, 16'h4aef 	:	val_out <= 16'hfb71;
         16'h4af0, 16'h4af1, 16'h4af2, 16'h4af3, 16'h4af4, 16'h4af5, 16'h4af6, 16'h4af7 	:	val_out <= 16'hfb6a;
         16'h4af8, 16'h4af9, 16'h4afa, 16'h4afb, 16'h4afc, 16'h4afd, 16'h4afe, 16'h4aff 	:	val_out <= 16'hfb63;
         16'h4b00, 16'h4b01, 16'h4b02, 16'h4b03, 16'h4b04, 16'h4b05, 16'h4b06, 16'h4b07 	:	val_out <= 16'hfb5d;
         16'h4b08, 16'h4b09, 16'h4b0a, 16'h4b0b, 16'h4b0c, 16'h4b0d, 16'h4b0e, 16'h4b0f 	:	val_out <= 16'hfb56;
         16'h4b10, 16'h4b11, 16'h4b12, 16'h4b13, 16'h4b14, 16'h4b15, 16'h4b16, 16'h4b17 	:	val_out <= 16'hfb4f;
         16'h4b18, 16'h4b19, 16'h4b1a, 16'h4b1b, 16'h4b1c, 16'h4b1d, 16'h4b1e, 16'h4b1f 	:	val_out <= 16'hfb48;
         16'h4b20, 16'h4b21, 16'h4b22, 16'h4b23, 16'h4b24, 16'h4b25, 16'h4b26, 16'h4b27 	:	val_out <= 16'hfb42;
         16'h4b28, 16'h4b29, 16'h4b2a, 16'h4b2b, 16'h4b2c, 16'h4b2d, 16'h4b2e, 16'h4b2f 	:	val_out <= 16'hfb3b;
         16'h4b30, 16'h4b31, 16'h4b32, 16'h4b33, 16'h4b34, 16'h4b35, 16'h4b36, 16'h4b37 	:	val_out <= 16'hfb34;
         16'h4b38, 16'h4b39, 16'h4b3a, 16'h4b3b, 16'h4b3c, 16'h4b3d, 16'h4b3e, 16'h4b3f 	:	val_out <= 16'hfb2d;
         16'h4b40, 16'h4b41, 16'h4b42, 16'h4b43, 16'h4b44, 16'h4b45, 16'h4b46, 16'h4b47 	:	val_out <= 16'hfb26;
         16'h4b48, 16'h4b49, 16'h4b4a, 16'h4b4b, 16'h4b4c, 16'h4b4d, 16'h4b4e, 16'h4b4f 	:	val_out <= 16'hfb1f;
         16'h4b50, 16'h4b51, 16'h4b52, 16'h4b53, 16'h4b54, 16'h4b55, 16'h4b56, 16'h4b57 	:	val_out <= 16'hfb19;
         16'h4b58, 16'h4b59, 16'h4b5a, 16'h4b5b, 16'h4b5c, 16'h4b5d, 16'h4b5e, 16'h4b5f 	:	val_out <= 16'hfb12;
         16'h4b60, 16'h4b61, 16'h4b62, 16'h4b63, 16'h4b64, 16'h4b65, 16'h4b66, 16'h4b67 	:	val_out <= 16'hfb0b;
         16'h4b68, 16'h4b69, 16'h4b6a, 16'h4b6b, 16'h4b6c, 16'h4b6d, 16'h4b6e, 16'h4b6f 	:	val_out <= 16'hfb04;
         16'h4b70, 16'h4b71, 16'h4b72, 16'h4b73, 16'h4b74, 16'h4b75, 16'h4b76, 16'h4b77 	:	val_out <= 16'hfafd;
         16'h4b78, 16'h4b79, 16'h4b7a, 16'h4b7b, 16'h4b7c, 16'h4b7d, 16'h4b7e, 16'h4b7f 	:	val_out <= 16'hfaf6;
         16'h4b80, 16'h4b81, 16'h4b82, 16'h4b83, 16'h4b84, 16'h4b85, 16'h4b86, 16'h4b87 	:	val_out <= 16'hfaef;
         16'h4b88, 16'h4b89, 16'h4b8a, 16'h4b8b, 16'h4b8c, 16'h4b8d, 16'h4b8e, 16'h4b8f 	:	val_out <= 16'hfae8;
         16'h4b90, 16'h4b91, 16'h4b92, 16'h4b93, 16'h4b94, 16'h4b95, 16'h4b96, 16'h4b97 	:	val_out <= 16'hfae1;
         16'h4b98, 16'h4b99, 16'h4b9a, 16'h4b9b, 16'h4b9c, 16'h4b9d, 16'h4b9e, 16'h4b9f 	:	val_out <= 16'hfada;
         16'h4ba0, 16'h4ba1, 16'h4ba2, 16'h4ba3, 16'h4ba4, 16'h4ba5, 16'h4ba6, 16'h4ba7 	:	val_out <= 16'hfad3;
         16'h4ba8, 16'h4ba9, 16'h4baa, 16'h4bab, 16'h4bac, 16'h4bad, 16'h4bae, 16'h4baf 	:	val_out <= 16'hfacc;
         16'h4bb0, 16'h4bb1, 16'h4bb2, 16'h4bb3, 16'h4bb4, 16'h4bb5, 16'h4bb6, 16'h4bb7 	:	val_out <= 16'hfac5;
         16'h4bb8, 16'h4bb9, 16'h4bba, 16'h4bbb, 16'h4bbc, 16'h4bbd, 16'h4bbe, 16'h4bbf 	:	val_out <= 16'hfabd;
         16'h4bc0, 16'h4bc1, 16'h4bc2, 16'h4bc3, 16'h4bc4, 16'h4bc5, 16'h4bc6, 16'h4bc7 	:	val_out <= 16'hfab6;
         16'h4bc8, 16'h4bc9, 16'h4bca, 16'h4bcb, 16'h4bcc, 16'h4bcd, 16'h4bce, 16'h4bcf 	:	val_out <= 16'hfaaf;
         16'h4bd0, 16'h4bd1, 16'h4bd2, 16'h4bd3, 16'h4bd4, 16'h4bd5, 16'h4bd6, 16'h4bd7 	:	val_out <= 16'hfaa8;
         16'h4bd8, 16'h4bd9, 16'h4bda, 16'h4bdb, 16'h4bdc, 16'h4bdd, 16'h4bde, 16'h4bdf 	:	val_out <= 16'hfaa1;
         16'h4be0, 16'h4be1, 16'h4be2, 16'h4be3, 16'h4be4, 16'h4be5, 16'h4be6, 16'h4be7 	:	val_out <= 16'hfa9a;
         16'h4be8, 16'h4be9, 16'h4bea, 16'h4beb, 16'h4bec, 16'h4bed, 16'h4bee, 16'h4bef 	:	val_out <= 16'hfa92;
         16'h4bf0, 16'h4bf1, 16'h4bf2, 16'h4bf3, 16'h4bf4, 16'h4bf5, 16'h4bf6, 16'h4bf7 	:	val_out <= 16'hfa8b;
         16'h4bf8, 16'h4bf9, 16'h4bfa, 16'h4bfb, 16'h4bfc, 16'h4bfd, 16'h4bfe, 16'h4bff 	:	val_out <= 16'hfa84;
         16'h4c00, 16'h4c01, 16'h4c02, 16'h4c03, 16'h4c04, 16'h4c05, 16'h4c06, 16'h4c07 	:	val_out <= 16'hfa7d;
         16'h4c08, 16'h4c09, 16'h4c0a, 16'h4c0b, 16'h4c0c, 16'h4c0d, 16'h4c0e, 16'h4c0f 	:	val_out <= 16'hfa75;
         16'h4c10, 16'h4c11, 16'h4c12, 16'h4c13, 16'h4c14, 16'h4c15, 16'h4c16, 16'h4c17 	:	val_out <= 16'hfa6e;
         16'h4c18, 16'h4c19, 16'h4c1a, 16'h4c1b, 16'h4c1c, 16'h4c1d, 16'h4c1e, 16'h4c1f 	:	val_out <= 16'hfa67;
         16'h4c20, 16'h4c21, 16'h4c22, 16'h4c23, 16'h4c24, 16'h4c25, 16'h4c26, 16'h4c27 	:	val_out <= 16'hfa5f;
         16'h4c28, 16'h4c29, 16'h4c2a, 16'h4c2b, 16'h4c2c, 16'h4c2d, 16'h4c2e, 16'h4c2f 	:	val_out <= 16'hfa58;
         16'h4c30, 16'h4c31, 16'h4c32, 16'h4c33, 16'h4c34, 16'h4c35, 16'h4c36, 16'h4c37 	:	val_out <= 16'hfa50;
         16'h4c38, 16'h4c39, 16'h4c3a, 16'h4c3b, 16'h4c3c, 16'h4c3d, 16'h4c3e, 16'h4c3f 	:	val_out <= 16'hfa49;
         16'h4c40, 16'h4c41, 16'h4c42, 16'h4c43, 16'h4c44, 16'h4c45, 16'h4c46, 16'h4c47 	:	val_out <= 16'hfa42;
         16'h4c48, 16'h4c49, 16'h4c4a, 16'h4c4b, 16'h4c4c, 16'h4c4d, 16'h4c4e, 16'h4c4f 	:	val_out <= 16'hfa3a;
         16'h4c50, 16'h4c51, 16'h4c52, 16'h4c53, 16'h4c54, 16'h4c55, 16'h4c56, 16'h4c57 	:	val_out <= 16'hfa33;
         16'h4c58, 16'h4c59, 16'h4c5a, 16'h4c5b, 16'h4c5c, 16'h4c5d, 16'h4c5e, 16'h4c5f 	:	val_out <= 16'hfa2b;
         16'h4c60, 16'h4c61, 16'h4c62, 16'h4c63, 16'h4c64, 16'h4c65, 16'h4c66, 16'h4c67 	:	val_out <= 16'hfa24;
         16'h4c68, 16'h4c69, 16'h4c6a, 16'h4c6b, 16'h4c6c, 16'h4c6d, 16'h4c6e, 16'h4c6f 	:	val_out <= 16'hfa1c;
         16'h4c70, 16'h4c71, 16'h4c72, 16'h4c73, 16'h4c74, 16'h4c75, 16'h4c76, 16'h4c77 	:	val_out <= 16'hfa15;
         16'h4c78, 16'h4c79, 16'h4c7a, 16'h4c7b, 16'h4c7c, 16'h4c7d, 16'h4c7e, 16'h4c7f 	:	val_out <= 16'hfa0d;
         16'h4c80, 16'h4c81, 16'h4c82, 16'h4c83, 16'h4c84, 16'h4c85, 16'h4c86, 16'h4c87 	:	val_out <= 16'hfa05;
         16'h4c88, 16'h4c89, 16'h4c8a, 16'h4c8b, 16'h4c8c, 16'h4c8d, 16'h4c8e, 16'h4c8f 	:	val_out <= 16'hf9fe;
         16'h4c90, 16'h4c91, 16'h4c92, 16'h4c93, 16'h4c94, 16'h4c95, 16'h4c96, 16'h4c97 	:	val_out <= 16'hf9f6;
         16'h4c98, 16'h4c99, 16'h4c9a, 16'h4c9b, 16'h4c9c, 16'h4c9d, 16'h4c9e, 16'h4c9f 	:	val_out <= 16'hf9ef;
         16'h4ca0, 16'h4ca1, 16'h4ca2, 16'h4ca3, 16'h4ca4, 16'h4ca5, 16'h4ca6, 16'h4ca7 	:	val_out <= 16'hf9e7;
         16'h4ca8, 16'h4ca9, 16'h4caa, 16'h4cab, 16'h4cac, 16'h4cad, 16'h4cae, 16'h4caf 	:	val_out <= 16'hf9df;
         16'h4cb0, 16'h4cb1, 16'h4cb2, 16'h4cb3, 16'h4cb4, 16'h4cb5, 16'h4cb6, 16'h4cb7 	:	val_out <= 16'hf9d8;
         16'h4cb8, 16'h4cb9, 16'h4cba, 16'h4cbb, 16'h4cbc, 16'h4cbd, 16'h4cbe, 16'h4cbf 	:	val_out <= 16'hf9d0;
         16'h4cc0, 16'h4cc1, 16'h4cc2, 16'h4cc3, 16'h4cc4, 16'h4cc5, 16'h4cc6, 16'h4cc7 	:	val_out <= 16'hf9c8;
         16'h4cc8, 16'h4cc9, 16'h4cca, 16'h4ccb, 16'h4ccc, 16'h4ccd, 16'h4cce, 16'h4ccf 	:	val_out <= 16'hf9c0;
         16'h4cd0, 16'h4cd1, 16'h4cd2, 16'h4cd3, 16'h4cd4, 16'h4cd5, 16'h4cd6, 16'h4cd7 	:	val_out <= 16'hf9b9;
         16'h4cd8, 16'h4cd9, 16'h4cda, 16'h4cdb, 16'h4cdc, 16'h4cdd, 16'h4cde, 16'h4cdf 	:	val_out <= 16'hf9b1;
         16'h4ce0, 16'h4ce1, 16'h4ce2, 16'h4ce3, 16'h4ce4, 16'h4ce5, 16'h4ce6, 16'h4ce7 	:	val_out <= 16'hf9a9;
         16'h4ce8, 16'h4ce9, 16'h4cea, 16'h4ceb, 16'h4cec, 16'h4ced, 16'h4cee, 16'h4cef 	:	val_out <= 16'hf9a1;
         16'h4cf0, 16'h4cf1, 16'h4cf2, 16'h4cf3, 16'h4cf4, 16'h4cf5, 16'h4cf6, 16'h4cf7 	:	val_out <= 16'hf999;
         16'h4cf8, 16'h4cf9, 16'h4cfa, 16'h4cfb, 16'h4cfc, 16'h4cfd, 16'h4cfe, 16'h4cff 	:	val_out <= 16'hf992;
         16'h4d00, 16'h4d01, 16'h4d02, 16'h4d03, 16'h4d04, 16'h4d05, 16'h4d06, 16'h4d07 	:	val_out <= 16'hf98a;
         16'h4d08, 16'h4d09, 16'h4d0a, 16'h4d0b, 16'h4d0c, 16'h4d0d, 16'h4d0e, 16'h4d0f 	:	val_out <= 16'hf982;
         16'h4d10, 16'h4d11, 16'h4d12, 16'h4d13, 16'h4d14, 16'h4d15, 16'h4d16, 16'h4d17 	:	val_out <= 16'hf97a;
         16'h4d18, 16'h4d19, 16'h4d1a, 16'h4d1b, 16'h4d1c, 16'h4d1d, 16'h4d1e, 16'h4d1f 	:	val_out <= 16'hf972;
         16'h4d20, 16'h4d21, 16'h4d22, 16'h4d23, 16'h4d24, 16'h4d25, 16'h4d26, 16'h4d27 	:	val_out <= 16'hf96a;
         16'h4d28, 16'h4d29, 16'h4d2a, 16'h4d2b, 16'h4d2c, 16'h4d2d, 16'h4d2e, 16'h4d2f 	:	val_out <= 16'hf962;
         16'h4d30, 16'h4d31, 16'h4d32, 16'h4d33, 16'h4d34, 16'h4d35, 16'h4d36, 16'h4d37 	:	val_out <= 16'hf95a;
         16'h4d38, 16'h4d39, 16'h4d3a, 16'h4d3b, 16'h4d3c, 16'h4d3d, 16'h4d3e, 16'h4d3f 	:	val_out <= 16'hf952;
         16'h4d40, 16'h4d41, 16'h4d42, 16'h4d43, 16'h4d44, 16'h4d45, 16'h4d46, 16'h4d47 	:	val_out <= 16'hf94a;
         16'h4d48, 16'h4d49, 16'h4d4a, 16'h4d4b, 16'h4d4c, 16'h4d4d, 16'h4d4e, 16'h4d4f 	:	val_out <= 16'hf942;
         16'h4d50, 16'h4d51, 16'h4d52, 16'h4d53, 16'h4d54, 16'h4d55, 16'h4d56, 16'h4d57 	:	val_out <= 16'hf93a;
         16'h4d58, 16'h4d59, 16'h4d5a, 16'h4d5b, 16'h4d5c, 16'h4d5d, 16'h4d5e, 16'h4d5f 	:	val_out <= 16'hf932;
         16'h4d60, 16'h4d61, 16'h4d62, 16'h4d63, 16'h4d64, 16'h4d65, 16'h4d66, 16'h4d67 	:	val_out <= 16'hf92a;
         16'h4d68, 16'h4d69, 16'h4d6a, 16'h4d6b, 16'h4d6c, 16'h4d6d, 16'h4d6e, 16'h4d6f 	:	val_out <= 16'hf922;
         16'h4d70, 16'h4d71, 16'h4d72, 16'h4d73, 16'h4d74, 16'h4d75, 16'h4d76, 16'h4d77 	:	val_out <= 16'hf919;
         16'h4d78, 16'h4d79, 16'h4d7a, 16'h4d7b, 16'h4d7c, 16'h4d7d, 16'h4d7e, 16'h4d7f 	:	val_out <= 16'hf911;
         16'h4d80, 16'h4d81, 16'h4d82, 16'h4d83, 16'h4d84, 16'h4d85, 16'h4d86, 16'h4d87 	:	val_out <= 16'hf909;
         16'h4d88, 16'h4d89, 16'h4d8a, 16'h4d8b, 16'h4d8c, 16'h4d8d, 16'h4d8e, 16'h4d8f 	:	val_out <= 16'hf901;
         16'h4d90, 16'h4d91, 16'h4d92, 16'h4d93, 16'h4d94, 16'h4d95, 16'h4d96, 16'h4d97 	:	val_out <= 16'hf8f9;
         16'h4d98, 16'h4d99, 16'h4d9a, 16'h4d9b, 16'h4d9c, 16'h4d9d, 16'h4d9e, 16'h4d9f 	:	val_out <= 16'hf8f1;
         16'h4da0, 16'h4da1, 16'h4da2, 16'h4da3, 16'h4da4, 16'h4da5, 16'h4da6, 16'h4da7 	:	val_out <= 16'hf8e8;
         16'h4da8, 16'h4da9, 16'h4daa, 16'h4dab, 16'h4dac, 16'h4dad, 16'h4dae, 16'h4daf 	:	val_out <= 16'hf8e0;
         16'h4db0, 16'h4db1, 16'h4db2, 16'h4db3, 16'h4db4, 16'h4db5, 16'h4db6, 16'h4db7 	:	val_out <= 16'hf8d8;
         16'h4db8, 16'h4db9, 16'h4dba, 16'h4dbb, 16'h4dbc, 16'h4dbd, 16'h4dbe, 16'h4dbf 	:	val_out <= 16'hf8cf;
         16'h4dc0, 16'h4dc1, 16'h4dc2, 16'h4dc3, 16'h4dc4, 16'h4dc5, 16'h4dc6, 16'h4dc7 	:	val_out <= 16'hf8c7;
         16'h4dc8, 16'h4dc9, 16'h4dca, 16'h4dcb, 16'h4dcc, 16'h4dcd, 16'h4dce, 16'h4dcf 	:	val_out <= 16'hf8bf;
         16'h4dd0, 16'h4dd1, 16'h4dd2, 16'h4dd3, 16'h4dd4, 16'h4dd5, 16'h4dd6, 16'h4dd7 	:	val_out <= 16'hf8b6;
         16'h4dd8, 16'h4dd9, 16'h4dda, 16'h4ddb, 16'h4ddc, 16'h4ddd, 16'h4dde, 16'h4ddf 	:	val_out <= 16'hf8ae;
         16'h4de0, 16'h4de1, 16'h4de2, 16'h4de3, 16'h4de4, 16'h4de5, 16'h4de6, 16'h4de7 	:	val_out <= 16'hf8a6;
         16'h4de8, 16'h4de9, 16'h4dea, 16'h4deb, 16'h4dec, 16'h4ded, 16'h4dee, 16'h4def 	:	val_out <= 16'hf89d;
         16'h4df0, 16'h4df1, 16'h4df2, 16'h4df3, 16'h4df4, 16'h4df5, 16'h4df6, 16'h4df7 	:	val_out <= 16'hf895;
         16'h4df8, 16'h4df9, 16'h4dfa, 16'h4dfb, 16'h4dfc, 16'h4dfd, 16'h4dfe, 16'h4dff 	:	val_out <= 16'hf88c;
         16'h4e00, 16'h4e01, 16'h4e02, 16'h4e03, 16'h4e04, 16'h4e05, 16'h4e06, 16'h4e07 	:	val_out <= 16'hf884;
         16'h4e08, 16'h4e09, 16'h4e0a, 16'h4e0b, 16'h4e0c, 16'h4e0d, 16'h4e0e, 16'h4e0f 	:	val_out <= 16'hf87c;
         16'h4e10, 16'h4e11, 16'h4e12, 16'h4e13, 16'h4e14, 16'h4e15, 16'h4e16, 16'h4e17 	:	val_out <= 16'hf873;
         16'h4e18, 16'h4e19, 16'h4e1a, 16'h4e1b, 16'h4e1c, 16'h4e1d, 16'h4e1e, 16'h4e1f 	:	val_out <= 16'hf86b;
         16'h4e20, 16'h4e21, 16'h4e22, 16'h4e23, 16'h4e24, 16'h4e25, 16'h4e26, 16'h4e27 	:	val_out <= 16'hf862;
         16'h4e28, 16'h4e29, 16'h4e2a, 16'h4e2b, 16'h4e2c, 16'h4e2d, 16'h4e2e, 16'h4e2f 	:	val_out <= 16'hf859;
         16'h4e30, 16'h4e31, 16'h4e32, 16'h4e33, 16'h4e34, 16'h4e35, 16'h4e36, 16'h4e37 	:	val_out <= 16'hf851;
         16'h4e38, 16'h4e39, 16'h4e3a, 16'h4e3b, 16'h4e3c, 16'h4e3d, 16'h4e3e, 16'h4e3f 	:	val_out <= 16'hf848;
         16'h4e40, 16'h4e41, 16'h4e42, 16'h4e43, 16'h4e44, 16'h4e45, 16'h4e46, 16'h4e47 	:	val_out <= 16'hf840;
         16'h4e48, 16'h4e49, 16'h4e4a, 16'h4e4b, 16'h4e4c, 16'h4e4d, 16'h4e4e, 16'h4e4f 	:	val_out <= 16'hf837;
         16'h4e50, 16'h4e51, 16'h4e52, 16'h4e53, 16'h4e54, 16'h4e55, 16'h4e56, 16'h4e57 	:	val_out <= 16'hf82e;
         16'h4e58, 16'h4e59, 16'h4e5a, 16'h4e5b, 16'h4e5c, 16'h4e5d, 16'h4e5e, 16'h4e5f 	:	val_out <= 16'hf826;
         16'h4e60, 16'h4e61, 16'h4e62, 16'h4e63, 16'h4e64, 16'h4e65, 16'h4e66, 16'h4e67 	:	val_out <= 16'hf81d;
         16'h4e68, 16'h4e69, 16'h4e6a, 16'h4e6b, 16'h4e6c, 16'h4e6d, 16'h4e6e, 16'h4e6f 	:	val_out <= 16'hf814;
         16'h4e70, 16'h4e71, 16'h4e72, 16'h4e73, 16'h4e74, 16'h4e75, 16'h4e76, 16'h4e77 	:	val_out <= 16'hf80c;
         16'h4e78, 16'h4e79, 16'h4e7a, 16'h4e7b, 16'h4e7c, 16'h4e7d, 16'h4e7e, 16'h4e7f 	:	val_out <= 16'hf803;
         16'h4e80, 16'h4e81, 16'h4e82, 16'h4e83, 16'h4e84, 16'h4e85, 16'h4e86, 16'h4e87 	:	val_out <= 16'hf7fa;
         16'h4e88, 16'h4e89, 16'h4e8a, 16'h4e8b, 16'h4e8c, 16'h4e8d, 16'h4e8e, 16'h4e8f 	:	val_out <= 16'hf7f1;
         16'h4e90, 16'h4e91, 16'h4e92, 16'h4e93, 16'h4e94, 16'h4e95, 16'h4e96, 16'h4e97 	:	val_out <= 16'hf7e9;
         16'h4e98, 16'h4e99, 16'h4e9a, 16'h4e9b, 16'h4e9c, 16'h4e9d, 16'h4e9e, 16'h4e9f 	:	val_out <= 16'hf7e0;
         16'h4ea0, 16'h4ea1, 16'h4ea2, 16'h4ea3, 16'h4ea4, 16'h4ea5, 16'h4ea6, 16'h4ea7 	:	val_out <= 16'hf7d7;
         16'h4ea8, 16'h4ea9, 16'h4eaa, 16'h4eab, 16'h4eac, 16'h4ead, 16'h4eae, 16'h4eaf 	:	val_out <= 16'hf7ce;
         16'h4eb0, 16'h4eb1, 16'h4eb2, 16'h4eb3, 16'h4eb4, 16'h4eb5, 16'h4eb6, 16'h4eb7 	:	val_out <= 16'hf7c5;
         16'h4eb8, 16'h4eb9, 16'h4eba, 16'h4ebb, 16'h4ebc, 16'h4ebd, 16'h4ebe, 16'h4ebf 	:	val_out <= 16'hf7bc;
         16'h4ec0, 16'h4ec1, 16'h4ec2, 16'h4ec3, 16'h4ec4, 16'h4ec5, 16'h4ec6, 16'h4ec7 	:	val_out <= 16'hf7b4;
         16'h4ec8, 16'h4ec9, 16'h4eca, 16'h4ecb, 16'h4ecc, 16'h4ecd, 16'h4ece, 16'h4ecf 	:	val_out <= 16'hf7ab;
         16'h4ed0, 16'h4ed1, 16'h4ed2, 16'h4ed3, 16'h4ed4, 16'h4ed5, 16'h4ed6, 16'h4ed7 	:	val_out <= 16'hf7a2;
         16'h4ed8, 16'h4ed9, 16'h4eda, 16'h4edb, 16'h4edc, 16'h4edd, 16'h4ede, 16'h4edf 	:	val_out <= 16'hf799;
         16'h4ee0, 16'h4ee1, 16'h4ee2, 16'h4ee3, 16'h4ee4, 16'h4ee5, 16'h4ee6, 16'h4ee7 	:	val_out <= 16'hf790;
         16'h4ee8, 16'h4ee9, 16'h4eea, 16'h4eeb, 16'h4eec, 16'h4eed, 16'h4eee, 16'h4eef 	:	val_out <= 16'hf787;
         16'h4ef0, 16'h4ef1, 16'h4ef2, 16'h4ef3, 16'h4ef4, 16'h4ef5, 16'h4ef6, 16'h4ef7 	:	val_out <= 16'hf77e;
         16'h4ef8, 16'h4ef9, 16'h4efa, 16'h4efb, 16'h4efc, 16'h4efd, 16'h4efe, 16'h4eff 	:	val_out <= 16'hf775;
         16'h4f00, 16'h4f01, 16'h4f02, 16'h4f03, 16'h4f04, 16'h4f05, 16'h4f06, 16'h4f07 	:	val_out <= 16'hf76c;
         16'h4f08, 16'h4f09, 16'h4f0a, 16'h4f0b, 16'h4f0c, 16'h4f0d, 16'h4f0e, 16'h4f0f 	:	val_out <= 16'hf763;
         16'h4f10, 16'h4f11, 16'h4f12, 16'h4f13, 16'h4f14, 16'h4f15, 16'h4f16, 16'h4f17 	:	val_out <= 16'hf75a;
         16'h4f18, 16'h4f19, 16'h4f1a, 16'h4f1b, 16'h4f1c, 16'h4f1d, 16'h4f1e, 16'h4f1f 	:	val_out <= 16'hf751;
         16'h4f20, 16'h4f21, 16'h4f22, 16'h4f23, 16'h4f24, 16'h4f25, 16'h4f26, 16'h4f27 	:	val_out <= 16'hf747;
         16'h4f28, 16'h4f29, 16'h4f2a, 16'h4f2b, 16'h4f2c, 16'h4f2d, 16'h4f2e, 16'h4f2f 	:	val_out <= 16'hf73e;
         16'h4f30, 16'h4f31, 16'h4f32, 16'h4f33, 16'h4f34, 16'h4f35, 16'h4f36, 16'h4f37 	:	val_out <= 16'hf735;
         16'h4f38, 16'h4f39, 16'h4f3a, 16'h4f3b, 16'h4f3c, 16'h4f3d, 16'h4f3e, 16'h4f3f 	:	val_out <= 16'hf72c;
         16'h4f40, 16'h4f41, 16'h4f42, 16'h4f43, 16'h4f44, 16'h4f45, 16'h4f46, 16'h4f47 	:	val_out <= 16'hf723;
         16'h4f48, 16'h4f49, 16'h4f4a, 16'h4f4b, 16'h4f4c, 16'h4f4d, 16'h4f4e, 16'h4f4f 	:	val_out <= 16'hf71a;
         16'h4f50, 16'h4f51, 16'h4f52, 16'h4f53, 16'h4f54, 16'h4f55, 16'h4f56, 16'h4f57 	:	val_out <= 16'hf710;
         16'h4f58, 16'h4f59, 16'h4f5a, 16'h4f5b, 16'h4f5c, 16'h4f5d, 16'h4f5e, 16'h4f5f 	:	val_out <= 16'hf707;
         16'h4f60, 16'h4f61, 16'h4f62, 16'h4f63, 16'h4f64, 16'h4f65, 16'h4f66, 16'h4f67 	:	val_out <= 16'hf6fe;
         16'h4f68, 16'h4f69, 16'h4f6a, 16'h4f6b, 16'h4f6c, 16'h4f6d, 16'h4f6e, 16'h4f6f 	:	val_out <= 16'hf6f5;
         16'h4f70, 16'h4f71, 16'h4f72, 16'h4f73, 16'h4f74, 16'h4f75, 16'h4f76, 16'h4f77 	:	val_out <= 16'hf6eb;
         16'h4f78, 16'h4f79, 16'h4f7a, 16'h4f7b, 16'h4f7c, 16'h4f7d, 16'h4f7e, 16'h4f7f 	:	val_out <= 16'hf6e2;
         16'h4f80, 16'h4f81, 16'h4f82, 16'h4f83, 16'h4f84, 16'h4f85, 16'h4f86, 16'h4f87 	:	val_out <= 16'hf6d9;
         16'h4f88, 16'h4f89, 16'h4f8a, 16'h4f8b, 16'h4f8c, 16'h4f8d, 16'h4f8e, 16'h4f8f 	:	val_out <= 16'hf6cf;
         16'h4f90, 16'h4f91, 16'h4f92, 16'h4f93, 16'h4f94, 16'h4f95, 16'h4f96, 16'h4f97 	:	val_out <= 16'hf6c6;
         16'h4f98, 16'h4f99, 16'h4f9a, 16'h4f9b, 16'h4f9c, 16'h4f9d, 16'h4f9e, 16'h4f9f 	:	val_out <= 16'hf6bd;
         16'h4fa0, 16'h4fa1, 16'h4fa2, 16'h4fa3, 16'h4fa4, 16'h4fa5, 16'h4fa6, 16'h4fa7 	:	val_out <= 16'hf6b3;
         16'h4fa8, 16'h4fa9, 16'h4faa, 16'h4fab, 16'h4fac, 16'h4fad, 16'h4fae, 16'h4faf 	:	val_out <= 16'hf6aa;
         16'h4fb0, 16'h4fb1, 16'h4fb2, 16'h4fb3, 16'h4fb4, 16'h4fb5, 16'h4fb6, 16'h4fb7 	:	val_out <= 16'hf6a0;
         16'h4fb8, 16'h4fb9, 16'h4fba, 16'h4fbb, 16'h4fbc, 16'h4fbd, 16'h4fbe, 16'h4fbf 	:	val_out <= 16'hf697;
         16'h4fc0, 16'h4fc1, 16'h4fc2, 16'h4fc3, 16'h4fc4, 16'h4fc5, 16'h4fc6, 16'h4fc7 	:	val_out <= 16'hf68e;
         16'h4fc8, 16'h4fc9, 16'h4fca, 16'h4fcb, 16'h4fcc, 16'h4fcd, 16'h4fce, 16'h4fcf 	:	val_out <= 16'hf684;
         16'h4fd0, 16'h4fd1, 16'h4fd2, 16'h4fd3, 16'h4fd4, 16'h4fd5, 16'h4fd6, 16'h4fd7 	:	val_out <= 16'hf67b;
         16'h4fd8, 16'h4fd9, 16'h4fda, 16'h4fdb, 16'h4fdc, 16'h4fdd, 16'h4fde, 16'h4fdf 	:	val_out <= 16'hf671;
         16'h4fe0, 16'h4fe1, 16'h4fe2, 16'h4fe3, 16'h4fe4, 16'h4fe5, 16'h4fe6, 16'h4fe7 	:	val_out <= 16'hf668;
         16'h4fe8, 16'h4fe9, 16'h4fea, 16'h4feb, 16'h4fec, 16'h4fed, 16'h4fee, 16'h4fef 	:	val_out <= 16'hf65e;
         16'h4ff0, 16'h4ff1, 16'h4ff2, 16'h4ff3, 16'h4ff4, 16'h4ff5, 16'h4ff6, 16'h4ff7 	:	val_out <= 16'hf654;
         16'h4ff8, 16'h4ff9, 16'h4ffa, 16'h4ffb, 16'h4ffc, 16'h4ffd, 16'h4ffe, 16'h4fff 	:	val_out <= 16'hf64b;
         16'h5000, 16'h5001, 16'h5002, 16'h5003, 16'h5004, 16'h5005, 16'h5006, 16'h5007 	:	val_out <= 16'hf641;
         16'h5008, 16'h5009, 16'h500a, 16'h500b, 16'h500c, 16'h500d, 16'h500e, 16'h500f 	:	val_out <= 16'hf638;
         16'h5010, 16'h5011, 16'h5012, 16'h5013, 16'h5014, 16'h5015, 16'h5016, 16'h5017 	:	val_out <= 16'hf62e;
         16'h5018, 16'h5019, 16'h501a, 16'h501b, 16'h501c, 16'h501d, 16'h501e, 16'h501f 	:	val_out <= 16'hf624;
         16'h5020, 16'h5021, 16'h5022, 16'h5023, 16'h5024, 16'h5025, 16'h5026, 16'h5027 	:	val_out <= 16'hf61b;
         16'h5028, 16'h5029, 16'h502a, 16'h502b, 16'h502c, 16'h502d, 16'h502e, 16'h502f 	:	val_out <= 16'hf611;
         16'h5030, 16'h5031, 16'h5032, 16'h5033, 16'h5034, 16'h5035, 16'h5036, 16'h5037 	:	val_out <= 16'hf607;
         16'h5038, 16'h5039, 16'h503a, 16'h503b, 16'h503c, 16'h503d, 16'h503e, 16'h503f 	:	val_out <= 16'hf5fd;
         16'h5040, 16'h5041, 16'h5042, 16'h5043, 16'h5044, 16'h5045, 16'h5046, 16'h5047 	:	val_out <= 16'hf5f4;
         16'h5048, 16'h5049, 16'h504a, 16'h504b, 16'h504c, 16'h504d, 16'h504e, 16'h504f 	:	val_out <= 16'hf5ea;
         16'h5050, 16'h5051, 16'h5052, 16'h5053, 16'h5054, 16'h5055, 16'h5056, 16'h5057 	:	val_out <= 16'hf5e0;
         16'h5058, 16'h5059, 16'h505a, 16'h505b, 16'h505c, 16'h505d, 16'h505e, 16'h505f 	:	val_out <= 16'hf5d6;
         16'h5060, 16'h5061, 16'h5062, 16'h5063, 16'h5064, 16'h5065, 16'h5066, 16'h5067 	:	val_out <= 16'hf5cc;
         16'h5068, 16'h5069, 16'h506a, 16'h506b, 16'h506c, 16'h506d, 16'h506e, 16'h506f 	:	val_out <= 16'hf5c3;
         16'h5070, 16'h5071, 16'h5072, 16'h5073, 16'h5074, 16'h5075, 16'h5076, 16'h5077 	:	val_out <= 16'hf5b9;
         16'h5078, 16'h5079, 16'h507a, 16'h507b, 16'h507c, 16'h507d, 16'h507e, 16'h507f 	:	val_out <= 16'hf5af;
         16'h5080, 16'h5081, 16'h5082, 16'h5083, 16'h5084, 16'h5085, 16'h5086, 16'h5087 	:	val_out <= 16'hf5a5;
         16'h5088, 16'h5089, 16'h508a, 16'h508b, 16'h508c, 16'h508d, 16'h508e, 16'h508f 	:	val_out <= 16'hf59b;
         16'h5090, 16'h5091, 16'h5092, 16'h5093, 16'h5094, 16'h5095, 16'h5096, 16'h5097 	:	val_out <= 16'hf591;
         16'h5098, 16'h5099, 16'h509a, 16'h509b, 16'h509c, 16'h509d, 16'h509e, 16'h509f 	:	val_out <= 16'hf587;
         16'h50a0, 16'h50a1, 16'h50a2, 16'h50a3, 16'h50a4, 16'h50a5, 16'h50a6, 16'h50a7 	:	val_out <= 16'hf57d;
         16'h50a8, 16'h50a9, 16'h50aa, 16'h50ab, 16'h50ac, 16'h50ad, 16'h50ae, 16'h50af 	:	val_out <= 16'hf573;
         16'h50b0, 16'h50b1, 16'h50b2, 16'h50b3, 16'h50b4, 16'h50b5, 16'h50b6, 16'h50b7 	:	val_out <= 16'hf569;
         16'h50b8, 16'h50b9, 16'h50ba, 16'h50bb, 16'h50bc, 16'h50bd, 16'h50be, 16'h50bf 	:	val_out <= 16'hf55f;
         16'h50c0, 16'h50c1, 16'h50c2, 16'h50c3, 16'h50c4, 16'h50c5, 16'h50c6, 16'h50c7 	:	val_out <= 16'hf555;
         16'h50c8, 16'h50c9, 16'h50ca, 16'h50cb, 16'h50cc, 16'h50cd, 16'h50ce, 16'h50cf 	:	val_out <= 16'hf54b;
         16'h50d0, 16'h50d1, 16'h50d2, 16'h50d3, 16'h50d4, 16'h50d5, 16'h50d6, 16'h50d7 	:	val_out <= 16'hf541;
         16'h50d8, 16'h50d9, 16'h50da, 16'h50db, 16'h50dc, 16'h50dd, 16'h50de, 16'h50df 	:	val_out <= 16'hf537;
         16'h50e0, 16'h50e1, 16'h50e2, 16'h50e3, 16'h50e4, 16'h50e5, 16'h50e6, 16'h50e7 	:	val_out <= 16'hf52d;
         16'h50e8, 16'h50e9, 16'h50ea, 16'h50eb, 16'h50ec, 16'h50ed, 16'h50ee, 16'h50ef 	:	val_out <= 16'hf523;
         16'h50f0, 16'h50f1, 16'h50f2, 16'h50f3, 16'h50f4, 16'h50f5, 16'h50f6, 16'h50f7 	:	val_out <= 16'hf519;
         16'h50f8, 16'h50f9, 16'h50fa, 16'h50fb, 16'h50fc, 16'h50fd, 16'h50fe, 16'h50ff 	:	val_out <= 16'hf50f;
         16'h5100, 16'h5101, 16'h5102, 16'h5103, 16'h5104, 16'h5105, 16'h5106, 16'h5107 	:	val_out <= 16'hf504;
         16'h5108, 16'h5109, 16'h510a, 16'h510b, 16'h510c, 16'h510d, 16'h510e, 16'h510f 	:	val_out <= 16'hf4fa;
         16'h5110, 16'h5111, 16'h5112, 16'h5113, 16'h5114, 16'h5115, 16'h5116, 16'h5117 	:	val_out <= 16'hf4f0;
         16'h5118, 16'h5119, 16'h511a, 16'h511b, 16'h511c, 16'h511d, 16'h511e, 16'h511f 	:	val_out <= 16'hf4e6;
         16'h5120, 16'h5121, 16'h5122, 16'h5123, 16'h5124, 16'h5125, 16'h5126, 16'h5127 	:	val_out <= 16'hf4db;
         16'h5128, 16'h5129, 16'h512a, 16'h512b, 16'h512c, 16'h512d, 16'h512e, 16'h512f 	:	val_out <= 16'hf4d1;
         16'h5130, 16'h5131, 16'h5132, 16'h5133, 16'h5134, 16'h5135, 16'h5136, 16'h5137 	:	val_out <= 16'hf4c7;
         16'h5138, 16'h5139, 16'h513a, 16'h513b, 16'h513c, 16'h513d, 16'h513e, 16'h513f 	:	val_out <= 16'hf4bd;
         16'h5140, 16'h5141, 16'h5142, 16'h5143, 16'h5144, 16'h5145, 16'h5146, 16'h5147 	:	val_out <= 16'hf4b2;
         16'h5148, 16'h5149, 16'h514a, 16'h514b, 16'h514c, 16'h514d, 16'h514e, 16'h514f 	:	val_out <= 16'hf4a8;
         16'h5150, 16'h5151, 16'h5152, 16'h5153, 16'h5154, 16'h5155, 16'h5156, 16'h5157 	:	val_out <= 16'hf49e;
         16'h5158, 16'h5159, 16'h515a, 16'h515b, 16'h515c, 16'h515d, 16'h515e, 16'h515f 	:	val_out <= 16'hf493;
         16'h5160, 16'h5161, 16'h5162, 16'h5163, 16'h5164, 16'h5165, 16'h5166, 16'h5167 	:	val_out <= 16'hf489;
         16'h5168, 16'h5169, 16'h516a, 16'h516b, 16'h516c, 16'h516d, 16'h516e, 16'h516f 	:	val_out <= 16'hf47e;
         16'h5170, 16'h5171, 16'h5172, 16'h5173, 16'h5174, 16'h5175, 16'h5176, 16'h5177 	:	val_out <= 16'hf474;
         16'h5178, 16'h5179, 16'h517a, 16'h517b, 16'h517c, 16'h517d, 16'h517e, 16'h517f 	:	val_out <= 16'hf46a;
         16'h5180, 16'h5181, 16'h5182, 16'h5183, 16'h5184, 16'h5185, 16'h5186, 16'h5187 	:	val_out <= 16'hf45f;
         16'h5188, 16'h5189, 16'h518a, 16'h518b, 16'h518c, 16'h518d, 16'h518e, 16'h518f 	:	val_out <= 16'hf455;
         16'h5190, 16'h5191, 16'h5192, 16'h5193, 16'h5194, 16'h5195, 16'h5196, 16'h5197 	:	val_out <= 16'hf44a;
         16'h5198, 16'h5199, 16'h519a, 16'h519b, 16'h519c, 16'h519d, 16'h519e, 16'h519f 	:	val_out <= 16'hf440;
         16'h51a0, 16'h51a1, 16'h51a2, 16'h51a3, 16'h51a4, 16'h51a5, 16'h51a6, 16'h51a7 	:	val_out <= 16'hf435;
         16'h51a8, 16'h51a9, 16'h51aa, 16'h51ab, 16'h51ac, 16'h51ad, 16'h51ae, 16'h51af 	:	val_out <= 16'hf42b;
         16'h51b0, 16'h51b1, 16'h51b2, 16'h51b3, 16'h51b4, 16'h51b5, 16'h51b6, 16'h51b7 	:	val_out <= 16'hf420;
         16'h51b8, 16'h51b9, 16'h51ba, 16'h51bb, 16'h51bc, 16'h51bd, 16'h51be, 16'h51bf 	:	val_out <= 16'hf415;
         16'h51c0, 16'h51c1, 16'h51c2, 16'h51c3, 16'h51c4, 16'h51c5, 16'h51c6, 16'h51c7 	:	val_out <= 16'hf40b;
         16'h51c8, 16'h51c9, 16'h51ca, 16'h51cb, 16'h51cc, 16'h51cd, 16'h51ce, 16'h51cf 	:	val_out <= 16'hf400;
         16'h51d0, 16'h51d1, 16'h51d2, 16'h51d3, 16'h51d4, 16'h51d5, 16'h51d6, 16'h51d7 	:	val_out <= 16'hf3f6;
         16'h51d8, 16'h51d9, 16'h51da, 16'h51db, 16'h51dc, 16'h51dd, 16'h51de, 16'h51df 	:	val_out <= 16'hf3eb;
         16'h51e0, 16'h51e1, 16'h51e2, 16'h51e3, 16'h51e4, 16'h51e5, 16'h51e6, 16'h51e7 	:	val_out <= 16'hf3e0;
         16'h51e8, 16'h51e9, 16'h51ea, 16'h51eb, 16'h51ec, 16'h51ed, 16'h51ee, 16'h51ef 	:	val_out <= 16'hf3d6;
         16'h51f0, 16'h51f1, 16'h51f2, 16'h51f3, 16'h51f4, 16'h51f5, 16'h51f6, 16'h51f7 	:	val_out <= 16'hf3cb;
         16'h51f8, 16'h51f9, 16'h51fa, 16'h51fb, 16'h51fc, 16'h51fd, 16'h51fe, 16'h51ff 	:	val_out <= 16'hf3c0;
         16'h5200, 16'h5201, 16'h5202, 16'h5203, 16'h5204, 16'h5205, 16'h5206, 16'h5207 	:	val_out <= 16'hf3b5;
         16'h5208, 16'h5209, 16'h520a, 16'h520b, 16'h520c, 16'h520d, 16'h520e, 16'h520f 	:	val_out <= 16'hf3ab;
         16'h5210, 16'h5211, 16'h5212, 16'h5213, 16'h5214, 16'h5215, 16'h5216, 16'h5217 	:	val_out <= 16'hf3a0;
         16'h5218, 16'h5219, 16'h521a, 16'h521b, 16'h521c, 16'h521d, 16'h521e, 16'h521f 	:	val_out <= 16'hf395;
         16'h5220, 16'h5221, 16'h5222, 16'h5223, 16'h5224, 16'h5225, 16'h5226, 16'h5227 	:	val_out <= 16'hf38a;
         16'h5228, 16'h5229, 16'h522a, 16'h522b, 16'h522c, 16'h522d, 16'h522e, 16'h522f 	:	val_out <= 16'hf37f;
         16'h5230, 16'h5231, 16'h5232, 16'h5233, 16'h5234, 16'h5235, 16'h5236, 16'h5237 	:	val_out <= 16'hf375;
         16'h5238, 16'h5239, 16'h523a, 16'h523b, 16'h523c, 16'h523d, 16'h523e, 16'h523f 	:	val_out <= 16'hf36a;
         16'h5240, 16'h5241, 16'h5242, 16'h5243, 16'h5244, 16'h5245, 16'h5246, 16'h5247 	:	val_out <= 16'hf35f;
         16'h5248, 16'h5249, 16'h524a, 16'h524b, 16'h524c, 16'h524d, 16'h524e, 16'h524f 	:	val_out <= 16'hf354;
         16'h5250, 16'h5251, 16'h5252, 16'h5253, 16'h5254, 16'h5255, 16'h5256, 16'h5257 	:	val_out <= 16'hf349;
         16'h5258, 16'h5259, 16'h525a, 16'h525b, 16'h525c, 16'h525d, 16'h525e, 16'h525f 	:	val_out <= 16'hf33e;
         16'h5260, 16'h5261, 16'h5262, 16'h5263, 16'h5264, 16'h5265, 16'h5266, 16'h5267 	:	val_out <= 16'hf333;
         16'h5268, 16'h5269, 16'h526a, 16'h526b, 16'h526c, 16'h526d, 16'h526e, 16'h526f 	:	val_out <= 16'hf328;
         16'h5270, 16'h5271, 16'h5272, 16'h5273, 16'h5274, 16'h5275, 16'h5276, 16'h5277 	:	val_out <= 16'hf31d;
         16'h5278, 16'h5279, 16'h527a, 16'h527b, 16'h527c, 16'h527d, 16'h527e, 16'h527f 	:	val_out <= 16'hf312;
         16'h5280, 16'h5281, 16'h5282, 16'h5283, 16'h5284, 16'h5285, 16'h5286, 16'h5287 	:	val_out <= 16'hf307;
         16'h5288, 16'h5289, 16'h528a, 16'h528b, 16'h528c, 16'h528d, 16'h528e, 16'h528f 	:	val_out <= 16'hf2fc;
         16'h5290, 16'h5291, 16'h5292, 16'h5293, 16'h5294, 16'h5295, 16'h5296, 16'h5297 	:	val_out <= 16'hf2f1;
         16'h5298, 16'h5299, 16'h529a, 16'h529b, 16'h529c, 16'h529d, 16'h529e, 16'h529f 	:	val_out <= 16'hf2e6;
         16'h52a0, 16'h52a1, 16'h52a2, 16'h52a3, 16'h52a4, 16'h52a5, 16'h52a6, 16'h52a7 	:	val_out <= 16'hf2db;
         16'h52a8, 16'h52a9, 16'h52aa, 16'h52ab, 16'h52ac, 16'h52ad, 16'h52ae, 16'h52af 	:	val_out <= 16'hf2d0;
         16'h52b0, 16'h52b1, 16'h52b2, 16'h52b3, 16'h52b4, 16'h52b5, 16'h52b6, 16'h52b7 	:	val_out <= 16'hf2c5;
         16'h52b8, 16'h52b9, 16'h52ba, 16'h52bb, 16'h52bc, 16'h52bd, 16'h52be, 16'h52bf 	:	val_out <= 16'hf2ba;
         16'h52c0, 16'h52c1, 16'h52c2, 16'h52c3, 16'h52c4, 16'h52c5, 16'h52c6, 16'h52c7 	:	val_out <= 16'hf2af;
         16'h52c8, 16'h52c9, 16'h52ca, 16'h52cb, 16'h52cc, 16'h52cd, 16'h52ce, 16'h52cf 	:	val_out <= 16'hf2a3;
         16'h52d0, 16'h52d1, 16'h52d2, 16'h52d3, 16'h52d4, 16'h52d5, 16'h52d6, 16'h52d7 	:	val_out <= 16'hf298;
         16'h52d8, 16'h52d9, 16'h52da, 16'h52db, 16'h52dc, 16'h52dd, 16'h52de, 16'h52df 	:	val_out <= 16'hf28d;
         16'h52e0, 16'h52e1, 16'h52e2, 16'h52e3, 16'h52e4, 16'h52e5, 16'h52e6, 16'h52e7 	:	val_out <= 16'hf282;
         16'h52e8, 16'h52e9, 16'h52ea, 16'h52eb, 16'h52ec, 16'h52ed, 16'h52ee, 16'h52ef 	:	val_out <= 16'hf276;
         16'h52f0, 16'h52f1, 16'h52f2, 16'h52f3, 16'h52f4, 16'h52f5, 16'h52f6, 16'h52f7 	:	val_out <= 16'hf26b;
         16'h52f8, 16'h52f9, 16'h52fa, 16'h52fb, 16'h52fc, 16'h52fd, 16'h52fe, 16'h52ff 	:	val_out <= 16'hf260;
         16'h5300, 16'h5301, 16'h5302, 16'h5303, 16'h5304, 16'h5305, 16'h5306, 16'h5307 	:	val_out <= 16'hf255;
         16'h5308, 16'h5309, 16'h530a, 16'h530b, 16'h530c, 16'h530d, 16'h530e, 16'h530f 	:	val_out <= 16'hf249;
         16'h5310, 16'h5311, 16'h5312, 16'h5313, 16'h5314, 16'h5315, 16'h5316, 16'h5317 	:	val_out <= 16'hf23e;
         16'h5318, 16'h5319, 16'h531a, 16'h531b, 16'h531c, 16'h531d, 16'h531e, 16'h531f 	:	val_out <= 16'hf233;
         16'h5320, 16'h5321, 16'h5322, 16'h5323, 16'h5324, 16'h5325, 16'h5326, 16'h5327 	:	val_out <= 16'hf227;
         16'h5328, 16'h5329, 16'h532a, 16'h532b, 16'h532c, 16'h532d, 16'h532e, 16'h532f 	:	val_out <= 16'hf21c;
         16'h5330, 16'h5331, 16'h5332, 16'h5333, 16'h5334, 16'h5335, 16'h5336, 16'h5337 	:	val_out <= 16'hf211;
         16'h5338, 16'h5339, 16'h533a, 16'h533b, 16'h533c, 16'h533d, 16'h533e, 16'h533f 	:	val_out <= 16'hf205;
         16'h5340, 16'h5341, 16'h5342, 16'h5343, 16'h5344, 16'h5345, 16'h5346, 16'h5347 	:	val_out <= 16'hf1fa;
         16'h5348, 16'h5349, 16'h534a, 16'h534b, 16'h534c, 16'h534d, 16'h534e, 16'h534f 	:	val_out <= 16'hf1ee;
         16'h5350, 16'h5351, 16'h5352, 16'h5353, 16'h5354, 16'h5355, 16'h5356, 16'h5357 	:	val_out <= 16'hf1e3;
         16'h5358, 16'h5359, 16'h535a, 16'h535b, 16'h535c, 16'h535d, 16'h535e, 16'h535f 	:	val_out <= 16'hf1d7;
         16'h5360, 16'h5361, 16'h5362, 16'h5363, 16'h5364, 16'h5365, 16'h5366, 16'h5367 	:	val_out <= 16'hf1cc;
         16'h5368, 16'h5369, 16'h536a, 16'h536b, 16'h536c, 16'h536d, 16'h536e, 16'h536f 	:	val_out <= 16'hf1c0;
         16'h5370, 16'h5371, 16'h5372, 16'h5373, 16'h5374, 16'h5375, 16'h5376, 16'h5377 	:	val_out <= 16'hf1b5;
         16'h5378, 16'h5379, 16'h537a, 16'h537b, 16'h537c, 16'h537d, 16'h537e, 16'h537f 	:	val_out <= 16'hf1a9;
         16'h5380, 16'h5381, 16'h5382, 16'h5383, 16'h5384, 16'h5385, 16'h5386, 16'h5387 	:	val_out <= 16'hf19e;
         16'h5388, 16'h5389, 16'h538a, 16'h538b, 16'h538c, 16'h538d, 16'h538e, 16'h538f 	:	val_out <= 16'hf192;
         16'h5390, 16'h5391, 16'h5392, 16'h5393, 16'h5394, 16'h5395, 16'h5396, 16'h5397 	:	val_out <= 16'hf186;
         16'h5398, 16'h5399, 16'h539a, 16'h539b, 16'h539c, 16'h539d, 16'h539e, 16'h539f 	:	val_out <= 16'hf17b;
         16'h53a0, 16'h53a1, 16'h53a2, 16'h53a3, 16'h53a4, 16'h53a5, 16'h53a6, 16'h53a7 	:	val_out <= 16'hf16f;
         16'h53a8, 16'h53a9, 16'h53aa, 16'h53ab, 16'h53ac, 16'h53ad, 16'h53ae, 16'h53af 	:	val_out <= 16'hf164;
         16'h53b0, 16'h53b1, 16'h53b2, 16'h53b3, 16'h53b4, 16'h53b5, 16'h53b6, 16'h53b7 	:	val_out <= 16'hf158;
         16'h53b8, 16'h53b9, 16'h53ba, 16'h53bb, 16'h53bc, 16'h53bd, 16'h53be, 16'h53bf 	:	val_out <= 16'hf14c;
         16'h53c0, 16'h53c1, 16'h53c2, 16'h53c3, 16'h53c4, 16'h53c5, 16'h53c6, 16'h53c7 	:	val_out <= 16'hf141;
         16'h53c8, 16'h53c9, 16'h53ca, 16'h53cb, 16'h53cc, 16'h53cd, 16'h53ce, 16'h53cf 	:	val_out <= 16'hf135;
         16'h53d0, 16'h53d1, 16'h53d2, 16'h53d3, 16'h53d4, 16'h53d5, 16'h53d6, 16'h53d7 	:	val_out <= 16'hf129;
         16'h53d8, 16'h53d9, 16'h53da, 16'h53db, 16'h53dc, 16'h53dd, 16'h53de, 16'h53df 	:	val_out <= 16'hf11d;
         16'h53e0, 16'h53e1, 16'h53e2, 16'h53e3, 16'h53e4, 16'h53e5, 16'h53e6, 16'h53e7 	:	val_out <= 16'hf112;
         16'h53e8, 16'h53e9, 16'h53ea, 16'h53eb, 16'h53ec, 16'h53ed, 16'h53ee, 16'h53ef 	:	val_out <= 16'hf106;
         16'h53f0, 16'h53f1, 16'h53f2, 16'h53f3, 16'h53f4, 16'h53f5, 16'h53f6, 16'h53f7 	:	val_out <= 16'hf0fa;
         16'h53f8, 16'h53f9, 16'h53fa, 16'h53fb, 16'h53fc, 16'h53fd, 16'h53fe, 16'h53ff 	:	val_out <= 16'hf0ee;
         16'h5400, 16'h5401, 16'h5402, 16'h5403, 16'h5404, 16'h5405, 16'h5406, 16'h5407 	:	val_out <= 16'hf0e2;
         16'h5408, 16'h5409, 16'h540a, 16'h540b, 16'h540c, 16'h540d, 16'h540e, 16'h540f 	:	val_out <= 16'hf0d6;
         16'h5410, 16'h5411, 16'h5412, 16'h5413, 16'h5414, 16'h5415, 16'h5416, 16'h5417 	:	val_out <= 16'hf0cb;
         16'h5418, 16'h5419, 16'h541a, 16'h541b, 16'h541c, 16'h541d, 16'h541e, 16'h541f 	:	val_out <= 16'hf0bf;
         16'h5420, 16'h5421, 16'h5422, 16'h5423, 16'h5424, 16'h5425, 16'h5426, 16'h5427 	:	val_out <= 16'hf0b3;
         16'h5428, 16'h5429, 16'h542a, 16'h542b, 16'h542c, 16'h542d, 16'h542e, 16'h542f 	:	val_out <= 16'hf0a7;
         16'h5430, 16'h5431, 16'h5432, 16'h5433, 16'h5434, 16'h5435, 16'h5436, 16'h5437 	:	val_out <= 16'hf09b;
         16'h5438, 16'h5439, 16'h543a, 16'h543b, 16'h543c, 16'h543d, 16'h543e, 16'h543f 	:	val_out <= 16'hf08f;
         16'h5440, 16'h5441, 16'h5442, 16'h5443, 16'h5444, 16'h5445, 16'h5446, 16'h5447 	:	val_out <= 16'hf083;
         16'h5448, 16'h5449, 16'h544a, 16'h544b, 16'h544c, 16'h544d, 16'h544e, 16'h544f 	:	val_out <= 16'hf077;
         16'h5450, 16'h5451, 16'h5452, 16'h5453, 16'h5454, 16'h5455, 16'h5456, 16'h5457 	:	val_out <= 16'hf06b;
         16'h5458, 16'h5459, 16'h545a, 16'h545b, 16'h545c, 16'h545d, 16'h545e, 16'h545f 	:	val_out <= 16'hf05f;
         16'h5460, 16'h5461, 16'h5462, 16'h5463, 16'h5464, 16'h5465, 16'h5466, 16'h5467 	:	val_out <= 16'hf053;
         16'h5468, 16'h5469, 16'h546a, 16'h546b, 16'h546c, 16'h546d, 16'h546e, 16'h546f 	:	val_out <= 16'hf047;
         16'h5470, 16'h5471, 16'h5472, 16'h5473, 16'h5474, 16'h5475, 16'h5476, 16'h5477 	:	val_out <= 16'hf03b;
         16'h5478, 16'h5479, 16'h547a, 16'h547b, 16'h547c, 16'h547d, 16'h547e, 16'h547f 	:	val_out <= 16'hf02f;
         16'h5480, 16'h5481, 16'h5482, 16'h5483, 16'h5484, 16'h5485, 16'h5486, 16'h5487 	:	val_out <= 16'hf023;
         16'h5488, 16'h5489, 16'h548a, 16'h548b, 16'h548c, 16'h548d, 16'h548e, 16'h548f 	:	val_out <= 16'hf016;
         16'h5490, 16'h5491, 16'h5492, 16'h5493, 16'h5494, 16'h5495, 16'h5496, 16'h5497 	:	val_out <= 16'hf00a;
         16'h5498, 16'h5499, 16'h549a, 16'h549b, 16'h549c, 16'h549d, 16'h549e, 16'h549f 	:	val_out <= 16'heffe;
         16'h54a0, 16'h54a1, 16'h54a2, 16'h54a3, 16'h54a4, 16'h54a5, 16'h54a6, 16'h54a7 	:	val_out <= 16'heff2;
         16'h54a8, 16'h54a9, 16'h54aa, 16'h54ab, 16'h54ac, 16'h54ad, 16'h54ae, 16'h54af 	:	val_out <= 16'hefe6;
         16'h54b0, 16'h54b1, 16'h54b2, 16'h54b3, 16'h54b4, 16'h54b5, 16'h54b6, 16'h54b7 	:	val_out <= 16'hefda;
         16'h54b8, 16'h54b9, 16'h54ba, 16'h54bb, 16'h54bc, 16'h54bd, 16'h54be, 16'h54bf 	:	val_out <= 16'hefcd;
         16'h54c0, 16'h54c1, 16'h54c2, 16'h54c3, 16'h54c4, 16'h54c5, 16'h54c6, 16'h54c7 	:	val_out <= 16'hefc1;
         16'h54c8, 16'h54c9, 16'h54ca, 16'h54cb, 16'h54cc, 16'h54cd, 16'h54ce, 16'h54cf 	:	val_out <= 16'hefb5;
         16'h54d0, 16'h54d1, 16'h54d2, 16'h54d3, 16'h54d4, 16'h54d5, 16'h54d6, 16'h54d7 	:	val_out <= 16'hefa9;
         16'h54d8, 16'h54d9, 16'h54da, 16'h54db, 16'h54dc, 16'h54dd, 16'h54de, 16'h54df 	:	val_out <= 16'hef9c;
         16'h54e0, 16'h54e1, 16'h54e2, 16'h54e3, 16'h54e4, 16'h54e5, 16'h54e6, 16'h54e7 	:	val_out <= 16'hef90;
         16'h54e8, 16'h54e9, 16'h54ea, 16'h54eb, 16'h54ec, 16'h54ed, 16'h54ee, 16'h54ef 	:	val_out <= 16'hef84;
         16'h54f0, 16'h54f1, 16'h54f2, 16'h54f3, 16'h54f4, 16'h54f5, 16'h54f6, 16'h54f7 	:	val_out <= 16'hef77;
         16'h54f8, 16'h54f9, 16'h54fa, 16'h54fb, 16'h54fc, 16'h54fd, 16'h54fe, 16'h54ff 	:	val_out <= 16'hef6b;
         16'h5500, 16'h5501, 16'h5502, 16'h5503, 16'h5504, 16'h5505, 16'h5506, 16'h5507 	:	val_out <= 16'hef5f;
         16'h5508, 16'h5509, 16'h550a, 16'h550b, 16'h550c, 16'h550d, 16'h550e, 16'h550f 	:	val_out <= 16'hef52;
         16'h5510, 16'h5511, 16'h5512, 16'h5513, 16'h5514, 16'h5515, 16'h5516, 16'h5517 	:	val_out <= 16'hef46;
         16'h5518, 16'h5519, 16'h551a, 16'h551b, 16'h551c, 16'h551d, 16'h551e, 16'h551f 	:	val_out <= 16'hef39;
         16'h5520, 16'h5521, 16'h5522, 16'h5523, 16'h5524, 16'h5525, 16'h5526, 16'h5527 	:	val_out <= 16'hef2d;
         16'h5528, 16'h5529, 16'h552a, 16'h552b, 16'h552c, 16'h552d, 16'h552e, 16'h552f 	:	val_out <= 16'hef20;
         16'h5530, 16'h5531, 16'h5532, 16'h5533, 16'h5534, 16'h5535, 16'h5536, 16'h5537 	:	val_out <= 16'hef14;
         16'h5538, 16'h5539, 16'h553a, 16'h553b, 16'h553c, 16'h553d, 16'h553e, 16'h553f 	:	val_out <= 16'hef07;
         16'h5540, 16'h5541, 16'h5542, 16'h5543, 16'h5544, 16'h5545, 16'h5546, 16'h5547 	:	val_out <= 16'heefb;
         16'h5548, 16'h5549, 16'h554a, 16'h554b, 16'h554c, 16'h554d, 16'h554e, 16'h554f 	:	val_out <= 16'heeee;
         16'h5550, 16'h5551, 16'h5552, 16'h5553, 16'h5554, 16'h5555, 16'h5556, 16'h5557 	:	val_out <= 16'heee2;
         16'h5558, 16'h5559, 16'h555a, 16'h555b, 16'h555c, 16'h555d, 16'h555e, 16'h555f 	:	val_out <= 16'heed5;
         16'h5560, 16'h5561, 16'h5562, 16'h5563, 16'h5564, 16'h5565, 16'h5566, 16'h5567 	:	val_out <= 16'heec9;
         16'h5568, 16'h5569, 16'h556a, 16'h556b, 16'h556c, 16'h556d, 16'h556e, 16'h556f 	:	val_out <= 16'heebc;
         16'h5570, 16'h5571, 16'h5572, 16'h5573, 16'h5574, 16'h5575, 16'h5576, 16'h5577 	:	val_out <= 16'heeaf;
         16'h5578, 16'h5579, 16'h557a, 16'h557b, 16'h557c, 16'h557d, 16'h557e, 16'h557f 	:	val_out <= 16'heea3;
         16'h5580, 16'h5581, 16'h5582, 16'h5583, 16'h5584, 16'h5585, 16'h5586, 16'h5587 	:	val_out <= 16'hee96;
         16'h5588, 16'h5589, 16'h558a, 16'h558b, 16'h558c, 16'h558d, 16'h558e, 16'h558f 	:	val_out <= 16'hee89;
         16'h5590, 16'h5591, 16'h5592, 16'h5593, 16'h5594, 16'h5595, 16'h5596, 16'h5597 	:	val_out <= 16'hee7d;
         16'h5598, 16'h5599, 16'h559a, 16'h559b, 16'h559c, 16'h559d, 16'h559e, 16'h559f 	:	val_out <= 16'hee70;
         16'h55a0, 16'h55a1, 16'h55a2, 16'h55a3, 16'h55a4, 16'h55a5, 16'h55a6, 16'h55a7 	:	val_out <= 16'hee63;
         16'h55a8, 16'h55a9, 16'h55aa, 16'h55ab, 16'h55ac, 16'h55ad, 16'h55ae, 16'h55af 	:	val_out <= 16'hee57;
         16'h55b0, 16'h55b1, 16'h55b2, 16'h55b3, 16'h55b4, 16'h55b5, 16'h55b6, 16'h55b7 	:	val_out <= 16'hee4a;
         16'h55b8, 16'h55b9, 16'h55ba, 16'h55bb, 16'h55bc, 16'h55bd, 16'h55be, 16'h55bf 	:	val_out <= 16'hee3d;
         16'h55c0, 16'h55c1, 16'h55c2, 16'h55c3, 16'h55c4, 16'h55c5, 16'h55c6, 16'h55c7 	:	val_out <= 16'hee30;
         16'h55c8, 16'h55c9, 16'h55ca, 16'h55cb, 16'h55cc, 16'h55cd, 16'h55ce, 16'h55cf 	:	val_out <= 16'hee24;
         16'h55d0, 16'h55d1, 16'h55d2, 16'h55d3, 16'h55d4, 16'h55d5, 16'h55d6, 16'h55d7 	:	val_out <= 16'hee17;
         16'h55d8, 16'h55d9, 16'h55da, 16'h55db, 16'h55dc, 16'h55dd, 16'h55de, 16'h55df 	:	val_out <= 16'hee0a;
         16'h55e0, 16'h55e1, 16'h55e2, 16'h55e3, 16'h55e4, 16'h55e5, 16'h55e6, 16'h55e7 	:	val_out <= 16'hedfd;
         16'h55e8, 16'h55e9, 16'h55ea, 16'h55eb, 16'h55ec, 16'h55ed, 16'h55ee, 16'h55ef 	:	val_out <= 16'hedf0;
         16'h55f0, 16'h55f1, 16'h55f2, 16'h55f3, 16'h55f4, 16'h55f5, 16'h55f6, 16'h55f7 	:	val_out <= 16'hede3;
         16'h55f8, 16'h55f9, 16'h55fa, 16'h55fb, 16'h55fc, 16'h55fd, 16'h55fe, 16'h55ff 	:	val_out <= 16'hedd6;
         16'h5600, 16'h5601, 16'h5602, 16'h5603, 16'h5604, 16'h5605, 16'h5606, 16'h5607 	:	val_out <= 16'hedca;
         16'h5608, 16'h5609, 16'h560a, 16'h560b, 16'h560c, 16'h560d, 16'h560e, 16'h560f 	:	val_out <= 16'hedbd;
         16'h5610, 16'h5611, 16'h5612, 16'h5613, 16'h5614, 16'h5615, 16'h5616, 16'h5617 	:	val_out <= 16'hedb0;
         16'h5618, 16'h5619, 16'h561a, 16'h561b, 16'h561c, 16'h561d, 16'h561e, 16'h561f 	:	val_out <= 16'heda3;
         16'h5620, 16'h5621, 16'h5622, 16'h5623, 16'h5624, 16'h5625, 16'h5626, 16'h5627 	:	val_out <= 16'hed96;
         16'h5628, 16'h5629, 16'h562a, 16'h562b, 16'h562c, 16'h562d, 16'h562e, 16'h562f 	:	val_out <= 16'hed89;
         16'h5630, 16'h5631, 16'h5632, 16'h5633, 16'h5634, 16'h5635, 16'h5636, 16'h5637 	:	val_out <= 16'hed7c;
         16'h5638, 16'h5639, 16'h563a, 16'h563b, 16'h563c, 16'h563d, 16'h563e, 16'h563f 	:	val_out <= 16'hed6f;
         16'h5640, 16'h5641, 16'h5642, 16'h5643, 16'h5644, 16'h5645, 16'h5646, 16'h5647 	:	val_out <= 16'hed62;
         16'h5648, 16'h5649, 16'h564a, 16'h564b, 16'h564c, 16'h564d, 16'h564e, 16'h564f 	:	val_out <= 16'hed55;
         16'h5650, 16'h5651, 16'h5652, 16'h5653, 16'h5654, 16'h5655, 16'h5656, 16'h5657 	:	val_out <= 16'hed48;
         16'h5658, 16'h5659, 16'h565a, 16'h565b, 16'h565c, 16'h565d, 16'h565e, 16'h565f 	:	val_out <= 16'hed3a;
         16'h5660, 16'h5661, 16'h5662, 16'h5663, 16'h5664, 16'h5665, 16'h5666, 16'h5667 	:	val_out <= 16'hed2d;
         16'h5668, 16'h5669, 16'h566a, 16'h566b, 16'h566c, 16'h566d, 16'h566e, 16'h566f 	:	val_out <= 16'hed20;
         16'h5670, 16'h5671, 16'h5672, 16'h5673, 16'h5674, 16'h5675, 16'h5676, 16'h5677 	:	val_out <= 16'hed13;
         16'h5678, 16'h5679, 16'h567a, 16'h567b, 16'h567c, 16'h567d, 16'h567e, 16'h567f 	:	val_out <= 16'hed06;
         16'h5680, 16'h5681, 16'h5682, 16'h5683, 16'h5684, 16'h5685, 16'h5686, 16'h5687 	:	val_out <= 16'hecf9;
         16'h5688, 16'h5689, 16'h568a, 16'h568b, 16'h568c, 16'h568d, 16'h568e, 16'h568f 	:	val_out <= 16'hecec;
         16'h5690, 16'h5691, 16'h5692, 16'h5693, 16'h5694, 16'h5695, 16'h5696, 16'h5697 	:	val_out <= 16'hecde;
         16'h5698, 16'h5699, 16'h569a, 16'h569b, 16'h569c, 16'h569d, 16'h569e, 16'h569f 	:	val_out <= 16'hecd1;
         16'h56a0, 16'h56a1, 16'h56a2, 16'h56a3, 16'h56a4, 16'h56a5, 16'h56a6, 16'h56a7 	:	val_out <= 16'hecc4;
         16'h56a8, 16'h56a9, 16'h56aa, 16'h56ab, 16'h56ac, 16'h56ad, 16'h56ae, 16'h56af 	:	val_out <= 16'hecb7;
         16'h56b0, 16'h56b1, 16'h56b2, 16'h56b3, 16'h56b4, 16'h56b5, 16'h56b6, 16'h56b7 	:	val_out <= 16'heca9;
         16'h56b8, 16'h56b9, 16'h56ba, 16'h56bb, 16'h56bc, 16'h56bd, 16'h56be, 16'h56bf 	:	val_out <= 16'hec9c;
         16'h56c0, 16'h56c1, 16'h56c2, 16'h56c3, 16'h56c4, 16'h56c5, 16'h56c6, 16'h56c7 	:	val_out <= 16'hec8f;
         16'h56c8, 16'h56c9, 16'h56ca, 16'h56cb, 16'h56cc, 16'h56cd, 16'h56ce, 16'h56cf 	:	val_out <= 16'hec81;
         16'h56d0, 16'h56d1, 16'h56d2, 16'h56d3, 16'h56d4, 16'h56d5, 16'h56d6, 16'h56d7 	:	val_out <= 16'hec74;
         16'h56d8, 16'h56d9, 16'h56da, 16'h56db, 16'h56dc, 16'h56dd, 16'h56de, 16'h56df 	:	val_out <= 16'hec67;
         16'h56e0, 16'h56e1, 16'h56e2, 16'h56e3, 16'h56e4, 16'h56e5, 16'h56e6, 16'h56e7 	:	val_out <= 16'hec59;
         16'h56e8, 16'h56e9, 16'h56ea, 16'h56eb, 16'h56ec, 16'h56ed, 16'h56ee, 16'h56ef 	:	val_out <= 16'hec4c;
         16'h56f0, 16'h56f1, 16'h56f2, 16'h56f3, 16'h56f4, 16'h56f5, 16'h56f6, 16'h56f7 	:	val_out <= 16'hec3f;
         16'h56f8, 16'h56f9, 16'h56fa, 16'h56fb, 16'h56fc, 16'h56fd, 16'h56fe, 16'h56ff 	:	val_out <= 16'hec31;
         16'h5700, 16'h5701, 16'h5702, 16'h5703, 16'h5704, 16'h5705, 16'h5706, 16'h5707 	:	val_out <= 16'hec24;
         16'h5708, 16'h5709, 16'h570a, 16'h570b, 16'h570c, 16'h570d, 16'h570e, 16'h570f 	:	val_out <= 16'hec16;
         16'h5710, 16'h5711, 16'h5712, 16'h5713, 16'h5714, 16'h5715, 16'h5716, 16'h5717 	:	val_out <= 16'hec09;
         16'h5718, 16'h5719, 16'h571a, 16'h571b, 16'h571c, 16'h571d, 16'h571e, 16'h571f 	:	val_out <= 16'hebfb;
         16'h5720, 16'h5721, 16'h5722, 16'h5723, 16'h5724, 16'h5725, 16'h5726, 16'h5727 	:	val_out <= 16'hebee;
         16'h5728, 16'h5729, 16'h572a, 16'h572b, 16'h572c, 16'h572d, 16'h572e, 16'h572f 	:	val_out <= 16'hebe0;
         16'h5730, 16'h5731, 16'h5732, 16'h5733, 16'h5734, 16'h5735, 16'h5736, 16'h5737 	:	val_out <= 16'hebd3;
         16'h5738, 16'h5739, 16'h573a, 16'h573b, 16'h573c, 16'h573d, 16'h573e, 16'h573f 	:	val_out <= 16'hebc5;
         16'h5740, 16'h5741, 16'h5742, 16'h5743, 16'h5744, 16'h5745, 16'h5746, 16'h5747 	:	val_out <= 16'hebb8;
         16'h5748, 16'h5749, 16'h574a, 16'h574b, 16'h574c, 16'h574d, 16'h574e, 16'h574f 	:	val_out <= 16'hebaa;
         16'h5750, 16'h5751, 16'h5752, 16'h5753, 16'h5754, 16'h5755, 16'h5756, 16'h5757 	:	val_out <= 16'heb9c;
         16'h5758, 16'h5759, 16'h575a, 16'h575b, 16'h575c, 16'h575d, 16'h575e, 16'h575f 	:	val_out <= 16'heb8f;
         16'h5760, 16'h5761, 16'h5762, 16'h5763, 16'h5764, 16'h5765, 16'h5766, 16'h5767 	:	val_out <= 16'heb81;
         16'h5768, 16'h5769, 16'h576a, 16'h576b, 16'h576c, 16'h576d, 16'h576e, 16'h576f 	:	val_out <= 16'heb73;
         16'h5770, 16'h5771, 16'h5772, 16'h5773, 16'h5774, 16'h5775, 16'h5776, 16'h5777 	:	val_out <= 16'heb66;
         16'h5778, 16'h5779, 16'h577a, 16'h577b, 16'h577c, 16'h577d, 16'h577e, 16'h577f 	:	val_out <= 16'heb58;
         16'h5780, 16'h5781, 16'h5782, 16'h5783, 16'h5784, 16'h5785, 16'h5786, 16'h5787 	:	val_out <= 16'heb4a;
         16'h5788, 16'h5789, 16'h578a, 16'h578b, 16'h578c, 16'h578d, 16'h578e, 16'h578f 	:	val_out <= 16'heb3d;
         16'h5790, 16'h5791, 16'h5792, 16'h5793, 16'h5794, 16'h5795, 16'h5796, 16'h5797 	:	val_out <= 16'heb2f;
         16'h5798, 16'h5799, 16'h579a, 16'h579b, 16'h579c, 16'h579d, 16'h579e, 16'h579f 	:	val_out <= 16'heb21;
         16'h57a0, 16'h57a1, 16'h57a2, 16'h57a3, 16'h57a4, 16'h57a5, 16'h57a6, 16'h57a7 	:	val_out <= 16'heb13;
         16'h57a8, 16'h57a9, 16'h57aa, 16'h57ab, 16'h57ac, 16'h57ad, 16'h57ae, 16'h57af 	:	val_out <= 16'heb06;
         16'h57b0, 16'h57b1, 16'h57b2, 16'h57b3, 16'h57b4, 16'h57b5, 16'h57b6, 16'h57b7 	:	val_out <= 16'heaf8;
         16'h57b8, 16'h57b9, 16'h57ba, 16'h57bb, 16'h57bc, 16'h57bd, 16'h57be, 16'h57bf 	:	val_out <= 16'heaea;
         16'h57c0, 16'h57c1, 16'h57c2, 16'h57c3, 16'h57c4, 16'h57c5, 16'h57c6, 16'h57c7 	:	val_out <= 16'headc;
         16'h57c8, 16'h57c9, 16'h57ca, 16'h57cb, 16'h57cc, 16'h57cd, 16'h57ce, 16'h57cf 	:	val_out <= 16'heace;
         16'h57d0, 16'h57d1, 16'h57d2, 16'h57d3, 16'h57d4, 16'h57d5, 16'h57d6, 16'h57d7 	:	val_out <= 16'heac1;
         16'h57d8, 16'h57d9, 16'h57da, 16'h57db, 16'h57dc, 16'h57dd, 16'h57de, 16'h57df 	:	val_out <= 16'heab3;
         16'h57e0, 16'h57e1, 16'h57e2, 16'h57e3, 16'h57e4, 16'h57e5, 16'h57e6, 16'h57e7 	:	val_out <= 16'heaa5;
         16'h57e8, 16'h57e9, 16'h57ea, 16'h57eb, 16'h57ec, 16'h57ed, 16'h57ee, 16'h57ef 	:	val_out <= 16'hea97;
         16'h57f0, 16'h57f1, 16'h57f2, 16'h57f3, 16'h57f4, 16'h57f5, 16'h57f6, 16'h57f7 	:	val_out <= 16'hea89;
         16'h57f8, 16'h57f9, 16'h57fa, 16'h57fb, 16'h57fc, 16'h57fd, 16'h57fe, 16'h57ff 	:	val_out <= 16'hea7b;
         16'h5800, 16'h5801, 16'h5802, 16'h5803, 16'h5804, 16'h5805, 16'h5806, 16'h5807 	:	val_out <= 16'hea6d;
         16'h5808, 16'h5809, 16'h580a, 16'h580b, 16'h580c, 16'h580d, 16'h580e, 16'h580f 	:	val_out <= 16'hea5f;
         16'h5810, 16'h5811, 16'h5812, 16'h5813, 16'h5814, 16'h5815, 16'h5816, 16'h5817 	:	val_out <= 16'hea51;
         16'h5818, 16'h5819, 16'h581a, 16'h581b, 16'h581c, 16'h581d, 16'h581e, 16'h581f 	:	val_out <= 16'hea43;
         16'h5820, 16'h5821, 16'h5822, 16'h5823, 16'h5824, 16'h5825, 16'h5826, 16'h5827 	:	val_out <= 16'hea35;
         16'h5828, 16'h5829, 16'h582a, 16'h582b, 16'h582c, 16'h582d, 16'h582e, 16'h582f 	:	val_out <= 16'hea27;
         16'h5830, 16'h5831, 16'h5832, 16'h5833, 16'h5834, 16'h5835, 16'h5836, 16'h5837 	:	val_out <= 16'hea19;
         16'h5838, 16'h5839, 16'h583a, 16'h583b, 16'h583c, 16'h583d, 16'h583e, 16'h583f 	:	val_out <= 16'hea0b;
         16'h5840, 16'h5841, 16'h5842, 16'h5843, 16'h5844, 16'h5845, 16'h5846, 16'h5847 	:	val_out <= 16'he9fd;
         16'h5848, 16'h5849, 16'h584a, 16'h584b, 16'h584c, 16'h584d, 16'h584e, 16'h584f 	:	val_out <= 16'he9ef;
         16'h5850, 16'h5851, 16'h5852, 16'h5853, 16'h5854, 16'h5855, 16'h5856, 16'h5857 	:	val_out <= 16'he9e1;
         16'h5858, 16'h5859, 16'h585a, 16'h585b, 16'h585c, 16'h585d, 16'h585e, 16'h585f 	:	val_out <= 16'he9d3;
         16'h5860, 16'h5861, 16'h5862, 16'h5863, 16'h5864, 16'h5865, 16'h5866, 16'h5867 	:	val_out <= 16'he9c4;
         16'h5868, 16'h5869, 16'h586a, 16'h586b, 16'h586c, 16'h586d, 16'h586e, 16'h586f 	:	val_out <= 16'he9b6;
         16'h5870, 16'h5871, 16'h5872, 16'h5873, 16'h5874, 16'h5875, 16'h5876, 16'h5877 	:	val_out <= 16'he9a8;
         16'h5878, 16'h5879, 16'h587a, 16'h587b, 16'h587c, 16'h587d, 16'h587e, 16'h587f 	:	val_out <= 16'he99a;
         16'h5880, 16'h5881, 16'h5882, 16'h5883, 16'h5884, 16'h5885, 16'h5886, 16'h5887 	:	val_out <= 16'he98c;
         16'h5888, 16'h5889, 16'h588a, 16'h588b, 16'h588c, 16'h588d, 16'h588e, 16'h588f 	:	val_out <= 16'he97d;
         16'h5890, 16'h5891, 16'h5892, 16'h5893, 16'h5894, 16'h5895, 16'h5896, 16'h5897 	:	val_out <= 16'he96f;
         16'h5898, 16'h5899, 16'h589a, 16'h589b, 16'h589c, 16'h589d, 16'h589e, 16'h589f 	:	val_out <= 16'he961;
         16'h58a0, 16'h58a1, 16'h58a2, 16'h58a3, 16'h58a4, 16'h58a5, 16'h58a6, 16'h58a7 	:	val_out <= 16'he953;
         16'h58a8, 16'h58a9, 16'h58aa, 16'h58ab, 16'h58ac, 16'h58ad, 16'h58ae, 16'h58af 	:	val_out <= 16'he944;
         16'h58b0, 16'h58b1, 16'h58b2, 16'h58b3, 16'h58b4, 16'h58b5, 16'h58b6, 16'h58b7 	:	val_out <= 16'he936;
         16'h58b8, 16'h58b9, 16'h58ba, 16'h58bb, 16'h58bc, 16'h58bd, 16'h58be, 16'h58bf 	:	val_out <= 16'he928;
         16'h58c0, 16'h58c1, 16'h58c2, 16'h58c3, 16'h58c4, 16'h58c5, 16'h58c6, 16'h58c7 	:	val_out <= 16'he919;
         16'h58c8, 16'h58c9, 16'h58ca, 16'h58cb, 16'h58cc, 16'h58cd, 16'h58ce, 16'h58cf 	:	val_out <= 16'he90b;
         16'h58d0, 16'h58d1, 16'h58d2, 16'h58d3, 16'h58d4, 16'h58d5, 16'h58d6, 16'h58d7 	:	val_out <= 16'he8fd;
         16'h58d8, 16'h58d9, 16'h58da, 16'h58db, 16'h58dc, 16'h58dd, 16'h58de, 16'h58df 	:	val_out <= 16'he8ee;
         16'h58e0, 16'h58e1, 16'h58e2, 16'h58e3, 16'h58e4, 16'h58e5, 16'h58e6, 16'h58e7 	:	val_out <= 16'he8e0;
         16'h58e8, 16'h58e9, 16'h58ea, 16'h58eb, 16'h58ec, 16'h58ed, 16'h58ee, 16'h58ef 	:	val_out <= 16'he8d1;
         16'h58f0, 16'h58f1, 16'h58f2, 16'h58f3, 16'h58f4, 16'h58f5, 16'h58f6, 16'h58f7 	:	val_out <= 16'he8c3;
         16'h58f8, 16'h58f9, 16'h58fa, 16'h58fb, 16'h58fc, 16'h58fd, 16'h58fe, 16'h58ff 	:	val_out <= 16'he8b5;
         16'h5900, 16'h5901, 16'h5902, 16'h5903, 16'h5904, 16'h5905, 16'h5906, 16'h5907 	:	val_out <= 16'he8a6;
         16'h5908, 16'h5909, 16'h590a, 16'h590b, 16'h590c, 16'h590d, 16'h590e, 16'h590f 	:	val_out <= 16'he898;
         16'h5910, 16'h5911, 16'h5912, 16'h5913, 16'h5914, 16'h5915, 16'h5916, 16'h5917 	:	val_out <= 16'he889;
         16'h5918, 16'h5919, 16'h591a, 16'h591b, 16'h591c, 16'h591d, 16'h591e, 16'h591f 	:	val_out <= 16'he87b;
         16'h5920, 16'h5921, 16'h5922, 16'h5923, 16'h5924, 16'h5925, 16'h5926, 16'h5927 	:	val_out <= 16'he86c;
         16'h5928, 16'h5929, 16'h592a, 16'h592b, 16'h592c, 16'h592d, 16'h592e, 16'h592f 	:	val_out <= 16'he85e;
         16'h5930, 16'h5931, 16'h5932, 16'h5933, 16'h5934, 16'h5935, 16'h5936, 16'h5937 	:	val_out <= 16'he84f;
         16'h5938, 16'h5939, 16'h593a, 16'h593b, 16'h593c, 16'h593d, 16'h593e, 16'h593f 	:	val_out <= 16'he840;
         16'h5940, 16'h5941, 16'h5942, 16'h5943, 16'h5944, 16'h5945, 16'h5946, 16'h5947 	:	val_out <= 16'he832;
         16'h5948, 16'h5949, 16'h594a, 16'h594b, 16'h594c, 16'h594d, 16'h594e, 16'h594f 	:	val_out <= 16'he823;
         16'h5950, 16'h5951, 16'h5952, 16'h5953, 16'h5954, 16'h5955, 16'h5956, 16'h5957 	:	val_out <= 16'he815;
         16'h5958, 16'h5959, 16'h595a, 16'h595b, 16'h595c, 16'h595d, 16'h595e, 16'h595f 	:	val_out <= 16'he806;
         16'h5960, 16'h5961, 16'h5962, 16'h5963, 16'h5964, 16'h5965, 16'h5966, 16'h5967 	:	val_out <= 16'he7f7;
         16'h5968, 16'h5969, 16'h596a, 16'h596b, 16'h596c, 16'h596d, 16'h596e, 16'h596f 	:	val_out <= 16'he7e9;
         16'h5970, 16'h5971, 16'h5972, 16'h5973, 16'h5974, 16'h5975, 16'h5976, 16'h5977 	:	val_out <= 16'he7da;
         16'h5978, 16'h5979, 16'h597a, 16'h597b, 16'h597c, 16'h597d, 16'h597e, 16'h597f 	:	val_out <= 16'he7cb;
         16'h5980, 16'h5981, 16'h5982, 16'h5983, 16'h5984, 16'h5985, 16'h5986, 16'h5987 	:	val_out <= 16'he7bd;
         16'h5988, 16'h5989, 16'h598a, 16'h598b, 16'h598c, 16'h598d, 16'h598e, 16'h598f 	:	val_out <= 16'he7ae;
         16'h5990, 16'h5991, 16'h5992, 16'h5993, 16'h5994, 16'h5995, 16'h5996, 16'h5997 	:	val_out <= 16'he79f;
         16'h5998, 16'h5999, 16'h599a, 16'h599b, 16'h599c, 16'h599d, 16'h599e, 16'h599f 	:	val_out <= 16'he790;
         16'h59a0, 16'h59a1, 16'h59a2, 16'h59a3, 16'h59a4, 16'h59a5, 16'h59a6, 16'h59a7 	:	val_out <= 16'he782;
         16'h59a8, 16'h59a9, 16'h59aa, 16'h59ab, 16'h59ac, 16'h59ad, 16'h59ae, 16'h59af 	:	val_out <= 16'he773;
         16'h59b0, 16'h59b1, 16'h59b2, 16'h59b3, 16'h59b4, 16'h59b5, 16'h59b6, 16'h59b7 	:	val_out <= 16'he764;
         16'h59b8, 16'h59b9, 16'h59ba, 16'h59bb, 16'h59bc, 16'h59bd, 16'h59be, 16'h59bf 	:	val_out <= 16'he755;
         16'h59c0, 16'h59c1, 16'h59c2, 16'h59c3, 16'h59c4, 16'h59c5, 16'h59c6, 16'h59c7 	:	val_out <= 16'he746;
         16'h59c8, 16'h59c9, 16'h59ca, 16'h59cb, 16'h59cc, 16'h59cd, 16'h59ce, 16'h59cf 	:	val_out <= 16'he737;
         16'h59d0, 16'h59d1, 16'h59d2, 16'h59d3, 16'h59d4, 16'h59d5, 16'h59d6, 16'h59d7 	:	val_out <= 16'he729;
         16'h59d8, 16'h59d9, 16'h59da, 16'h59db, 16'h59dc, 16'h59dd, 16'h59de, 16'h59df 	:	val_out <= 16'he71a;
         16'h59e0, 16'h59e1, 16'h59e2, 16'h59e3, 16'h59e4, 16'h59e5, 16'h59e6, 16'h59e7 	:	val_out <= 16'he70b;
         16'h59e8, 16'h59e9, 16'h59ea, 16'h59eb, 16'h59ec, 16'h59ed, 16'h59ee, 16'h59ef 	:	val_out <= 16'he6fc;
         16'h59f0, 16'h59f1, 16'h59f2, 16'h59f3, 16'h59f4, 16'h59f5, 16'h59f6, 16'h59f7 	:	val_out <= 16'he6ed;
         16'h59f8, 16'h59f9, 16'h59fa, 16'h59fb, 16'h59fc, 16'h59fd, 16'h59fe, 16'h59ff 	:	val_out <= 16'he6de;
         16'h5a00, 16'h5a01, 16'h5a02, 16'h5a03, 16'h5a04, 16'h5a05, 16'h5a06, 16'h5a07 	:	val_out <= 16'he6cf;
         16'h5a08, 16'h5a09, 16'h5a0a, 16'h5a0b, 16'h5a0c, 16'h5a0d, 16'h5a0e, 16'h5a0f 	:	val_out <= 16'he6c0;
         16'h5a10, 16'h5a11, 16'h5a12, 16'h5a13, 16'h5a14, 16'h5a15, 16'h5a16, 16'h5a17 	:	val_out <= 16'he6b1;
         16'h5a18, 16'h5a19, 16'h5a1a, 16'h5a1b, 16'h5a1c, 16'h5a1d, 16'h5a1e, 16'h5a1f 	:	val_out <= 16'he6a2;
         16'h5a20, 16'h5a21, 16'h5a22, 16'h5a23, 16'h5a24, 16'h5a25, 16'h5a26, 16'h5a27 	:	val_out <= 16'he693;
         16'h5a28, 16'h5a29, 16'h5a2a, 16'h5a2b, 16'h5a2c, 16'h5a2d, 16'h5a2e, 16'h5a2f 	:	val_out <= 16'he684;
         16'h5a30, 16'h5a31, 16'h5a32, 16'h5a33, 16'h5a34, 16'h5a35, 16'h5a36, 16'h5a37 	:	val_out <= 16'he675;
         16'h5a38, 16'h5a39, 16'h5a3a, 16'h5a3b, 16'h5a3c, 16'h5a3d, 16'h5a3e, 16'h5a3f 	:	val_out <= 16'he666;
         16'h5a40, 16'h5a41, 16'h5a42, 16'h5a43, 16'h5a44, 16'h5a45, 16'h5a46, 16'h5a47 	:	val_out <= 16'he657;
         16'h5a48, 16'h5a49, 16'h5a4a, 16'h5a4b, 16'h5a4c, 16'h5a4d, 16'h5a4e, 16'h5a4f 	:	val_out <= 16'he648;
         16'h5a50, 16'h5a51, 16'h5a52, 16'h5a53, 16'h5a54, 16'h5a55, 16'h5a56, 16'h5a57 	:	val_out <= 16'he639;
         16'h5a58, 16'h5a59, 16'h5a5a, 16'h5a5b, 16'h5a5c, 16'h5a5d, 16'h5a5e, 16'h5a5f 	:	val_out <= 16'he629;
         16'h5a60, 16'h5a61, 16'h5a62, 16'h5a63, 16'h5a64, 16'h5a65, 16'h5a66, 16'h5a67 	:	val_out <= 16'he61a;
         16'h5a68, 16'h5a69, 16'h5a6a, 16'h5a6b, 16'h5a6c, 16'h5a6d, 16'h5a6e, 16'h5a6f 	:	val_out <= 16'he60b;
         16'h5a70, 16'h5a71, 16'h5a72, 16'h5a73, 16'h5a74, 16'h5a75, 16'h5a76, 16'h5a77 	:	val_out <= 16'he5fc;
         16'h5a78, 16'h5a79, 16'h5a7a, 16'h5a7b, 16'h5a7c, 16'h5a7d, 16'h5a7e, 16'h5a7f 	:	val_out <= 16'he5ed;
         16'h5a80, 16'h5a81, 16'h5a82, 16'h5a83, 16'h5a84, 16'h5a85, 16'h5a86, 16'h5a87 	:	val_out <= 16'he5dd;
         16'h5a88, 16'h5a89, 16'h5a8a, 16'h5a8b, 16'h5a8c, 16'h5a8d, 16'h5a8e, 16'h5a8f 	:	val_out <= 16'he5ce;
         16'h5a90, 16'h5a91, 16'h5a92, 16'h5a93, 16'h5a94, 16'h5a95, 16'h5a96, 16'h5a97 	:	val_out <= 16'he5bf;
         16'h5a98, 16'h5a99, 16'h5a9a, 16'h5a9b, 16'h5a9c, 16'h5a9d, 16'h5a9e, 16'h5a9f 	:	val_out <= 16'he5b0;
         16'h5aa0, 16'h5aa1, 16'h5aa2, 16'h5aa3, 16'h5aa4, 16'h5aa5, 16'h5aa6, 16'h5aa7 	:	val_out <= 16'he5a0;
         16'h5aa8, 16'h5aa9, 16'h5aaa, 16'h5aab, 16'h5aac, 16'h5aad, 16'h5aae, 16'h5aaf 	:	val_out <= 16'he591;
         16'h5ab0, 16'h5ab1, 16'h5ab2, 16'h5ab3, 16'h5ab4, 16'h5ab5, 16'h5ab6, 16'h5ab7 	:	val_out <= 16'he582;
         16'h5ab8, 16'h5ab9, 16'h5aba, 16'h5abb, 16'h5abc, 16'h5abd, 16'h5abe, 16'h5abf 	:	val_out <= 16'he573;
         16'h5ac0, 16'h5ac1, 16'h5ac2, 16'h5ac3, 16'h5ac4, 16'h5ac5, 16'h5ac6, 16'h5ac7 	:	val_out <= 16'he563;
         16'h5ac8, 16'h5ac9, 16'h5aca, 16'h5acb, 16'h5acc, 16'h5acd, 16'h5ace, 16'h5acf 	:	val_out <= 16'he554;
         16'h5ad0, 16'h5ad1, 16'h5ad2, 16'h5ad3, 16'h5ad4, 16'h5ad5, 16'h5ad6, 16'h5ad7 	:	val_out <= 16'he545;
         16'h5ad8, 16'h5ad9, 16'h5ada, 16'h5adb, 16'h5adc, 16'h5add, 16'h5ade, 16'h5adf 	:	val_out <= 16'he535;
         16'h5ae0, 16'h5ae1, 16'h5ae2, 16'h5ae3, 16'h5ae4, 16'h5ae5, 16'h5ae6, 16'h5ae7 	:	val_out <= 16'he526;
         16'h5ae8, 16'h5ae9, 16'h5aea, 16'h5aeb, 16'h5aec, 16'h5aed, 16'h5aee, 16'h5aef 	:	val_out <= 16'he516;
         16'h5af0, 16'h5af1, 16'h5af2, 16'h5af3, 16'h5af4, 16'h5af5, 16'h5af6, 16'h5af7 	:	val_out <= 16'he507;
         16'h5af8, 16'h5af9, 16'h5afa, 16'h5afb, 16'h5afc, 16'h5afd, 16'h5afe, 16'h5aff 	:	val_out <= 16'he4f7;
         16'h5b00, 16'h5b01, 16'h5b02, 16'h5b03, 16'h5b04, 16'h5b05, 16'h5b06, 16'h5b07 	:	val_out <= 16'he4e8;
         16'h5b08, 16'h5b09, 16'h5b0a, 16'h5b0b, 16'h5b0c, 16'h5b0d, 16'h5b0e, 16'h5b0f 	:	val_out <= 16'he4d9;
         16'h5b10, 16'h5b11, 16'h5b12, 16'h5b13, 16'h5b14, 16'h5b15, 16'h5b16, 16'h5b17 	:	val_out <= 16'he4c9;
         16'h5b18, 16'h5b19, 16'h5b1a, 16'h5b1b, 16'h5b1c, 16'h5b1d, 16'h5b1e, 16'h5b1f 	:	val_out <= 16'he4ba;
         16'h5b20, 16'h5b21, 16'h5b22, 16'h5b23, 16'h5b24, 16'h5b25, 16'h5b26, 16'h5b27 	:	val_out <= 16'he4aa;
         16'h5b28, 16'h5b29, 16'h5b2a, 16'h5b2b, 16'h5b2c, 16'h5b2d, 16'h5b2e, 16'h5b2f 	:	val_out <= 16'he49b;
         16'h5b30, 16'h5b31, 16'h5b32, 16'h5b33, 16'h5b34, 16'h5b35, 16'h5b36, 16'h5b37 	:	val_out <= 16'he48b;
         16'h5b38, 16'h5b39, 16'h5b3a, 16'h5b3b, 16'h5b3c, 16'h5b3d, 16'h5b3e, 16'h5b3f 	:	val_out <= 16'he47b;
         16'h5b40, 16'h5b41, 16'h5b42, 16'h5b43, 16'h5b44, 16'h5b45, 16'h5b46, 16'h5b47 	:	val_out <= 16'he46c;
         16'h5b48, 16'h5b49, 16'h5b4a, 16'h5b4b, 16'h5b4c, 16'h5b4d, 16'h5b4e, 16'h5b4f 	:	val_out <= 16'he45c;
         16'h5b50, 16'h5b51, 16'h5b52, 16'h5b53, 16'h5b54, 16'h5b55, 16'h5b56, 16'h5b57 	:	val_out <= 16'he44d;
         16'h5b58, 16'h5b59, 16'h5b5a, 16'h5b5b, 16'h5b5c, 16'h5b5d, 16'h5b5e, 16'h5b5f 	:	val_out <= 16'he43d;
         16'h5b60, 16'h5b61, 16'h5b62, 16'h5b63, 16'h5b64, 16'h5b65, 16'h5b66, 16'h5b67 	:	val_out <= 16'he42d;
         16'h5b68, 16'h5b69, 16'h5b6a, 16'h5b6b, 16'h5b6c, 16'h5b6d, 16'h5b6e, 16'h5b6f 	:	val_out <= 16'he41e;
         16'h5b70, 16'h5b71, 16'h5b72, 16'h5b73, 16'h5b74, 16'h5b75, 16'h5b76, 16'h5b77 	:	val_out <= 16'he40e;
         16'h5b78, 16'h5b79, 16'h5b7a, 16'h5b7b, 16'h5b7c, 16'h5b7d, 16'h5b7e, 16'h5b7f 	:	val_out <= 16'he3fe;
         16'h5b80, 16'h5b81, 16'h5b82, 16'h5b83, 16'h5b84, 16'h5b85, 16'h5b86, 16'h5b87 	:	val_out <= 16'he3ef;
         16'h5b88, 16'h5b89, 16'h5b8a, 16'h5b8b, 16'h5b8c, 16'h5b8d, 16'h5b8e, 16'h5b8f 	:	val_out <= 16'he3df;
         16'h5b90, 16'h5b91, 16'h5b92, 16'h5b93, 16'h5b94, 16'h5b95, 16'h5b96, 16'h5b97 	:	val_out <= 16'he3cf;
         16'h5b98, 16'h5b99, 16'h5b9a, 16'h5b9b, 16'h5b9c, 16'h5b9d, 16'h5b9e, 16'h5b9f 	:	val_out <= 16'he3c0;
         16'h5ba0, 16'h5ba1, 16'h5ba2, 16'h5ba3, 16'h5ba4, 16'h5ba5, 16'h5ba6, 16'h5ba7 	:	val_out <= 16'he3b0;
         16'h5ba8, 16'h5ba9, 16'h5baa, 16'h5bab, 16'h5bac, 16'h5bad, 16'h5bae, 16'h5baf 	:	val_out <= 16'he3a0;
         16'h5bb0, 16'h5bb1, 16'h5bb2, 16'h5bb3, 16'h5bb4, 16'h5bb5, 16'h5bb6, 16'h5bb7 	:	val_out <= 16'he390;
         16'h5bb8, 16'h5bb9, 16'h5bba, 16'h5bbb, 16'h5bbc, 16'h5bbd, 16'h5bbe, 16'h5bbf 	:	val_out <= 16'he380;
         16'h5bc0, 16'h5bc1, 16'h5bc2, 16'h5bc3, 16'h5bc4, 16'h5bc5, 16'h5bc6, 16'h5bc7 	:	val_out <= 16'he371;
         16'h5bc8, 16'h5bc9, 16'h5bca, 16'h5bcb, 16'h5bcc, 16'h5bcd, 16'h5bce, 16'h5bcf 	:	val_out <= 16'he361;
         16'h5bd0, 16'h5bd1, 16'h5bd2, 16'h5bd3, 16'h5bd4, 16'h5bd5, 16'h5bd6, 16'h5bd7 	:	val_out <= 16'he351;
         16'h5bd8, 16'h5bd9, 16'h5bda, 16'h5bdb, 16'h5bdc, 16'h5bdd, 16'h5bde, 16'h5bdf 	:	val_out <= 16'he341;
         16'h5be0, 16'h5be1, 16'h5be2, 16'h5be3, 16'h5be4, 16'h5be5, 16'h5be6, 16'h5be7 	:	val_out <= 16'he331;
         16'h5be8, 16'h5be9, 16'h5bea, 16'h5beb, 16'h5bec, 16'h5bed, 16'h5bee, 16'h5bef 	:	val_out <= 16'he321;
         16'h5bf0, 16'h5bf1, 16'h5bf2, 16'h5bf3, 16'h5bf4, 16'h5bf5, 16'h5bf6, 16'h5bf7 	:	val_out <= 16'he311;
         16'h5bf8, 16'h5bf9, 16'h5bfa, 16'h5bfb, 16'h5bfc, 16'h5bfd, 16'h5bfe, 16'h5bff 	:	val_out <= 16'he301;
         16'h5c00, 16'h5c01, 16'h5c02, 16'h5c03, 16'h5c04, 16'h5c05, 16'h5c06, 16'h5c07 	:	val_out <= 16'he2f2;
         16'h5c08, 16'h5c09, 16'h5c0a, 16'h5c0b, 16'h5c0c, 16'h5c0d, 16'h5c0e, 16'h5c0f 	:	val_out <= 16'he2e2;
         16'h5c10, 16'h5c11, 16'h5c12, 16'h5c13, 16'h5c14, 16'h5c15, 16'h5c16, 16'h5c17 	:	val_out <= 16'he2d2;
         16'h5c18, 16'h5c19, 16'h5c1a, 16'h5c1b, 16'h5c1c, 16'h5c1d, 16'h5c1e, 16'h5c1f 	:	val_out <= 16'he2c2;
         16'h5c20, 16'h5c21, 16'h5c22, 16'h5c23, 16'h5c24, 16'h5c25, 16'h5c26, 16'h5c27 	:	val_out <= 16'he2b2;
         16'h5c28, 16'h5c29, 16'h5c2a, 16'h5c2b, 16'h5c2c, 16'h5c2d, 16'h5c2e, 16'h5c2f 	:	val_out <= 16'he2a2;
         16'h5c30, 16'h5c31, 16'h5c32, 16'h5c33, 16'h5c34, 16'h5c35, 16'h5c36, 16'h5c37 	:	val_out <= 16'he292;
         16'h5c38, 16'h5c39, 16'h5c3a, 16'h5c3b, 16'h5c3c, 16'h5c3d, 16'h5c3e, 16'h5c3f 	:	val_out <= 16'he282;
         16'h5c40, 16'h5c41, 16'h5c42, 16'h5c43, 16'h5c44, 16'h5c45, 16'h5c46, 16'h5c47 	:	val_out <= 16'he271;
         16'h5c48, 16'h5c49, 16'h5c4a, 16'h5c4b, 16'h5c4c, 16'h5c4d, 16'h5c4e, 16'h5c4f 	:	val_out <= 16'he261;
         16'h5c50, 16'h5c51, 16'h5c52, 16'h5c53, 16'h5c54, 16'h5c55, 16'h5c56, 16'h5c57 	:	val_out <= 16'he251;
         16'h5c58, 16'h5c59, 16'h5c5a, 16'h5c5b, 16'h5c5c, 16'h5c5d, 16'h5c5e, 16'h5c5f 	:	val_out <= 16'he241;
         16'h5c60, 16'h5c61, 16'h5c62, 16'h5c63, 16'h5c64, 16'h5c65, 16'h5c66, 16'h5c67 	:	val_out <= 16'he231;
         16'h5c68, 16'h5c69, 16'h5c6a, 16'h5c6b, 16'h5c6c, 16'h5c6d, 16'h5c6e, 16'h5c6f 	:	val_out <= 16'he221;
         16'h5c70, 16'h5c71, 16'h5c72, 16'h5c73, 16'h5c74, 16'h5c75, 16'h5c76, 16'h5c77 	:	val_out <= 16'he211;
         16'h5c78, 16'h5c79, 16'h5c7a, 16'h5c7b, 16'h5c7c, 16'h5c7d, 16'h5c7e, 16'h5c7f 	:	val_out <= 16'he201;
         16'h5c80, 16'h5c81, 16'h5c82, 16'h5c83, 16'h5c84, 16'h5c85, 16'h5c86, 16'h5c87 	:	val_out <= 16'he1f1;
         16'h5c88, 16'h5c89, 16'h5c8a, 16'h5c8b, 16'h5c8c, 16'h5c8d, 16'h5c8e, 16'h5c8f 	:	val_out <= 16'he1e0;
         16'h5c90, 16'h5c91, 16'h5c92, 16'h5c93, 16'h5c94, 16'h5c95, 16'h5c96, 16'h5c97 	:	val_out <= 16'he1d0;
         16'h5c98, 16'h5c99, 16'h5c9a, 16'h5c9b, 16'h5c9c, 16'h5c9d, 16'h5c9e, 16'h5c9f 	:	val_out <= 16'he1c0;
         16'h5ca0, 16'h5ca1, 16'h5ca2, 16'h5ca3, 16'h5ca4, 16'h5ca5, 16'h5ca6, 16'h5ca7 	:	val_out <= 16'he1b0;
         16'h5ca8, 16'h5ca9, 16'h5caa, 16'h5cab, 16'h5cac, 16'h5cad, 16'h5cae, 16'h5caf 	:	val_out <= 16'he19f;
         16'h5cb0, 16'h5cb1, 16'h5cb2, 16'h5cb3, 16'h5cb4, 16'h5cb5, 16'h5cb6, 16'h5cb7 	:	val_out <= 16'he18f;
         16'h5cb8, 16'h5cb9, 16'h5cba, 16'h5cbb, 16'h5cbc, 16'h5cbd, 16'h5cbe, 16'h5cbf 	:	val_out <= 16'he17f;
         16'h5cc0, 16'h5cc1, 16'h5cc2, 16'h5cc3, 16'h5cc4, 16'h5cc5, 16'h5cc6, 16'h5cc7 	:	val_out <= 16'he16f;
         16'h5cc8, 16'h5cc9, 16'h5cca, 16'h5ccb, 16'h5ccc, 16'h5ccd, 16'h5cce, 16'h5ccf 	:	val_out <= 16'he15e;
         16'h5cd0, 16'h5cd1, 16'h5cd2, 16'h5cd3, 16'h5cd4, 16'h5cd5, 16'h5cd6, 16'h5cd7 	:	val_out <= 16'he14e;
         16'h5cd8, 16'h5cd9, 16'h5cda, 16'h5cdb, 16'h5cdc, 16'h5cdd, 16'h5cde, 16'h5cdf 	:	val_out <= 16'he13e;
         16'h5ce0, 16'h5ce1, 16'h5ce2, 16'h5ce3, 16'h5ce4, 16'h5ce5, 16'h5ce6, 16'h5ce7 	:	val_out <= 16'he12d;
         16'h5ce8, 16'h5ce9, 16'h5cea, 16'h5ceb, 16'h5cec, 16'h5ced, 16'h5cee, 16'h5cef 	:	val_out <= 16'he11d;
         16'h5cf0, 16'h5cf1, 16'h5cf2, 16'h5cf3, 16'h5cf4, 16'h5cf5, 16'h5cf6, 16'h5cf7 	:	val_out <= 16'he10d;
         16'h5cf8, 16'h5cf9, 16'h5cfa, 16'h5cfb, 16'h5cfc, 16'h5cfd, 16'h5cfe, 16'h5cff 	:	val_out <= 16'he0fc;
         16'h5d00, 16'h5d01, 16'h5d02, 16'h5d03, 16'h5d04, 16'h5d05, 16'h5d06, 16'h5d07 	:	val_out <= 16'he0ec;
         16'h5d08, 16'h5d09, 16'h5d0a, 16'h5d0b, 16'h5d0c, 16'h5d0d, 16'h5d0e, 16'h5d0f 	:	val_out <= 16'he0db;
         16'h5d10, 16'h5d11, 16'h5d12, 16'h5d13, 16'h5d14, 16'h5d15, 16'h5d16, 16'h5d17 	:	val_out <= 16'he0cb;
         16'h5d18, 16'h5d19, 16'h5d1a, 16'h5d1b, 16'h5d1c, 16'h5d1d, 16'h5d1e, 16'h5d1f 	:	val_out <= 16'he0ba;
         16'h5d20, 16'h5d21, 16'h5d22, 16'h5d23, 16'h5d24, 16'h5d25, 16'h5d26, 16'h5d27 	:	val_out <= 16'he0aa;
         16'h5d28, 16'h5d29, 16'h5d2a, 16'h5d2b, 16'h5d2c, 16'h5d2d, 16'h5d2e, 16'h5d2f 	:	val_out <= 16'he099;
         16'h5d30, 16'h5d31, 16'h5d32, 16'h5d33, 16'h5d34, 16'h5d35, 16'h5d36, 16'h5d37 	:	val_out <= 16'he089;
         16'h5d38, 16'h5d39, 16'h5d3a, 16'h5d3b, 16'h5d3c, 16'h5d3d, 16'h5d3e, 16'h5d3f 	:	val_out <= 16'he078;
         16'h5d40, 16'h5d41, 16'h5d42, 16'h5d43, 16'h5d44, 16'h5d45, 16'h5d46, 16'h5d47 	:	val_out <= 16'he068;
         16'h5d48, 16'h5d49, 16'h5d4a, 16'h5d4b, 16'h5d4c, 16'h5d4d, 16'h5d4e, 16'h5d4f 	:	val_out <= 16'he057;
         16'h5d50, 16'h5d51, 16'h5d52, 16'h5d53, 16'h5d54, 16'h5d55, 16'h5d56, 16'h5d57 	:	val_out <= 16'he047;
         16'h5d58, 16'h5d59, 16'h5d5a, 16'h5d5b, 16'h5d5c, 16'h5d5d, 16'h5d5e, 16'h5d5f 	:	val_out <= 16'he036;
         16'h5d60, 16'h5d61, 16'h5d62, 16'h5d63, 16'h5d64, 16'h5d65, 16'h5d66, 16'h5d67 	:	val_out <= 16'he026;
         16'h5d68, 16'h5d69, 16'h5d6a, 16'h5d6b, 16'h5d6c, 16'h5d6d, 16'h5d6e, 16'h5d6f 	:	val_out <= 16'he015;
         16'h5d70, 16'h5d71, 16'h5d72, 16'h5d73, 16'h5d74, 16'h5d75, 16'h5d76, 16'h5d77 	:	val_out <= 16'he004;
         16'h5d78, 16'h5d79, 16'h5d7a, 16'h5d7b, 16'h5d7c, 16'h5d7d, 16'h5d7e, 16'h5d7f 	:	val_out <= 16'hdff4;
         16'h5d80, 16'h5d81, 16'h5d82, 16'h5d83, 16'h5d84, 16'h5d85, 16'h5d86, 16'h5d87 	:	val_out <= 16'hdfe3;
         16'h5d88, 16'h5d89, 16'h5d8a, 16'h5d8b, 16'h5d8c, 16'h5d8d, 16'h5d8e, 16'h5d8f 	:	val_out <= 16'hdfd3;
         16'h5d90, 16'h5d91, 16'h5d92, 16'h5d93, 16'h5d94, 16'h5d95, 16'h5d96, 16'h5d97 	:	val_out <= 16'hdfc2;
         16'h5d98, 16'h5d99, 16'h5d9a, 16'h5d9b, 16'h5d9c, 16'h5d9d, 16'h5d9e, 16'h5d9f 	:	val_out <= 16'hdfb1;
         16'h5da0, 16'h5da1, 16'h5da2, 16'h5da3, 16'h5da4, 16'h5da5, 16'h5da6, 16'h5da7 	:	val_out <= 16'hdfa0;
         16'h5da8, 16'h5da9, 16'h5daa, 16'h5dab, 16'h5dac, 16'h5dad, 16'h5dae, 16'h5daf 	:	val_out <= 16'hdf90;
         16'h5db0, 16'h5db1, 16'h5db2, 16'h5db3, 16'h5db4, 16'h5db5, 16'h5db6, 16'h5db7 	:	val_out <= 16'hdf7f;
         16'h5db8, 16'h5db9, 16'h5dba, 16'h5dbb, 16'h5dbc, 16'h5dbd, 16'h5dbe, 16'h5dbf 	:	val_out <= 16'hdf6e;
         16'h5dc0, 16'h5dc1, 16'h5dc2, 16'h5dc3, 16'h5dc4, 16'h5dc5, 16'h5dc6, 16'h5dc7 	:	val_out <= 16'hdf5e;
         16'h5dc8, 16'h5dc9, 16'h5dca, 16'h5dcb, 16'h5dcc, 16'h5dcd, 16'h5dce, 16'h5dcf 	:	val_out <= 16'hdf4d;
         16'h5dd0, 16'h5dd1, 16'h5dd2, 16'h5dd3, 16'h5dd4, 16'h5dd5, 16'h5dd6, 16'h5dd7 	:	val_out <= 16'hdf3c;
         16'h5dd8, 16'h5dd9, 16'h5dda, 16'h5ddb, 16'h5ddc, 16'h5ddd, 16'h5dde, 16'h5ddf 	:	val_out <= 16'hdf2b;
         16'h5de0, 16'h5de1, 16'h5de2, 16'h5de3, 16'h5de4, 16'h5de5, 16'h5de6, 16'h5de7 	:	val_out <= 16'hdf1a;
         16'h5de8, 16'h5de9, 16'h5dea, 16'h5deb, 16'h5dec, 16'h5ded, 16'h5dee, 16'h5def 	:	val_out <= 16'hdf0a;
         16'h5df0, 16'h5df1, 16'h5df2, 16'h5df3, 16'h5df4, 16'h5df5, 16'h5df6, 16'h5df7 	:	val_out <= 16'hdef9;
         16'h5df8, 16'h5df9, 16'h5dfa, 16'h5dfb, 16'h5dfc, 16'h5dfd, 16'h5dfe, 16'h5dff 	:	val_out <= 16'hdee8;
         16'h5e00, 16'h5e01, 16'h5e02, 16'h5e03, 16'h5e04, 16'h5e05, 16'h5e06, 16'h5e07 	:	val_out <= 16'hded7;
         16'h5e08, 16'h5e09, 16'h5e0a, 16'h5e0b, 16'h5e0c, 16'h5e0d, 16'h5e0e, 16'h5e0f 	:	val_out <= 16'hdec6;
         16'h5e10, 16'h5e11, 16'h5e12, 16'h5e13, 16'h5e14, 16'h5e15, 16'h5e16, 16'h5e17 	:	val_out <= 16'hdeb5;
         16'h5e18, 16'h5e19, 16'h5e1a, 16'h5e1b, 16'h5e1c, 16'h5e1d, 16'h5e1e, 16'h5e1f 	:	val_out <= 16'hdea4;
         16'h5e20, 16'h5e21, 16'h5e22, 16'h5e23, 16'h5e24, 16'h5e25, 16'h5e26, 16'h5e27 	:	val_out <= 16'hde93;
         16'h5e28, 16'h5e29, 16'h5e2a, 16'h5e2b, 16'h5e2c, 16'h5e2d, 16'h5e2e, 16'h5e2f 	:	val_out <= 16'hde82;
         16'h5e30, 16'h5e31, 16'h5e32, 16'h5e33, 16'h5e34, 16'h5e35, 16'h5e36, 16'h5e37 	:	val_out <= 16'hde71;
         16'h5e38, 16'h5e39, 16'h5e3a, 16'h5e3b, 16'h5e3c, 16'h5e3d, 16'h5e3e, 16'h5e3f 	:	val_out <= 16'hde60;
         16'h5e40, 16'h5e41, 16'h5e42, 16'h5e43, 16'h5e44, 16'h5e45, 16'h5e46, 16'h5e47 	:	val_out <= 16'hde50;
         16'h5e48, 16'h5e49, 16'h5e4a, 16'h5e4b, 16'h5e4c, 16'h5e4d, 16'h5e4e, 16'h5e4f 	:	val_out <= 16'hde3f;
         16'h5e50, 16'h5e51, 16'h5e52, 16'h5e53, 16'h5e54, 16'h5e55, 16'h5e56, 16'h5e57 	:	val_out <= 16'hde2d;
         16'h5e58, 16'h5e59, 16'h5e5a, 16'h5e5b, 16'h5e5c, 16'h5e5d, 16'h5e5e, 16'h5e5f 	:	val_out <= 16'hde1c;
         16'h5e60, 16'h5e61, 16'h5e62, 16'h5e63, 16'h5e64, 16'h5e65, 16'h5e66, 16'h5e67 	:	val_out <= 16'hde0b;
         16'h5e68, 16'h5e69, 16'h5e6a, 16'h5e6b, 16'h5e6c, 16'h5e6d, 16'h5e6e, 16'h5e6f 	:	val_out <= 16'hddfa;
         16'h5e70, 16'h5e71, 16'h5e72, 16'h5e73, 16'h5e74, 16'h5e75, 16'h5e76, 16'h5e77 	:	val_out <= 16'hdde9;
         16'h5e78, 16'h5e79, 16'h5e7a, 16'h5e7b, 16'h5e7c, 16'h5e7d, 16'h5e7e, 16'h5e7f 	:	val_out <= 16'hddd8;
         16'h5e80, 16'h5e81, 16'h5e82, 16'h5e83, 16'h5e84, 16'h5e85, 16'h5e86, 16'h5e87 	:	val_out <= 16'hddc7;
         16'h5e88, 16'h5e89, 16'h5e8a, 16'h5e8b, 16'h5e8c, 16'h5e8d, 16'h5e8e, 16'h5e8f 	:	val_out <= 16'hddb6;
         16'h5e90, 16'h5e91, 16'h5e92, 16'h5e93, 16'h5e94, 16'h5e95, 16'h5e96, 16'h5e97 	:	val_out <= 16'hdda5;
         16'h5e98, 16'h5e99, 16'h5e9a, 16'h5e9b, 16'h5e9c, 16'h5e9d, 16'h5e9e, 16'h5e9f 	:	val_out <= 16'hdd94;
         16'h5ea0, 16'h5ea1, 16'h5ea2, 16'h5ea3, 16'h5ea4, 16'h5ea5, 16'h5ea6, 16'h5ea7 	:	val_out <= 16'hdd83;
         16'h5ea8, 16'h5ea9, 16'h5eaa, 16'h5eab, 16'h5eac, 16'h5ead, 16'h5eae, 16'h5eaf 	:	val_out <= 16'hdd71;
         16'h5eb0, 16'h5eb1, 16'h5eb2, 16'h5eb3, 16'h5eb4, 16'h5eb5, 16'h5eb6, 16'h5eb7 	:	val_out <= 16'hdd60;
         16'h5eb8, 16'h5eb9, 16'h5eba, 16'h5ebb, 16'h5ebc, 16'h5ebd, 16'h5ebe, 16'h5ebf 	:	val_out <= 16'hdd4f;
         16'h5ec0, 16'h5ec1, 16'h5ec2, 16'h5ec3, 16'h5ec4, 16'h5ec5, 16'h5ec6, 16'h5ec7 	:	val_out <= 16'hdd3e;
         16'h5ec8, 16'h5ec9, 16'h5eca, 16'h5ecb, 16'h5ecc, 16'h5ecd, 16'h5ece, 16'h5ecf 	:	val_out <= 16'hdd2d;
         16'h5ed0, 16'h5ed1, 16'h5ed2, 16'h5ed3, 16'h5ed4, 16'h5ed5, 16'h5ed6, 16'h5ed7 	:	val_out <= 16'hdd1b;
         16'h5ed8, 16'h5ed9, 16'h5eda, 16'h5edb, 16'h5edc, 16'h5edd, 16'h5ede, 16'h5edf 	:	val_out <= 16'hdd0a;
         16'h5ee0, 16'h5ee1, 16'h5ee2, 16'h5ee3, 16'h5ee4, 16'h5ee5, 16'h5ee6, 16'h5ee7 	:	val_out <= 16'hdcf9;
         16'h5ee8, 16'h5ee9, 16'h5eea, 16'h5eeb, 16'h5eec, 16'h5eed, 16'h5eee, 16'h5eef 	:	val_out <= 16'hdce8;
         16'h5ef0, 16'h5ef1, 16'h5ef2, 16'h5ef3, 16'h5ef4, 16'h5ef5, 16'h5ef6, 16'h5ef7 	:	val_out <= 16'hdcd6;
         16'h5ef8, 16'h5ef9, 16'h5efa, 16'h5efb, 16'h5efc, 16'h5efd, 16'h5efe, 16'h5eff 	:	val_out <= 16'hdcc5;
         16'h5f00, 16'h5f01, 16'h5f02, 16'h5f03, 16'h5f04, 16'h5f05, 16'h5f06, 16'h5f07 	:	val_out <= 16'hdcb4;
         16'h5f08, 16'h5f09, 16'h5f0a, 16'h5f0b, 16'h5f0c, 16'h5f0d, 16'h5f0e, 16'h5f0f 	:	val_out <= 16'hdca2;
         16'h5f10, 16'h5f11, 16'h5f12, 16'h5f13, 16'h5f14, 16'h5f15, 16'h5f16, 16'h5f17 	:	val_out <= 16'hdc91;
         16'h5f18, 16'h5f19, 16'h5f1a, 16'h5f1b, 16'h5f1c, 16'h5f1d, 16'h5f1e, 16'h5f1f 	:	val_out <= 16'hdc80;
         16'h5f20, 16'h5f21, 16'h5f22, 16'h5f23, 16'h5f24, 16'h5f25, 16'h5f26, 16'h5f27 	:	val_out <= 16'hdc6e;
         16'h5f28, 16'h5f29, 16'h5f2a, 16'h5f2b, 16'h5f2c, 16'h5f2d, 16'h5f2e, 16'h5f2f 	:	val_out <= 16'hdc5d;
         16'h5f30, 16'h5f31, 16'h5f32, 16'h5f33, 16'h5f34, 16'h5f35, 16'h5f36, 16'h5f37 	:	val_out <= 16'hdc4b;
         16'h5f38, 16'h5f39, 16'h5f3a, 16'h5f3b, 16'h5f3c, 16'h5f3d, 16'h5f3e, 16'h5f3f 	:	val_out <= 16'hdc3a;
         16'h5f40, 16'h5f41, 16'h5f42, 16'h5f43, 16'h5f44, 16'h5f45, 16'h5f46, 16'h5f47 	:	val_out <= 16'hdc29;
         16'h5f48, 16'h5f49, 16'h5f4a, 16'h5f4b, 16'h5f4c, 16'h5f4d, 16'h5f4e, 16'h5f4f 	:	val_out <= 16'hdc17;
         16'h5f50, 16'h5f51, 16'h5f52, 16'h5f53, 16'h5f54, 16'h5f55, 16'h5f56, 16'h5f57 	:	val_out <= 16'hdc06;
         16'h5f58, 16'h5f59, 16'h5f5a, 16'h5f5b, 16'h5f5c, 16'h5f5d, 16'h5f5e, 16'h5f5f 	:	val_out <= 16'hdbf4;
         16'h5f60, 16'h5f61, 16'h5f62, 16'h5f63, 16'h5f64, 16'h5f65, 16'h5f66, 16'h5f67 	:	val_out <= 16'hdbe3;
         16'h5f68, 16'h5f69, 16'h5f6a, 16'h5f6b, 16'h5f6c, 16'h5f6d, 16'h5f6e, 16'h5f6f 	:	val_out <= 16'hdbd1;
         16'h5f70, 16'h5f71, 16'h5f72, 16'h5f73, 16'h5f74, 16'h5f75, 16'h5f76, 16'h5f77 	:	val_out <= 16'hdbc0;
         16'h5f78, 16'h5f79, 16'h5f7a, 16'h5f7b, 16'h5f7c, 16'h5f7d, 16'h5f7e, 16'h5f7f 	:	val_out <= 16'hdbae;
         16'h5f80, 16'h5f81, 16'h5f82, 16'h5f83, 16'h5f84, 16'h5f85, 16'h5f86, 16'h5f87 	:	val_out <= 16'hdb9d;
         16'h5f88, 16'h5f89, 16'h5f8a, 16'h5f8b, 16'h5f8c, 16'h5f8d, 16'h5f8e, 16'h5f8f 	:	val_out <= 16'hdb8b;
         16'h5f90, 16'h5f91, 16'h5f92, 16'h5f93, 16'h5f94, 16'h5f95, 16'h5f96, 16'h5f97 	:	val_out <= 16'hdb79;
         16'h5f98, 16'h5f99, 16'h5f9a, 16'h5f9b, 16'h5f9c, 16'h5f9d, 16'h5f9e, 16'h5f9f 	:	val_out <= 16'hdb68;
         16'h5fa0, 16'h5fa1, 16'h5fa2, 16'h5fa3, 16'h5fa4, 16'h5fa5, 16'h5fa6, 16'h5fa7 	:	val_out <= 16'hdb56;
         16'h5fa8, 16'h5fa9, 16'h5faa, 16'h5fab, 16'h5fac, 16'h5fad, 16'h5fae, 16'h5faf 	:	val_out <= 16'hdb45;
         16'h5fb0, 16'h5fb1, 16'h5fb2, 16'h5fb3, 16'h5fb4, 16'h5fb5, 16'h5fb6, 16'h5fb7 	:	val_out <= 16'hdb33;
         16'h5fb8, 16'h5fb9, 16'h5fba, 16'h5fbb, 16'h5fbc, 16'h5fbd, 16'h5fbe, 16'h5fbf 	:	val_out <= 16'hdb21;
         16'h5fc0, 16'h5fc1, 16'h5fc2, 16'h5fc3, 16'h5fc4, 16'h5fc5, 16'h5fc6, 16'h5fc7 	:	val_out <= 16'hdb10;
         16'h5fc8, 16'h5fc9, 16'h5fca, 16'h5fcb, 16'h5fcc, 16'h5fcd, 16'h5fce, 16'h5fcf 	:	val_out <= 16'hdafe;
         16'h5fd0, 16'h5fd1, 16'h5fd2, 16'h5fd3, 16'h5fd4, 16'h5fd5, 16'h5fd6, 16'h5fd7 	:	val_out <= 16'hdaec;
         16'h5fd8, 16'h5fd9, 16'h5fda, 16'h5fdb, 16'h5fdc, 16'h5fdd, 16'h5fde, 16'h5fdf 	:	val_out <= 16'hdadb;
         16'h5fe0, 16'h5fe1, 16'h5fe2, 16'h5fe3, 16'h5fe4, 16'h5fe5, 16'h5fe6, 16'h5fe7 	:	val_out <= 16'hdac9;
         16'h5fe8, 16'h5fe9, 16'h5fea, 16'h5feb, 16'h5fec, 16'h5fed, 16'h5fee, 16'h5fef 	:	val_out <= 16'hdab7;
         16'h5ff0, 16'h5ff1, 16'h5ff2, 16'h5ff3, 16'h5ff4, 16'h5ff5, 16'h5ff6, 16'h5ff7 	:	val_out <= 16'hdaa5;
         16'h5ff8, 16'h5ff9, 16'h5ffa, 16'h5ffb, 16'h5ffc, 16'h5ffd, 16'h5ffe, 16'h5fff 	:	val_out <= 16'hda94;
         16'h6000, 16'h6001, 16'h6002, 16'h6003, 16'h6004, 16'h6005, 16'h6006, 16'h6007 	:	val_out <= 16'hda82;
         16'h6008, 16'h6009, 16'h600a, 16'h600b, 16'h600c, 16'h600d, 16'h600e, 16'h600f 	:	val_out <= 16'hda70;
         16'h6010, 16'h6011, 16'h6012, 16'h6013, 16'h6014, 16'h6015, 16'h6016, 16'h6017 	:	val_out <= 16'hda5e;
         16'h6018, 16'h6019, 16'h601a, 16'h601b, 16'h601c, 16'h601d, 16'h601e, 16'h601f 	:	val_out <= 16'hda4d;
         16'h6020, 16'h6021, 16'h6022, 16'h6023, 16'h6024, 16'h6025, 16'h6026, 16'h6027 	:	val_out <= 16'hda3b;
         16'h6028, 16'h6029, 16'h602a, 16'h602b, 16'h602c, 16'h602d, 16'h602e, 16'h602f 	:	val_out <= 16'hda29;
         16'h6030, 16'h6031, 16'h6032, 16'h6033, 16'h6034, 16'h6035, 16'h6036, 16'h6037 	:	val_out <= 16'hda17;
         16'h6038, 16'h6039, 16'h603a, 16'h603b, 16'h603c, 16'h603d, 16'h603e, 16'h603f 	:	val_out <= 16'hda05;
         16'h6040, 16'h6041, 16'h6042, 16'h6043, 16'h6044, 16'h6045, 16'h6046, 16'h6047 	:	val_out <= 16'hd9f3;
         16'h6048, 16'h6049, 16'h604a, 16'h604b, 16'h604c, 16'h604d, 16'h604e, 16'h604f 	:	val_out <= 16'hd9e1;
         16'h6050, 16'h6051, 16'h6052, 16'h6053, 16'h6054, 16'h6055, 16'h6056, 16'h6057 	:	val_out <= 16'hd9d0;
         16'h6058, 16'h6059, 16'h605a, 16'h605b, 16'h605c, 16'h605d, 16'h605e, 16'h605f 	:	val_out <= 16'hd9be;
         16'h6060, 16'h6061, 16'h6062, 16'h6063, 16'h6064, 16'h6065, 16'h6066, 16'h6067 	:	val_out <= 16'hd9ac;
         16'h6068, 16'h6069, 16'h606a, 16'h606b, 16'h606c, 16'h606d, 16'h606e, 16'h606f 	:	val_out <= 16'hd99a;
         16'h6070, 16'h6071, 16'h6072, 16'h6073, 16'h6074, 16'h6075, 16'h6076, 16'h6077 	:	val_out <= 16'hd988;
         16'h6078, 16'h6079, 16'h607a, 16'h607b, 16'h607c, 16'h607d, 16'h607e, 16'h607f 	:	val_out <= 16'hd976;
         16'h6080, 16'h6081, 16'h6082, 16'h6083, 16'h6084, 16'h6085, 16'h6086, 16'h6087 	:	val_out <= 16'hd964;
         16'h6088, 16'h6089, 16'h608a, 16'h608b, 16'h608c, 16'h608d, 16'h608e, 16'h608f 	:	val_out <= 16'hd952;
         16'h6090, 16'h6091, 16'h6092, 16'h6093, 16'h6094, 16'h6095, 16'h6096, 16'h6097 	:	val_out <= 16'hd940;
         16'h6098, 16'h6099, 16'h609a, 16'h609b, 16'h609c, 16'h609d, 16'h609e, 16'h609f 	:	val_out <= 16'hd92e;
         16'h60a0, 16'h60a1, 16'h60a2, 16'h60a3, 16'h60a4, 16'h60a5, 16'h60a6, 16'h60a7 	:	val_out <= 16'hd91c;
         16'h60a8, 16'h60a9, 16'h60aa, 16'h60ab, 16'h60ac, 16'h60ad, 16'h60ae, 16'h60af 	:	val_out <= 16'hd90a;
         16'h60b0, 16'h60b1, 16'h60b2, 16'h60b3, 16'h60b4, 16'h60b5, 16'h60b6, 16'h60b7 	:	val_out <= 16'hd8f8;
         16'h60b8, 16'h60b9, 16'h60ba, 16'h60bb, 16'h60bc, 16'h60bd, 16'h60be, 16'h60bf 	:	val_out <= 16'hd8e6;
         16'h60c0, 16'h60c1, 16'h60c2, 16'h60c3, 16'h60c4, 16'h60c5, 16'h60c6, 16'h60c7 	:	val_out <= 16'hd8d4;
         16'h60c8, 16'h60c9, 16'h60ca, 16'h60cb, 16'h60cc, 16'h60cd, 16'h60ce, 16'h60cf 	:	val_out <= 16'hd8c1;
         16'h60d0, 16'h60d1, 16'h60d2, 16'h60d3, 16'h60d4, 16'h60d5, 16'h60d6, 16'h60d7 	:	val_out <= 16'hd8af;
         16'h60d8, 16'h60d9, 16'h60da, 16'h60db, 16'h60dc, 16'h60dd, 16'h60de, 16'h60df 	:	val_out <= 16'hd89d;
         16'h60e0, 16'h60e1, 16'h60e2, 16'h60e3, 16'h60e4, 16'h60e5, 16'h60e6, 16'h60e7 	:	val_out <= 16'hd88b;
         16'h60e8, 16'h60e9, 16'h60ea, 16'h60eb, 16'h60ec, 16'h60ed, 16'h60ee, 16'h60ef 	:	val_out <= 16'hd879;
         16'h60f0, 16'h60f1, 16'h60f2, 16'h60f3, 16'h60f4, 16'h60f5, 16'h60f6, 16'h60f7 	:	val_out <= 16'hd867;
         16'h60f8, 16'h60f9, 16'h60fa, 16'h60fb, 16'h60fc, 16'h60fd, 16'h60fe, 16'h60ff 	:	val_out <= 16'hd855;
         16'h6100, 16'h6101, 16'h6102, 16'h6103, 16'h6104, 16'h6105, 16'h6106, 16'h6107 	:	val_out <= 16'hd842;
         16'h6108, 16'h6109, 16'h610a, 16'h610b, 16'h610c, 16'h610d, 16'h610e, 16'h610f 	:	val_out <= 16'hd830;
         16'h6110, 16'h6111, 16'h6112, 16'h6113, 16'h6114, 16'h6115, 16'h6116, 16'h6117 	:	val_out <= 16'hd81e;
         16'h6118, 16'h6119, 16'h611a, 16'h611b, 16'h611c, 16'h611d, 16'h611e, 16'h611f 	:	val_out <= 16'hd80c;
         16'h6120, 16'h6121, 16'h6122, 16'h6123, 16'h6124, 16'h6125, 16'h6126, 16'h6127 	:	val_out <= 16'hd7f9;
         16'h6128, 16'h6129, 16'h612a, 16'h612b, 16'h612c, 16'h612d, 16'h612e, 16'h612f 	:	val_out <= 16'hd7e7;
         16'h6130, 16'h6131, 16'h6132, 16'h6133, 16'h6134, 16'h6135, 16'h6136, 16'h6137 	:	val_out <= 16'hd7d5;
         16'h6138, 16'h6139, 16'h613a, 16'h613b, 16'h613c, 16'h613d, 16'h613e, 16'h613f 	:	val_out <= 16'hd7c3;
         16'h6140, 16'h6141, 16'h6142, 16'h6143, 16'h6144, 16'h6145, 16'h6146, 16'h6147 	:	val_out <= 16'hd7b0;
         16'h6148, 16'h6149, 16'h614a, 16'h614b, 16'h614c, 16'h614d, 16'h614e, 16'h614f 	:	val_out <= 16'hd79e;
         16'h6150, 16'h6151, 16'h6152, 16'h6153, 16'h6154, 16'h6155, 16'h6156, 16'h6157 	:	val_out <= 16'hd78c;
         16'h6158, 16'h6159, 16'h615a, 16'h615b, 16'h615c, 16'h615d, 16'h615e, 16'h615f 	:	val_out <= 16'hd779;
         16'h6160, 16'h6161, 16'h6162, 16'h6163, 16'h6164, 16'h6165, 16'h6166, 16'h6167 	:	val_out <= 16'hd767;
         16'h6168, 16'h6169, 16'h616a, 16'h616b, 16'h616c, 16'h616d, 16'h616e, 16'h616f 	:	val_out <= 16'hd755;
         16'h6170, 16'h6171, 16'h6172, 16'h6173, 16'h6174, 16'h6175, 16'h6176, 16'h6177 	:	val_out <= 16'hd742;
         16'h6178, 16'h6179, 16'h617a, 16'h617b, 16'h617c, 16'h617d, 16'h617e, 16'h617f 	:	val_out <= 16'hd730;
         16'h6180, 16'h6181, 16'h6182, 16'h6183, 16'h6184, 16'h6185, 16'h6186, 16'h6187 	:	val_out <= 16'hd71d;
         16'h6188, 16'h6189, 16'h618a, 16'h618b, 16'h618c, 16'h618d, 16'h618e, 16'h618f 	:	val_out <= 16'hd70b;
         16'h6190, 16'h6191, 16'h6192, 16'h6193, 16'h6194, 16'h6195, 16'h6196, 16'h6197 	:	val_out <= 16'hd6f9;
         16'h6198, 16'h6199, 16'h619a, 16'h619b, 16'h619c, 16'h619d, 16'h619e, 16'h619f 	:	val_out <= 16'hd6e6;
         16'h61a0, 16'h61a1, 16'h61a2, 16'h61a3, 16'h61a4, 16'h61a5, 16'h61a6, 16'h61a7 	:	val_out <= 16'hd6d4;
         16'h61a8, 16'h61a9, 16'h61aa, 16'h61ab, 16'h61ac, 16'h61ad, 16'h61ae, 16'h61af 	:	val_out <= 16'hd6c1;
         16'h61b0, 16'h61b1, 16'h61b2, 16'h61b3, 16'h61b4, 16'h61b5, 16'h61b6, 16'h61b7 	:	val_out <= 16'hd6af;
         16'h61b8, 16'h61b9, 16'h61ba, 16'h61bb, 16'h61bc, 16'h61bd, 16'h61be, 16'h61bf 	:	val_out <= 16'hd69c;
         16'h61c0, 16'h61c1, 16'h61c2, 16'h61c3, 16'h61c4, 16'h61c5, 16'h61c6, 16'h61c7 	:	val_out <= 16'hd68a;
         16'h61c8, 16'h61c9, 16'h61ca, 16'h61cb, 16'h61cc, 16'h61cd, 16'h61ce, 16'h61cf 	:	val_out <= 16'hd677;
         16'h61d0, 16'h61d1, 16'h61d2, 16'h61d3, 16'h61d4, 16'h61d5, 16'h61d6, 16'h61d7 	:	val_out <= 16'hd665;
         16'h61d8, 16'h61d9, 16'h61da, 16'h61db, 16'h61dc, 16'h61dd, 16'h61de, 16'h61df 	:	val_out <= 16'hd652;
         16'h61e0, 16'h61e1, 16'h61e2, 16'h61e3, 16'h61e4, 16'h61e5, 16'h61e6, 16'h61e7 	:	val_out <= 16'hd640;
         16'h61e8, 16'h61e9, 16'h61ea, 16'h61eb, 16'h61ec, 16'h61ed, 16'h61ee, 16'h61ef 	:	val_out <= 16'hd62d;
         16'h61f0, 16'h61f1, 16'h61f2, 16'h61f3, 16'h61f4, 16'h61f5, 16'h61f6, 16'h61f7 	:	val_out <= 16'hd61a;
         16'h61f8, 16'h61f9, 16'h61fa, 16'h61fb, 16'h61fc, 16'h61fd, 16'h61fe, 16'h61ff 	:	val_out <= 16'hd608;
         16'h6200, 16'h6201, 16'h6202, 16'h6203, 16'h6204, 16'h6205, 16'h6206, 16'h6207 	:	val_out <= 16'hd5f5;
         16'h6208, 16'h6209, 16'h620a, 16'h620b, 16'h620c, 16'h620d, 16'h620e, 16'h620f 	:	val_out <= 16'hd5e3;
         16'h6210, 16'h6211, 16'h6212, 16'h6213, 16'h6214, 16'h6215, 16'h6216, 16'h6217 	:	val_out <= 16'hd5d0;
         16'h6218, 16'h6219, 16'h621a, 16'h621b, 16'h621c, 16'h621d, 16'h621e, 16'h621f 	:	val_out <= 16'hd5bd;
         16'h6220, 16'h6221, 16'h6222, 16'h6223, 16'h6224, 16'h6225, 16'h6226, 16'h6227 	:	val_out <= 16'hd5ab;
         16'h6228, 16'h6229, 16'h622a, 16'h622b, 16'h622c, 16'h622d, 16'h622e, 16'h622f 	:	val_out <= 16'hd598;
         16'h6230, 16'h6231, 16'h6232, 16'h6233, 16'h6234, 16'h6235, 16'h6236, 16'h6237 	:	val_out <= 16'hd585;
         16'h6238, 16'h6239, 16'h623a, 16'h623b, 16'h623c, 16'h623d, 16'h623e, 16'h623f 	:	val_out <= 16'hd572;
         16'h6240, 16'h6241, 16'h6242, 16'h6243, 16'h6244, 16'h6245, 16'h6246, 16'h6247 	:	val_out <= 16'hd560;
         16'h6248, 16'h6249, 16'h624a, 16'h624b, 16'h624c, 16'h624d, 16'h624e, 16'h624f 	:	val_out <= 16'hd54d;
         16'h6250, 16'h6251, 16'h6252, 16'h6253, 16'h6254, 16'h6255, 16'h6256, 16'h6257 	:	val_out <= 16'hd53a;
         16'h6258, 16'h6259, 16'h625a, 16'h625b, 16'h625c, 16'h625d, 16'h625e, 16'h625f 	:	val_out <= 16'hd528;
         16'h6260, 16'h6261, 16'h6262, 16'h6263, 16'h6264, 16'h6265, 16'h6266, 16'h6267 	:	val_out <= 16'hd515;
         16'h6268, 16'h6269, 16'h626a, 16'h626b, 16'h626c, 16'h626d, 16'h626e, 16'h626f 	:	val_out <= 16'hd502;
         16'h6270, 16'h6271, 16'h6272, 16'h6273, 16'h6274, 16'h6275, 16'h6276, 16'h6277 	:	val_out <= 16'hd4ef;
         16'h6278, 16'h6279, 16'h627a, 16'h627b, 16'h627c, 16'h627d, 16'h627e, 16'h627f 	:	val_out <= 16'hd4dc;
         16'h6280, 16'h6281, 16'h6282, 16'h6283, 16'h6284, 16'h6285, 16'h6286, 16'h6287 	:	val_out <= 16'hd4ca;
         16'h6288, 16'h6289, 16'h628a, 16'h628b, 16'h628c, 16'h628d, 16'h628e, 16'h628f 	:	val_out <= 16'hd4b7;
         16'h6290, 16'h6291, 16'h6292, 16'h6293, 16'h6294, 16'h6295, 16'h6296, 16'h6297 	:	val_out <= 16'hd4a4;
         16'h6298, 16'h6299, 16'h629a, 16'h629b, 16'h629c, 16'h629d, 16'h629e, 16'h629f 	:	val_out <= 16'hd491;
         16'h62a0, 16'h62a1, 16'h62a2, 16'h62a3, 16'h62a4, 16'h62a5, 16'h62a6, 16'h62a7 	:	val_out <= 16'hd47e;
         16'h62a8, 16'h62a9, 16'h62aa, 16'h62ab, 16'h62ac, 16'h62ad, 16'h62ae, 16'h62af 	:	val_out <= 16'hd46b;
         16'h62b0, 16'h62b1, 16'h62b2, 16'h62b3, 16'h62b4, 16'h62b5, 16'h62b6, 16'h62b7 	:	val_out <= 16'hd458;
         16'h62b8, 16'h62b9, 16'h62ba, 16'h62bb, 16'h62bc, 16'h62bd, 16'h62be, 16'h62bf 	:	val_out <= 16'hd445;
         16'h62c0, 16'h62c1, 16'h62c2, 16'h62c3, 16'h62c4, 16'h62c5, 16'h62c6, 16'h62c7 	:	val_out <= 16'hd433;
         16'h62c8, 16'h62c9, 16'h62ca, 16'h62cb, 16'h62cc, 16'h62cd, 16'h62ce, 16'h62cf 	:	val_out <= 16'hd420;
         16'h62d0, 16'h62d1, 16'h62d2, 16'h62d3, 16'h62d4, 16'h62d5, 16'h62d6, 16'h62d7 	:	val_out <= 16'hd40d;
         16'h62d8, 16'h62d9, 16'h62da, 16'h62db, 16'h62dc, 16'h62dd, 16'h62de, 16'h62df 	:	val_out <= 16'hd3fa;
         16'h62e0, 16'h62e1, 16'h62e2, 16'h62e3, 16'h62e4, 16'h62e5, 16'h62e6, 16'h62e7 	:	val_out <= 16'hd3e7;
         16'h62e8, 16'h62e9, 16'h62ea, 16'h62eb, 16'h62ec, 16'h62ed, 16'h62ee, 16'h62ef 	:	val_out <= 16'hd3d4;
         16'h62f0, 16'h62f1, 16'h62f2, 16'h62f3, 16'h62f4, 16'h62f5, 16'h62f6, 16'h62f7 	:	val_out <= 16'hd3c1;
         16'h62f8, 16'h62f9, 16'h62fa, 16'h62fb, 16'h62fc, 16'h62fd, 16'h62fe, 16'h62ff 	:	val_out <= 16'hd3ae;
         16'h6300, 16'h6301, 16'h6302, 16'h6303, 16'h6304, 16'h6305, 16'h6306, 16'h6307 	:	val_out <= 16'hd39b;
         16'h6308, 16'h6309, 16'h630a, 16'h630b, 16'h630c, 16'h630d, 16'h630e, 16'h630f 	:	val_out <= 16'hd388;
         16'h6310, 16'h6311, 16'h6312, 16'h6313, 16'h6314, 16'h6315, 16'h6316, 16'h6317 	:	val_out <= 16'hd375;
         16'h6318, 16'h6319, 16'h631a, 16'h631b, 16'h631c, 16'h631d, 16'h631e, 16'h631f 	:	val_out <= 16'hd362;
         16'h6320, 16'h6321, 16'h6322, 16'h6323, 16'h6324, 16'h6325, 16'h6326, 16'h6327 	:	val_out <= 16'hd34e;
         16'h6328, 16'h6329, 16'h632a, 16'h632b, 16'h632c, 16'h632d, 16'h632e, 16'h632f 	:	val_out <= 16'hd33b;
         16'h6330, 16'h6331, 16'h6332, 16'h6333, 16'h6334, 16'h6335, 16'h6336, 16'h6337 	:	val_out <= 16'hd328;
         16'h6338, 16'h6339, 16'h633a, 16'h633b, 16'h633c, 16'h633d, 16'h633e, 16'h633f 	:	val_out <= 16'hd315;
         16'h6340, 16'h6341, 16'h6342, 16'h6343, 16'h6344, 16'h6345, 16'h6346, 16'h6347 	:	val_out <= 16'hd302;
         16'h6348, 16'h6349, 16'h634a, 16'h634b, 16'h634c, 16'h634d, 16'h634e, 16'h634f 	:	val_out <= 16'hd2ef;
         16'h6350, 16'h6351, 16'h6352, 16'h6353, 16'h6354, 16'h6355, 16'h6356, 16'h6357 	:	val_out <= 16'hd2dc;
         16'h6358, 16'h6359, 16'h635a, 16'h635b, 16'h635c, 16'h635d, 16'h635e, 16'h635f 	:	val_out <= 16'hd2c9;
         16'h6360, 16'h6361, 16'h6362, 16'h6363, 16'h6364, 16'h6365, 16'h6366, 16'h6367 	:	val_out <= 16'hd2b5;
         16'h6368, 16'h6369, 16'h636a, 16'h636b, 16'h636c, 16'h636d, 16'h636e, 16'h636f 	:	val_out <= 16'hd2a2;
         16'h6370, 16'h6371, 16'h6372, 16'h6373, 16'h6374, 16'h6375, 16'h6376, 16'h6377 	:	val_out <= 16'hd28f;
         16'h6378, 16'h6379, 16'h637a, 16'h637b, 16'h637c, 16'h637d, 16'h637e, 16'h637f 	:	val_out <= 16'hd27c;
         16'h6380, 16'h6381, 16'h6382, 16'h6383, 16'h6384, 16'h6385, 16'h6386, 16'h6387 	:	val_out <= 16'hd269;
         16'h6388, 16'h6389, 16'h638a, 16'h638b, 16'h638c, 16'h638d, 16'h638e, 16'h638f 	:	val_out <= 16'hd255;
         16'h6390, 16'h6391, 16'h6392, 16'h6393, 16'h6394, 16'h6395, 16'h6396, 16'h6397 	:	val_out <= 16'hd242;
         16'h6398, 16'h6399, 16'h639a, 16'h639b, 16'h639c, 16'h639d, 16'h639e, 16'h639f 	:	val_out <= 16'hd22f;
         16'h63a0, 16'h63a1, 16'h63a2, 16'h63a3, 16'h63a4, 16'h63a5, 16'h63a6, 16'h63a7 	:	val_out <= 16'hd21c;
         16'h63a8, 16'h63a9, 16'h63aa, 16'h63ab, 16'h63ac, 16'h63ad, 16'h63ae, 16'h63af 	:	val_out <= 16'hd208;
         16'h63b0, 16'h63b1, 16'h63b2, 16'h63b3, 16'h63b4, 16'h63b5, 16'h63b6, 16'h63b7 	:	val_out <= 16'hd1f5;
         16'h63b8, 16'h63b9, 16'h63ba, 16'h63bb, 16'h63bc, 16'h63bd, 16'h63be, 16'h63bf 	:	val_out <= 16'hd1e2;
         16'h63c0, 16'h63c1, 16'h63c2, 16'h63c3, 16'h63c4, 16'h63c5, 16'h63c6, 16'h63c7 	:	val_out <= 16'hd1ce;
         16'h63c8, 16'h63c9, 16'h63ca, 16'h63cb, 16'h63cc, 16'h63cd, 16'h63ce, 16'h63cf 	:	val_out <= 16'hd1bb;
         16'h63d0, 16'h63d1, 16'h63d2, 16'h63d3, 16'h63d4, 16'h63d5, 16'h63d6, 16'h63d7 	:	val_out <= 16'hd1a8;
         16'h63d8, 16'h63d9, 16'h63da, 16'h63db, 16'h63dc, 16'h63dd, 16'h63de, 16'h63df 	:	val_out <= 16'hd194;
         16'h63e0, 16'h63e1, 16'h63e2, 16'h63e3, 16'h63e4, 16'h63e5, 16'h63e6, 16'h63e7 	:	val_out <= 16'hd181;
         16'h63e8, 16'h63e9, 16'h63ea, 16'h63eb, 16'h63ec, 16'h63ed, 16'h63ee, 16'h63ef 	:	val_out <= 16'hd16e;
         16'h63f0, 16'h63f1, 16'h63f2, 16'h63f3, 16'h63f4, 16'h63f5, 16'h63f6, 16'h63f7 	:	val_out <= 16'hd15a;
         16'h63f8, 16'h63f9, 16'h63fa, 16'h63fb, 16'h63fc, 16'h63fd, 16'h63fe, 16'h63ff 	:	val_out <= 16'hd147;
         16'h6400, 16'h6401, 16'h6402, 16'h6403, 16'h6404, 16'h6405, 16'h6406, 16'h6407 	:	val_out <= 16'hd133;
         16'h6408, 16'h6409, 16'h640a, 16'h640b, 16'h640c, 16'h640d, 16'h640e, 16'h640f 	:	val_out <= 16'hd120;
         16'h6410, 16'h6411, 16'h6412, 16'h6413, 16'h6414, 16'h6415, 16'h6416, 16'h6417 	:	val_out <= 16'hd10c;
         16'h6418, 16'h6419, 16'h641a, 16'h641b, 16'h641c, 16'h641d, 16'h641e, 16'h641f 	:	val_out <= 16'hd0f9;
         16'h6420, 16'h6421, 16'h6422, 16'h6423, 16'h6424, 16'h6425, 16'h6426, 16'h6427 	:	val_out <= 16'hd0e5;
         16'h6428, 16'h6429, 16'h642a, 16'h642b, 16'h642c, 16'h642d, 16'h642e, 16'h642f 	:	val_out <= 16'hd0d2;
         16'h6430, 16'h6431, 16'h6432, 16'h6433, 16'h6434, 16'h6435, 16'h6436, 16'h6437 	:	val_out <= 16'hd0bf;
         16'h6438, 16'h6439, 16'h643a, 16'h643b, 16'h643c, 16'h643d, 16'h643e, 16'h643f 	:	val_out <= 16'hd0ab;
         16'h6440, 16'h6441, 16'h6442, 16'h6443, 16'h6444, 16'h6445, 16'h6446, 16'h6447 	:	val_out <= 16'hd097;
         16'h6448, 16'h6449, 16'h644a, 16'h644b, 16'h644c, 16'h644d, 16'h644e, 16'h644f 	:	val_out <= 16'hd084;
         16'h6450, 16'h6451, 16'h6452, 16'h6453, 16'h6454, 16'h6455, 16'h6456, 16'h6457 	:	val_out <= 16'hd070;
         16'h6458, 16'h6459, 16'h645a, 16'h645b, 16'h645c, 16'h645d, 16'h645e, 16'h645f 	:	val_out <= 16'hd05d;
         16'h6460, 16'h6461, 16'h6462, 16'h6463, 16'h6464, 16'h6465, 16'h6466, 16'h6467 	:	val_out <= 16'hd049;
         16'h6468, 16'h6469, 16'h646a, 16'h646b, 16'h646c, 16'h646d, 16'h646e, 16'h646f 	:	val_out <= 16'hd036;
         16'h6470, 16'h6471, 16'h6472, 16'h6473, 16'h6474, 16'h6475, 16'h6476, 16'h6477 	:	val_out <= 16'hd022;
         16'h6478, 16'h6479, 16'h647a, 16'h647b, 16'h647c, 16'h647d, 16'h647e, 16'h647f 	:	val_out <= 16'hd00f;
         16'h6480, 16'h6481, 16'h6482, 16'h6483, 16'h6484, 16'h6485, 16'h6486, 16'h6487 	:	val_out <= 16'hcffb;
         16'h6488, 16'h6489, 16'h648a, 16'h648b, 16'h648c, 16'h648d, 16'h648e, 16'h648f 	:	val_out <= 16'hcfe7;
         16'h6490, 16'h6491, 16'h6492, 16'h6493, 16'h6494, 16'h6495, 16'h6496, 16'h6497 	:	val_out <= 16'hcfd4;
         16'h6498, 16'h6499, 16'h649a, 16'h649b, 16'h649c, 16'h649d, 16'h649e, 16'h649f 	:	val_out <= 16'hcfc0;
         16'h64a0, 16'h64a1, 16'h64a2, 16'h64a3, 16'h64a4, 16'h64a5, 16'h64a6, 16'h64a7 	:	val_out <= 16'hcfac;
         16'h64a8, 16'h64a9, 16'h64aa, 16'h64ab, 16'h64ac, 16'h64ad, 16'h64ae, 16'h64af 	:	val_out <= 16'hcf99;
         16'h64b0, 16'h64b1, 16'h64b2, 16'h64b3, 16'h64b4, 16'h64b5, 16'h64b6, 16'h64b7 	:	val_out <= 16'hcf85;
         16'h64b8, 16'h64b9, 16'h64ba, 16'h64bb, 16'h64bc, 16'h64bd, 16'h64be, 16'h64bf 	:	val_out <= 16'hcf71;
         16'h64c0, 16'h64c1, 16'h64c2, 16'h64c3, 16'h64c4, 16'h64c5, 16'h64c6, 16'h64c7 	:	val_out <= 16'hcf5e;
         16'h64c8, 16'h64c9, 16'h64ca, 16'h64cb, 16'h64cc, 16'h64cd, 16'h64ce, 16'h64cf 	:	val_out <= 16'hcf4a;
         16'h64d0, 16'h64d1, 16'h64d2, 16'h64d3, 16'h64d4, 16'h64d5, 16'h64d6, 16'h64d7 	:	val_out <= 16'hcf36;
         16'h64d8, 16'h64d9, 16'h64da, 16'h64db, 16'h64dc, 16'h64dd, 16'h64de, 16'h64df 	:	val_out <= 16'hcf22;
         16'h64e0, 16'h64e1, 16'h64e2, 16'h64e3, 16'h64e4, 16'h64e5, 16'h64e6, 16'h64e7 	:	val_out <= 16'hcf0f;
         16'h64e8, 16'h64e9, 16'h64ea, 16'h64eb, 16'h64ec, 16'h64ed, 16'h64ee, 16'h64ef 	:	val_out <= 16'hcefb;
         16'h64f0, 16'h64f1, 16'h64f2, 16'h64f3, 16'h64f4, 16'h64f5, 16'h64f6, 16'h64f7 	:	val_out <= 16'hcee7;
         16'h64f8, 16'h64f9, 16'h64fa, 16'h64fb, 16'h64fc, 16'h64fd, 16'h64fe, 16'h64ff 	:	val_out <= 16'hced3;
         16'h6500, 16'h6501, 16'h6502, 16'h6503, 16'h6504, 16'h6505, 16'h6506, 16'h6507 	:	val_out <= 16'hcebf;
         16'h6508, 16'h6509, 16'h650a, 16'h650b, 16'h650c, 16'h650d, 16'h650e, 16'h650f 	:	val_out <= 16'hceac;
         16'h6510, 16'h6511, 16'h6512, 16'h6513, 16'h6514, 16'h6515, 16'h6516, 16'h6517 	:	val_out <= 16'hce98;
         16'h6518, 16'h6519, 16'h651a, 16'h651b, 16'h651c, 16'h651d, 16'h651e, 16'h651f 	:	val_out <= 16'hce84;
         16'h6520, 16'h6521, 16'h6522, 16'h6523, 16'h6524, 16'h6525, 16'h6526, 16'h6527 	:	val_out <= 16'hce70;
         16'h6528, 16'h6529, 16'h652a, 16'h652b, 16'h652c, 16'h652d, 16'h652e, 16'h652f 	:	val_out <= 16'hce5c;
         16'h6530, 16'h6531, 16'h6532, 16'h6533, 16'h6534, 16'h6535, 16'h6536, 16'h6537 	:	val_out <= 16'hce48;
         16'h6538, 16'h6539, 16'h653a, 16'h653b, 16'h653c, 16'h653d, 16'h653e, 16'h653f 	:	val_out <= 16'hce34;
         16'h6540, 16'h6541, 16'h6542, 16'h6543, 16'h6544, 16'h6545, 16'h6546, 16'h6547 	:	val_out <= 16'hce21;
         16'h6548, 16'h6549, 16'h654a, 16'h654b, 16'h654c, 16'h654d, 16'h654e, 16'h654f 	:	val_out <= 16'hce0d;
         16'h6550, 16'h6551, 16'h6552, 16'h6553, 16'h6554, 16'h6555, 16'h6556, 16'h6557 	:	val_out <= 16'hcdf9;
         16'h6558, 16'h6559, 16'h655a, 16'h655b, 16'h655c, 16'h655d, 16'h655e, 16'h655f 	:	val_out <= 16'hcde5;
         16'h6560, 16'h6561, 16'h6562, 16'h6563, 16'h6564, 16'h6565, 16'h6566, 16'h6567 	:	val_out <= 16'hcdd1;
         16'h6568, 16'h6569, 16'h656a, 16'h656b, 16'h656c, 16'h656d, 16'h656e, 16'h656f 	:	val_out <= 16'hcdbd;
         16'h6570, 16'h6571, 16'h6572, 16'h6573, 16'h6574, 16'h6575, 16'h6576, 16'h6577 	:	val_out <= 16'hcda9;
         16'h6578, 16'h6579, 16'h657a, 16'h657b, 16'h657c, 16'h657d, 16'h657e, 16'h657f 	:	val_out <= 16'hcd95;
         16'h6580, 16'h6581, 16'h6582, 16'h6583, 16'h6584, 16'h6585, 16'h6586, 16'h6587 	:	val_out <= 16'hcd81;
         16'h6588, 16'h6589, 16'h658a, 16'h658b, 16'h658c, 16'h658d, 16'h658e, 16'h658f 	:	val_out <= 16'hcd6d;
         16'h6590, 16'h6591, 16'h6592, 16'h6593, 16'h6594, 16'h6595, 16'h6596, 16'h6597 	:	val_out <= 16'hcd59;
         16'h6598, 16'h6599, 16'h659a, 16'h659b, 16'h659c, 16'h659d, 16'h659e, 16'h659f 	:	val_out <= 16'hcd45;
         16'h65a0, 16'h65a1, 16'h65a2, 16'h65a3, 16'h65a4, 16'h65a5, 16'h65a6, 16'h65a7 	:	val_out <= 16'hcd31;
         16'h65a8, 16'h65a9, 16'h65aa, 16'h65ab, 16'h65ac, 16'h65ad, 16'h65ae, 16'h65af 	:	val_out <= 16'hcd1d;
         16'h65b0, 16'h65b1, 16'h65b2, 16'h65b3, 16'h65b4, 16'h65b5, 16'h65b6, 16'h65b7 	:	val_out <= 16'hcd09;
         16'h65b8, 16'h65b9, 16'h65ba, 16'h65bb, 16'h65bc, 16'h65bd, 16'h65be, 16'h65bf 	:	val_out <= 16'hccf5;
         16'h65c0, 16'h65c1, 16'h65c2, 16'h65c3, 16'h65c4, 16'h65c5, 16'h65c6, 16'h65c7 	:	val_out <= 16'hcce1;
         16'h65c8, 16'h65c9, 16'h65ca, 16'h65cb, 16'h65cc, 16'h65cd, 16'h65ce, 16'h65cf 	:	val_out <= 16'hcccc;
         16'h65d0, 16'h65d1, 16'h65d2, 16'h65d3, 16'h65d4, 16'h65d5, 16'h65d6, 16'h65d7 	:	val_out <= 16'hccb8;
         16'h65d8, 16'h65d9, 16'h65da, 16'h65db, 16'h65dc, 16'h65dd, 16'h65de, 16'h65df 	:	val_out <= 16'hcca4;
         16'h65e0, 16'h65e1, 16'h65e2, 16'h65e3, 16'h65e4, 16'h65e5, 16'h65e6, 16'h65e7 	:	val_out <= 16'hcc90;
         16'h65e8, 16'h65e9, 16'h65ea, 16'h65eb, 16'h65ec, 16'h65ed, 16'h65ee, 16'h65ef 	:	val_out <= 16'hcc7c;
         16'h65f0, 16'h65f1, 16'h65f2, 16'h65f3, 16'h65f4, 16'h65f5, 16'h65f6, 16'h65f7 	:	val_out <= 16'hcc68;
         16'h65f8, 16'h65f9, 16'h65fa, 16'h65fb, 16'h65fc, 16'h65fd, 16'h65fe, 16'h65ff 	:	val_out <= 16'hcc54;
         16'h6600, 16'h6601, 16'h6602, 16'h6603, 16'h6604, 16'h6605, 16'h6606, 16'h6607 	:	val_out <= 16'hcc3f;
         16'h6608, 16'h6609, 16'h660a, 16'h660b, 16'h660c, 16'h660d, 16'h660e, 16'h660f 	:	val_out <= 16'hcc2b;
         16'h6610, 16'h6611, 16'h6612, 16'h6613, 16'h6614, 16'h6615, 16'h6616, 16'h6617 	:	val_out <= 16'hcc17;
         16'h6618, 16'h6619, 16'h661a, 16'h661b, 16'h661c, 16'h661d, 16'h661e, 16'h661f 	:	val_out <= 16'hcc03;
         16'h6620, 16'h6621, 16'h6622, 16'h6623, 16'h6624, 16'h6625, 16'h6626, 16'h6627 	:	val_out <= 16'hcbef;
         16'h6628, 16'h6629, 16'h662a, 16'h662b, 16'h662c, 16'h662d, 16'h662e, 16'h662f 	:	val_out <= 16'hcbda;
         16'h6630, 16'h6631, 16'h6632, 16'h6633, 16'h6634, 16'h6635, 16'h6636, 16'h6637 	:	val_out <= 16'hcbc6;
         16'h6638, 16'h6639, 16'h663a, 16'h663b, 16'h663c, 16'h663d, 16'h663e, 16'h663f 	:	val_out <= 16'hcbb2;
         16'h6640, 16'h6641, 16'h6642, 16'h6643, 16'h6644, 16'h6645, 16'h6646, 16'h6647 	:	val_out <= 16'hcb9e;
         16'h6648, 16'h6649, 16'h664a, 16'h664b, 16'h664c, 16'h664d, 16'h664e, 16'h664f 	:	val_out <= 16'hcb89;
         16'h6650, 16'h6651, 16'h6652, 16'h6653, 16'h6654, 16'h6655, 16'h6656, 16'h6657 	:	val_out <= 16'hcb75;
         16'h6658, 16'h6659, 16'h665a, 16'h665b, 16'h665c, 16'h665d, 16'h665e, 16'h665f 	:	val_out <= 16'hcb61;
         16'h6660, 16'h6661, 16'h6662, 16'h6663, 16'h6664, 16'h6665, 16'h6666, 16'h6667 	:	val_out <= 16'hcb4c;
         16'h6668, 16'h6669, 16'h666a, 16'h666b, 16'h666c, 16'h666d, 16'h666e, 16'h666f 	:	val_out <= 16'hcb38;
         16'h6670, 16'h6671, 16'h6672, 16'h6673, 16'h6674, 16'h6675, 16'h6676, 16'h6677 	:	val_out <= 16'hcb24;
         16'h6678, 16'h6679, 16'h667a, 16'h667b, 16'h667c, 16'h667d, 16'h667e, 16'h667f 	:	val_out <= 16'hcb0f;
         16'h6680, 16'h6681, 16'h6682, 16'h6683, 16'h6684, 16'h6685, 16'h6686, 16'h6687 	:	val_out <= 16'hcafb;
         16'h6688, 16'h6689, 16'h668a, 16'h668b, 16'h668c, 16'h668d, 16'h668e, 16'h668f 	:	val_out <= 16'hcae7;
         16'h6690, 16'h6691, 16'h6692, 16'h6693, 16'h6694, 16'h6695, 16'h6696, 16'h6697 	:	val_out <= 16'hcad2;
         16'h6698, 16'h6699, 16'h669a, 16'h669b, 16'h669c, 16'h669d, 16'h669e, 16'h669f 	:	val_out <= 16'hcabe;
         16'h66a0, 16'h66a1, 16'h66a2, 16'h66a3, 16'h66a4, 16'h66a5, 16'h66a6, 16'h66a7 	:	val_out <= 16'hcaa9;
         16'h66a8, 16'h66a9, 16'h66aa, 16'h66ab, 16'h66ac, 16'h66ad, 16'h66ae, 16'h66af 	:	val_out <= 16'hca95;
         16'h66b0, 16'h66b1, 16'h66b2, 16'h66b3, 16'h66b4, 16'h66b5, 16'h66b6, 16'h66b7 	:	val_out <= 16'hca81;
         16'h66b8, 16'h66b9, 16'h66ba, 16'h66bb, 16'h66bc, 16'h66bd, 16'h66be, 16'h66bf 	:	val_out <= 16'hca6c;
         16'h66c0, 16'h66c1, 16'h66c2, 16'h66c3, 16'h66c4, 16'h66c5, 16'h66c6, 16'h66c7 	:	val_out <= 16'hca58;
         16'h66c8, 16'h66c9, 16'h66ca, 16'h66cb, 16'h66cc, 16'h66cd, 16'h66ce, 16'h66cf 	:	val_out <= 16'hca43;
         16'h66d0, 16'h66d1, 16'h66d2, 16'h66d3, 16'h66d4, 16'h66d5, 16'h66d6, 16'h66d7 	:	val_out <= 16'hca2f;
         16'h66d8, 16'h66d9, 16'h66da, 16'h66db, 16'h66dc, 16'h66dd, 16'h66de, 16'h66df 	:	val_out <= 16'hca1a;
         16'h66e0, 16'h66e1, 16'h66e2, 16'h66e3, 16'h66e4, 16'h66e5, 16'h66e6, 16'h66e7 	:	val_out <= 16'hca06;
         16'h66e8, 16'h66e9, 16'h66ea, 16'h66eb, 16'h66ec, 16'h66ed, 16'h66ee, 16'h66ef 	:	val_out <= 16'hc9f1;
         16'h66f0, 16'h66f1, 16'h66f2, 16'h66f3, 16'h66f4, 16'h66f5, 16'h66f6, 16'h66f7 	:	val_out <= 16'hc9dd;
         16'h66f8, 16'h66f9, 16'h66fa, 16'h66fb, 16'h66fc, 16'h66fd, 16'h66fe, 16'h66ff 	:	val_out <= 16'hc9c8;
         16'h6700, 16'h6701, 16'h6702, 16'h6703, 16'h6704, 16'h6705, 16'h6706, 16'h6707 	:	val_out <= 16'hc9b4;
         16'h6708, 16'h6709, 16'h670a, 16'h670b, 16'h670c, 16'h670d, 16'h670e, 16'h670f 	:	val_out <= 16'hc99f;
         16'h6710, 16'h6711, 16'h6712, 16'h6713, 16'h6714, 16'h6715, 16'h6716, 16'h6717 	:	val_out <= 16'hc98a;
         16'h6718, 16'h6719, 16'h671a, 16'h671b, 16'h671c, 16'h671d, 16'h671e, 16'h671f 	:	val_out <= 16'hc976;
         16'h6720, 16'h6721, 16'h6722, 16'h6723, 16'h6724, 16'h6725, 16'h6726, 16'h6727 	:	val_out <= 16'hc961;
         16'h6728, 16'h6729, 16'h672a, 16'h672b, 16'h672c, 16'h672d, 16'h672e, 16'h672f 	:	val_out <= 16'hc94d;
         16'h6730, 16'h6731, 16'h6732, 16'h6733, 16'h6734, 16'h6735, 16'h6736, 16'h6737 	:	val_out <= 16'hc938;
         16'h6738, 16'h6739, 16'h673a, 16'h673b, 16'h673c, 16'h673d, 16'h673e, 16'h673f 	:	val_out <= 16'hc923;
         16'h6740, 16'h6741, 16'h6742, 16'h6743, 16'h6744, 16'h6745, 16'h6746, 16'h6747 	:	val_out <= 16'hc90f;
         16'h6748, 16'h6749, 16'h674a, 16'h674b, 16'h674c, 16'h674d, 16'h674e, 16'h674f 	:	val_out <= 16'hc8fa;
         16'h6750, 16'h6751, 16'h6752, 16'h6753, 16'h6754, 16'h6755, 16'h6756, 16'h6757 	:	val_out <= 16'hc8e6;
         16'h6758, 16'h6759, 16'h675a, 16'h675b, 16'h675c, 16'h675d, 16'h675e, 16'h675f 	:	val_out <= 16'hc8d1;
         16'h6760, 16'h6761, 16'h6762, 16'h6763, 16'h6764, 16'h6765, 16'h6766, 16'h6767 	:	val_out <= 16'hc8bc;
         16'h6768, 16'h6769, 16'h676a, 16'h676b, 16'h676c, 16'h676d, 16'h676e, 16'h676f 	:	val_out <= 16'hc8a8;
         16'h6770, 16'h6771, 16'h6772, 16'h6773, 16'h6774, 16'h6775, 16'h6776, 16'h6777 	:	val_out <= 16'hc893;
         16'h6778, 16'h6779, 16'h677a, 16'h677b, 16'h677c, 16'h677d, 16'h677e, 16'h677f 	:	val_out <= 16'hc87e;
         16'h6780, 16'h6781, 16'h6782, 16'h6783, 16'h6784, 16'h6785, 16'h6786, 16'h6787 	:	val_out <= 16'hc869;
         16'h6788, 16'h6789, 16'h678a, 16'h678b, 16'h678c, 16'h678d, 16'h678e, 16'h678f 	:	val_out <= 16'hc855;
         16'h6790, 16'h6791, 16'h6792, 16'h6793, 16'h6794, 16'h6795, 16'h6796, 16'h6797 	:	val_out <= 16'hc840;
         16'h6798, 16'h6799, 16'h679a, 16'h679b, 16'h679c, 16'h679d, 16'h679e, 16'h679f 	:	val_out <= 16'hc82b;
         16'h67a0, 16'h67a1, 16'h67a2, 16'h67a3, 16'h67a4, 16'h67a5, 16'h67a6, 16'h67a7 	:	val_out <= 16'hc816;
         16'h67a8, 16'h67a9, 16'h67aa, 16'h67ab, 16'h67ac, 16'h67ad, 16'h67ae, 16'h67af 	:	val_out <= 16'hc802;
         16'h67b0, 16'h67b1, 16'h67b2, 16'h67b3, 16'h67b4, 16'h67b5, 16'h67b6, 16'h67b7 	:	val_out <= 16'hc7ed;
         16'h67b8, 16'h67b9, 16'h67ba, 16'h67bb, 16'h67bc, 16'h67bd, 16'h67be, 16'h67bf 	:	val_out <= 16'hc7d8;
         16'h67c0, 16'h67c1, 16'h67c2, 16'h67c3, 16'h67c4, 16'h67c5, 16'h67c6, 16'h67c7 	:	val_out <= 16'hc7c3;
         16'h67c8, 16'h67c9, 16'h67ca, 16'h67cb, 16'h67cc, 16'h67cd, 16'h67ce, 16'h67cf 	:	val_out <= 16'hc7ae;
         16'h67d0, 16'h67d1, 16'h67d2, 16'h67d3, 16'h67d4, 16'h67d5, 16'h67d6, 16'h67d7 	:	val_out <= 16'hc79a;
         16'h67d8, 16'h67d9, 16'h67da, 16'h67db, 16'h67dc, 16'h67dd, 16'h67de, 16'h67df 	:	val_out <= 16'hc785;
         16'h67e0, 16'h67e1, 16'h67e2, 16'h67e3, 16'h67e4, 16'h67e5, 16'h67e6, 16'h67e7 	:	val_out <= 16'hc770;
         16'h67e8, 16'h67e9, 16'h67ea, 16'h67eb, 16'h67ec, 16'h67ed, 16'h67ee, 16'h67ef 	:	val_out <= 16'hc75b;
         16'h67f0, 16'h67f1, 16'h67f2, 16'h67f3, 16'h67f4, 16'h67f5, 16'h67f6, 16'h67f7 	:	val_out <= 16'hc746;
         16'h67f8, 16'h67f9, 16'h67fa, 16'h67fb, 16'h67fc, 16'h67fd, 16'h67fe, 16'h67ff 	:	val_out <= 16'hc731;
         16'h6800, 16'h6801, 16'h6802, 16'h6803, 16'h6804, 16'h6805, 16'h6806, 16'h6807 	:	val_out <= 16'hc71c;
         16'h6808, 16'h6809, 16'h680a, 16'h680b, 16'h680c, 16'h680d, 16'h680e, 16'h680f 	:	val_out <= 16'hc708;
         16'h6810, 16'h6811, 16'h6812, 16'h6813, 16'h6814, 16'h6815, 16'h6816, 16'h6817 	:	val_out <= 16'hc6f3;
         16'h6818, 16'h6819, 16'h681a, 16'h681b, 16'h681c, 16'h681d, 16'h681e, 16'h681f 	:	val_out <= 16'hc6de;
         16'h6820, 16'h6821, 16'h6822, 16'h6823, 16'h6824, 16'h6825, 16'h6826, 16'h6827 	:	val_out <= 16'hc6c9;
         16'h6828, 16'h6829, 16'h682a, 16'h682b, 16'h682c, 16'h682d, 16'h682e, 16'h682f 	:	val_out <= 16'hc6b4;
         16'h6830, 16'h6831, 16'h6832, 16'h6833, 16'h6834, 16'h6835, 16'h6836, 16'h6837 	:	val_out <= 16'hc69f;
         16'h6838, 16'h6839, 16'h683a, 16'h683b, 16'h683c, 16'h683d, 16'h683e, 16'h683f 	:	val_out <= 16'hc68a;
         16'h6840, 16'h6841, 16'h6842, 16'h6843, 16'h6844, 16'h6845, 16'h6846, 16'h6847 	:	val_out <= 16'hc675;
         16'h6848, 16'h6849, 16'h684a, 16'h684b, 16'h684c, 16'h684d, 16'h684e, 16'h684f 	:	val_out <= 16'hc660;
         16'h6850, 16'h6851, 16'h6852, 16'h6853, 16'h6854, 16'h6855, 16'h6856, 16'h6857 	:	val_out <= 16'hc64b;
         16'h6858, 16'h6859, 16'h685a, 16'h685b, 16'h685c, 16'h685d, 16'h685e, 16'h685f 	:	val_out <= 16'hc636;
         16'h6860, 16'h6861, 16'h6862, 16'h6863, 16'h6864, 16'h6865, 16'h6866, 16'h6867 	:	val_out <= 16'hc621;
         16'h6868, 16'h6869, 16'h686a, 16'h686b, 16'h686c, 16'h686d, 16'h686e, 16'h686f 	:	val_out <= 16'hc60c;
         16'h6870, 16'h6871, 16'h6872, 16'h6873, 16'h6874, 16'h6875, 16'h6876, 16'h6877 	:	val_out <= 16'hc5f7;
         16'h6878, 16'h6879, 16'h687a, 16'h687b, 16'h687c, 16'h687d, 16'h687e, 16'h687f 	:	val_out <= 16'hc5e2;
         16'h6880, 16'h6881, 16'h6882, 16'h6883, 16'h6884, 16'h6885, 16'h6886, 16'h6887 	:	val_out <= 16'hc5cd;
         16'h6888, 16'h6889, 16'h688a, 16'h688b, 16'h688c, 16'h688d, 16'h688e, 16'h688f 	:	val_out <= 16'hc5b8;
         16'h6890, 16'h6891, 16'h6892, 16'h6893, 16'h6894, 16'h6895, 16'h6896, 16'h6897 	:	val_out <= 16'hc5a3;
         16'h6898, 16'h6899, 16'h689a, 16'h689b, 16'h689c, 16'h689d, 16'h689e, 16'h689f 	:	val_out <= 16'hc58d;
         16'h68a0, 16'h68a1, 16'h68a2, 16'h68a3, 16'h68a4, 16'h68a5, 16'h68a6, 16'h68a7 	:	val_out <= 16'hc578;
         16'h68a8, 16'h68a9, 16'h68aa, 16'h68ab, 16'h68ac, 16'h68ad, 16'h68ae, 16'h68af 	:	val_out <= 16'hc563;
         16'h68b0, 16'h68b1, 16'h68b2, 16'h68b3, 16'h68b4, 16'h68b5, 16'h68b6, 16'h68b7 	:	val_out <= 16'hc54e;
         16'h68b8, 16'h68b9, 16'h68ba, 16'h68bb, 16'h68bc, 16'h68bd, 16'h68be, 16'h68bf 	:	val_out <= 16'hc539;
         16'h68c0, 16'h68c1, 16'h68c2, 16'h68c3, 16'h68c4, 16'h68c5, 16'h68c6, 16'h68c7 	:	val_out <= 16'hc524;
         16'h68c8, 16'h68c9, 16'h68ca, 16'h68cb, 16'h68cc, 16'h68cd, 16'h68ce, 16'h68cf 	:	val_out <= 16'hc50f;
         16'h68d0, 16'h68d1, 16'h68d2, 16'h68d3, 16'h68d4, 16'h68d5, 16'h68d6, 16'h68d7 	:	val_out <= 16'hc4fa;
         16'h68d8, 16'h68d9, 16'h68da, 16'h68db, 16'h68dc, 16'h68dd, 16'h68de, 16'h68df 	:	val_out <= 16'hc4e4;
         16'h68e0, 16'h68e1, 16'h68e2, 16'h68e3, 16'h68e4, 16'h68e5, 16'h68e6, 16'h68e7 	:	val_out <= 16'hc4cf;
         16'h68e8, 16'h68e9, 16'h68ea, 16'h68eb, 16'h68ec, 16'h68ed, 16'h68ee, 16'h68ef 	:	val_out <= 16'hc4ba;
         16'h68f0, 16'h68f1, 16'h68f2, 16'h68f3, 16'h68f4, 16'h68f5, 16'h68f6, 16'h68f7 	:	val_out <= 16'hc4a5;
         16'h68f8, 16'h68f9, 16'h68fa, 16'h68fb, 16'h68fc, 16'h68fd, 16'h68fe, 16'h68ff 	:	val_out <= 16'hc490;
         16'h6900, 16'h6901, 16'h6902, 16'h6903, 16'h6904, 16'h6905, 16'h6906, 16'h6907 	:	val_out <= 16'hc47a;
         16'h6908, 16'h6909, 16'h690a, 16'h690b, 16'h690c, 16'h690d, 16'h690e, 16'h690f 	:	val_out <= 16'hc465;
         16'h6910, 16'h6911, 16'h6912, 16'h6913, 16'h6914, 16'h6915, 16'h6916, 16'h6917 	:	val_out <= 16'hc450;
         16'h6918, 16'h6919, 16'h691a, 16'h691b, 16'h691c, 16'h691d, 16'h691e, 16'h691f 	:	val_out <= 16'hc43b;
         16'h6920, 16'h6921, 16'h6922, 16'h6923, 16'h6924, 16'h6925, 16'h6926, 16'h6927 	:	val_out <= 16'hc425;
         16'h6928, 16'h6929, 16'h692a, 16'h692b, 16'h692c, 16'h692d, 16'h692e, 16'h692f 	:	val_out <= 16'hc410;
         16'h6930, 16'h6931, 16'h6932, 16'h6933, 16'h6934, 16'h6935, 16'h6936, 16'h6937 	:	val_out <= 16'hc3fb;
         16'h6938, 16'h6939, 16'h693a, 16'h693b, 16'h693c, 16'h693d, 16'h693e, 16'h693f 	:	val_out <= 16'hc3e5;
         16'h6940, 16'h6941, 16'h6942, 16'h6943, 16'h6944, 16'h6945, 16'h6946, 16'h6947 	:	val_out <= 16'hc3d0;
         16'h6948, 16'h6949, 16'h694a, 16'h694b, 16'h694c, 16'h694d, 16'h694e, 16'h694f 	:	val_out <= 16'hc3bb;
         16'h6950, 16'h6951, 16'h6952, 16'h6953, 16'h6954, 16'h6955, 16'h6956, 16'h6957 	:	val_out <= 16'hc3a5;
         16'h6958, 16'h6959, 16'h695a, 16'h695b, 16'h695c, 16'h695d, 16'h695e, 16'h695f 	:	val_out <= 16'hc390;
         16'h6960, 16'h6961, 16'h6962, 16'h6963, 16'h6964, 16'h6965, 16'h6966, 16'h6967 	:	val_out <= 16'hc37b;
         16'h6968, 16'h6969, 16'h696a, 16'h696b, 16'h696c, 16'h696d, 16'h696e, 16'h696f 	:	val_out <= 16'hc365;
         16'h6970, 16'h6971, 16'h6972, 16'h6973, 16'h6974, 16'h6975, 16'h6976, 16'h6977 	:	val_out <= 16'hc350;
         16'h6978, 16'h6979, 16'h697a, 16'h697b, 16'h697c, 16'h697d, 16'h697e, 16'h697f 	:	val_out <= 16'hc33b;
         16'h6980, 16'h6981, 16'h6982, 16'h6983, 16'h6984, 16'h6985, 16'h6986, 16'h6987 	:	val_out <= 16'hc325;
         16'h6988, 16'h6989, 16'h698a, 16'h698b, 16'h698c, 16'h698d, 16'h698e, 16'h698f 	:	val_out <= 16'hc310;
         16'h6990, 16'h6991, 16'h6992, 16'h6993, 16'h6994, 16'h6995, 16'h6996, 16'h6997 	:	val_out <= 16'hc2fa;
         16'h6998, 16'h6999, 16'h699a, 16'h699b, 16'h699c, 16'h699d, 16'h699e, 16'h699f 	:	val_out <= 16'hc2e5;
         16'h69a0, 16'h69a1, 16'h69a2, 16'h69a3, 16'h69a4, 16'h69a5, 16'h69a6, 16'h69a7 	:	val_out <= 16'hc2d0;
         16'h69a8, 16'h69a9, 16'h69aa, 16'h69ab, 16'h69ac, 16'h69ad, 16'h69ae, 16'h69af 	:	val_out <= 16'hc2ba;
         16'h69b0, 16'h69b1, 16'h69b2, 16'h69b3, 16'h69b4, 16'h69b5, 16'h69b6, 16'h69b7 	:	val_out <= 16'hc2a5;
         16'h69b8, 16'h69b9, 16'h69ba, 16'h69bb, 16'h69bc, 16'h69bd, 16'h69be, 16'h69bf 	:	val_out <= 16'hc28f;
         16'h69c0, 16'h69c1, 16'h69c2, 16'h69c3, 16'h69c4, 16'h69c5, 16'h69c6, 16'h69c7 	:	val_out <= 16'hc27a;
         16'h69c8, 16'h69c9, 16'h69ca, 16'h69cb, 16'h69cc, 16'h69cd, 16'h69ce, 16'h69cf 	:	val_out <= 16'hc264;
         16'h69d0, 16'h69d1, 16'h69d2, 16'h69d3, 16'h69d4, 16'h69d5, 16'h69d6, 16'h69d7 	:	val_out <= 16'hc24f;
         16'h69d8, 16'h69d9, 16'h69da, 16'h69db, 16'h69dc, 16'h69dd, 16'h69de, 16'h69df 	:	val_out <= 16'hc239;
         16'h69e0, 16'h69e1, 16'h69e2, 16'h69e3, 16'h69e4, 16'h69e5, 16'h69e6, 16'h69e7 	:	val_out <= 16'hc224;
         16'h69e8, 16'h69e9, 16'h69ea, 16'h69eb, 16'h69ec, 16'h69ed, 16'h69ee, 16'h69ef 	:	val_out <= 16'hc20e;
         16'h69f0, 16'h69f1, 16'h69f2, 16'h69f3, 16'h69f4, 16'h69f5, 16'h69f6, 16'h69f7 	:	val_out <= 16'hc1f9;
         16'h69f8, 16'h69f9, 16'h69fa, 16'h69fb, 16'h69fc, 16'h69fd, 16'h69fe, 16'h69ff 	:	val_out <= 16'hc1e3;
         16'h6a00, 16'h6a01, 16'h6a02, 16'h6a03, 16'h6a04, 16'h6a05, 16'h6a06, 16'h6a07 	:	val_out <= 16'hc1ce;
         16'h6a08, 16'h6a09, 16'h6a0a, 16'h6a0b, 16'h6a0c, 16'h6a0d, 16'h6a0e, 16'h6a0f 	:	val_out <= 16'hc1b8;
         16'h6a10, 16'h6a11, 16'h6a12, 16'h6a13, 16'h6a14, 16'h6a15, 16'h6a16, 16'h6a17 	:	val_out <= 16'hc1a2;
         16'h6a18, 16'h6a19, 16'h6a1a, 16'h6a1b, 16'h6a1c, 16'h6a1d, 16'h6a1e, 16'h6a1f 	:	val_out <= 16'hc18d;
         16'h6a20, 16'h6a21, 16'h6a22, 16'h6a23, 16'h6a24, 16'h6a25, 16'h6a26, 16'h6a27 	:	val_out <= 16'hc177;
         16'h6a28, 16'h6a29, 16'h6a2a, 16'h6a2b, 16'h6a2c, 16'h6a2d, 16'h6a2e, 16'h6a2f 	:	val_out <= 16'hc162;
         16'h6a30, 16'h6a31, 16'h6a32, 16'h6a33, 16'h6a34, 16'h6a35, 16'h6a36, 16'h6a37 	:	val_out <= 16'hc14c;
         16'h6a38, 16'h6a39, 16'h6a3a, 16'h6a3b, 16'h6a3c, 16'h6a3d, 16'h6a3e, 16'h6a3f 	:	val_out <= 16'hc136;
         16'h6a40, 16'h6a41, 16'h6a42, 16'h6a43, 16'h6a44, 16'h6a45, 16'h6a46, 16'h6a47 	:	val_out <= 16'hc121;
         16'h6a48, 16'h6a49, 16'h6a4a, 16'h6a4b, 16'h6a4c, 16'h6a4d, 16'h6a4e, 16'h6a4f 	:	val_out <= 16'hc10b;
         16'h6a50, 16'h6a51, 16'h6a52, 16'h6a53, 16'h6a54, 16'h6a55, 16'h6a56, 16'h6a57 	:	val_out <= 16'hc0f6;
         16'h6a58, 16'h6a59, 16'h6a5a, 16'h6a5b, 16'h6a5c, 16'h6a5d, 16'h6a5e, 16'h6a5f 	:	val_out <= 16'hc0e0;
         16'h6a60, 16'h6a61, 16'h6a62, 16'h6a63, 16'h6a64, 16'h6a65, 16'h6a66, 16'h6a67 	:	val_out <= 16'hc0ca;
         16'h6a68, 16'h6a69, 16'h6a6a, 16'h6a6b, 16'h6a6c, 16'h6a6d, 16'h6a6e, 16'h6a6f 	:	val_out <= 16'hc0b5;
         16'h6a70, 16'h6a71, 16'h6a72, 16'h6a73, 16'h6a74, 16'h6a75, 16'h6a76, 16'h6a77 	:	val_out <= 16'hc09f;
         16'h6a78, 16'h6a79, 16'h6a7a, 16'h6a7b, 16'h6a7c, 16'h6a7d, 16'h6a7e, 16'h6a7f 	:	val_out <= 16'hc089;
         16'h6a80, 16'h6a81, 16'h6a82, 16'h6a83, 16'h6a84, 16'h6a85, 16'h6a86, 16'h6a87 	:	val_out <= 16'hc073;
         16'h6a88, 16'h6a89, 16'h6a8a, 16'h6a8b, 16'h6a8c, 16'h6a8d, 16'h6a8e, 16'h6a8f 	:	val_out <= 16'hc05e;
         16'h6a90, 16'h6a91, 16'h6a92, 16'h6a93, 16'h6a94, 16'h6a95, 16'h6a96, 16'h6a97 	:	val_out <= 16'hc048;
         16'h6a98, 16'h6a99, 16'h6a9a, 16'h6a9b, 16'h6a9c, 16'h6a9d, 16'h6a9e, 16'h6a9f 	:	val_out <= 16'hc032;
         16'h6aa0, 16'h6aa1, 16'h6aa2, 16'h6aa3, 16'h6aa4, 16'h6aa5, 16'h6aa6, 16'h6aa7 	:	val_out <= 16'hc01d;
         16'h6aa8, 16'h6aa9, 16'h6aaa, 16'h6aab, 16'h6aac, 16'h6aad, 16'h6aae, 16'h6aaf 	:	val_out <= 16'hc007;
         16'h6ab0, 16'h6ab1, 16'h6ab2, 16'h6ab3, 16'h6ab4, 16'h6ab5, 16'h6ab6, 16'h6ab7 	:	val_out <= 16'hbff1;
         16'h6ab8, 16'h6ab9, 16'h6aba, 16'h6abb, 16'h6abc, 16'h6abd, 16'h6abe, 16'h6abf 	:	val_out <= 16'hbfdb;
         16'h6ac0, 16'h6ac1, 16'h6ac2, 16'h6ac3, 16'h6ac4, 16'h6ac5, 16'h6ac6, 16'h6ac7 	:	val_out <= 16'hbfc5;
         16'h6ac8, 16'h6ac9, 16'h6aca, 16'h6acb, 16'h6acc, 16'h6acd, 16'h6ace, 16'h6acf 	:	val_out <= 16'hbfb0;
         16'h6ad0, 16'h6ad1, 16'h6ad2, 16'h6ad3, 16'h6ad4, 16'h6ad5, 16'h6ad6, 16'h6ad7 	:	val_out <= 16'hbf9a;
         16'h6ad8, 16'h6ad9, 16'h6ada, 16'h6adb, 16'h6adc, 16'h6add, 16'h6ade, 16'h6adf 	:	val_out <= 16'hbf84;
         16'h6ae0, 16'h6ae1, 16'h6ae2, 16'h6ae3, 16'h6ae4, 16'h6ae5, 16'h6ae6, 16'h6ae7 	:	val_out <= 16'hbf6e;
         16'h6ae8, 16'h6ae9, 16'h6aea, 16'h6aeb, 16'h6aec, 16'h6aed, 16'h6aee, 16'h6aef 	:	val_out <= 16'hbf58;
         16'h6af0, 16'h6af1, 16'h6af2, 16'h6af3, 16'h6af4, 16'h6af5, 16'h6af6, 16'h6af7 	:	val_out <= 16'hbf43;
         16'h6af8, 16'h6af9, 16'h6afa, 16'h6afb, 16'h6afc, 16'h6afd, 16'h6afe, 16'h6aff 	:	val_out <= 16'hbf2d;
         16'h6b00, 16'h6b01, 16'h6b02, 16'h6b03, 16'h6b04, 16'h6b05, 16'h6b06, 16'h6b07 	:	val_out <= 16'hbf17;
         16'h6b08, 16'h6b09, 16'h6b0a, 16'h6b0b, 16'h6b0c, 16'h6b0d, 16'h6b0e, 16'h6b0f 	:	val_out <= 16'hbf01;
         16'h6b10, 16'h6b11, 16'h6b12, 16'h6b13, 16'h6b14, 16'h6b15, 16'h6b16, 16'h6b17 	:	val_out <= 16'hbeeb;
         16'h6b18, 16'h6b19, 16'h6b1a, 16'h6b1b, 16'h6b1c, 16'h6b1d, 16'h6b1e, 16'h6b1f 	:	val_out <= 16'hbed5;
         16'h6b20, 16'h6b21, 16'h6b22, 16'h6b23, 16'h6b24, 16'h6b25, 16'h6b26, 16'h6b27 	:	val_out <= 16'hbebf;
         16'h6b28, 16'h6b29, 16'h6b2a, 16'h6b2b, 16'h6b2c, 16'h6b2d, 16'h6b2e, 16'h6b2f 	:	val_out <= 16'hbea9;
         16'h6b30, 16'h6b31, 16'h6b32, 16'h6b33, 16'h6b34, 16'h6b35, 16'h6b36, 16'h6b37 	:	val_out <= 16'hbe93;
         16'h6b38, 16'h6b39, 16'h6b3a, 16'h6b3b, 16'h6b3c, 16'h6b3d, 16'h6b3e, 16'h6b3f 	:	val_out <= 16'hbe7d;
         16'h6b40, 16'h6b41, 16'h6b42, 16'h6b43, 16'h6b44, 16'h6b45, 16'h6b46, 16'h6b47 	:	val_out <= 16'hbe68;
         16'h6b48, 16'h6b49, 16'h6b4a, 16'h6b4b, 16'h6b4c, 16'h6b4d, 16'h6b4e, 16'h6b4f 	:	val_out <= 16'hbe52;
         16'h6b50, 16'h6b51, 16'h6b52, 16'h6b53, 16'h6b54, 16'h6b55, 16'h6b56, 16'h6b57 	:	val_out <= 16'hbe3c;
         16'h6b58, 16'h6b59, 16'h6b5a, 16'h6b5b, 16'h6b5c, 16'h6b5d, 16'h6b5e, 16'h6b5f 	:	val_out <= 16'hbe26;
         16'h6b60, 16'h6b61, 16'h6b62, 16'h6b63, 16'h6b64, 16'h6b65, 16'h6b66, 16'h6b67 	:	val_out <= 16'hbe10;
         16'h6b68, 16'h6b69, 16'h6b6a, 16'h6b6b, 16'h6b6c, 16'h6b6d, 16'h6b6e, 16'h6b6f 	:	val_out <= 16'hbdfa;
         16'h6b70, 16'h6b71, 16'h6b72, 16'h6b73, 16'h6b74, 16'h6b75, 16'h6b76, 16'h6b77 	:	val_out <= 16'hbde4;
         16'h6b78, 16'h6b79, 16'h6b7a, 16'h6b7b, 16'h6b7c, 16'h6b7d, 16'h6b7e, 16'h6b7f 	:	val_out <= 16'hbdce;
         16'h6b80, 16'h6b81, 16'h6b82, 16'h6b83, 16'h6b84, 16'h6b85, 16'h6b86, 16'h6b87 	:	val_out <= 16'hbdb8;
         16'h6b88, 16'h6b89, 16'h6b8a, 16'h6b8b, 16'h6b8c, 16'h6b8d, 16'h6b8e, 16'h6b8f 	:	val_out <= 16'hbda2;
         16'h6b90, 16'h6b91, 16'h6b92, 16'h6b93, 16'h6b94, 16'h6b95, 16'h6b96, 16'h6b97 	:	val_out <= 16'hbd8c;
         16'h6b98, 16'h6b99, 16'h6b9a, 16'h6b9b, 16'h6b9c, 16'h6b9d, 16'h6b9e, 16'h6b9f 	:	val_out <= 16'hbd76;
         16'h6ba0, 16'h6ba1, 16'h6ba2, 16'h6ba3, 16'h6ba4, 16'h6ba5, 16'h6ba6, 16'h6ba7 	:	val_out <= 16'hbd60;
         16'h6ba8, 16'h6ba9, 16'h6baa, 16'h6bab, 16'h6bac, 16'h6bad, 16'h6bae, 16'h6baf 	:	val_out <= 16'hbd49;
         16'h6bb0, 16'h6bb1, 16'h6bb2, 16'h6bb3, 16'h6bb4, 16'h6bb5, 16'h6bb6, 16'h6bb7 	:	val_out <= 16'hbd33;
         16'h6bb8, 16'h6bb9, 16'h6bba, 16'h6bbb, 16'h6bbc, 16'h6bbd, 16'h6bbe, 16'h6bbf 	:	val_out <= 16'hbd1d;
         16'h6bc0, 16'h6bc1, 16'h6bc2, 16'h6bc3, 16'h6bc4, 16'h6bc5, 16'h6bc6, 16'h6bc7 	:	val_out <= 16'hbd07;
         16'h6bc8, 16'h6bc9, 16'h6bca, 16'h6bcb, 16'h6bcc, 16'h6bcd, 16'h6bce, 16'h6bcf 	:	val_out <= 16'hbcf1;
         16'h6bd0, 16'h6bd1, 16'h6bd2, 16'h6bd3, 16'h6bd4, 16'h6bd5, 16'h6bd6, 16'h6bd7 	:	val_out <= 16'hbcdb;
         16'h6bd8, 16'h6bd9, 16'h6bda, 16'h6bdb, 16'h6bdc, 16'h6bdd, 16'h6bde, 16'h6bdf 	:	val_out <= 16'hbcc5;
         16'h6be0, 16'h6be1, 16'h6be2, 16'h6be3, 16'h6be4, 16'h6be5, 16'h6be6, 16'h6be7 	:	val_out <= 16'hbcaf;
         16'h6be8, 16'h6be9, 16'h6bea, 16'h6beb, 16'h6bec, 16'h6bed, 16'h6bee, 16'h6bef 	:	val_out <= 16'hbc99;
         16'h6bf0, 16'h6bf1, 16'h6bf2, 16'h6bf3, 16'h6bf4, 16'h6bf5, 16'h6bf6, 16'h6bf7 	:	val_out <= 16'hbc83;
         16'h6bf8, 16'h6bf9, 16'h6bfa, 16'h6bfb, 16'h6bfc, 16'h6bfd, 16'h6bfe, 16'h6bff 	:	val_out <= 16'hbc6c;
         16'h6c00, 16'h6c01, 16'h6c02, 16'h6c03, 16'h6c04, 16'h6c05, 16'h6c06, 16'h6c07 	:	val_out <= 16'hbc56;
         16'h6c08, 16'h6c09, 16'h6c0a, 16'h6c0b, 16'h6c0c, 16'h6c0d, 16'h6c0e, 16'h6c0f 	:	val_out <= 16'hbc40;
         16'h6c10, 16'h6c11, 16'h6c12, 16'h6c13, 16'h6c14, 16'h6c15, 16'h6c16, 16'h6c17 	:	val_out <= 16'hbc2a;
         16'h6c18, 16'h6c19, 16'h6c1a, 16'h6c1b, 16'h6c1c, 16'h6c1d, 16'h6c1e, 16'h6c1f 	:	val_out <= 16'hbc14;
         16'h6c20, 16'h6c21, 16'h6c22, 16'h6c23, 16'h6c24, 16'h6c25, 16'h6c26, 16'h6c27 	:	val_out <= 16'hbbfd;
         16'h6c28, 16'h6c29, 16'h6c2a, 16'h6c2b, 16'h6c2c, 16'h6c2d, 16'h6c2e, 16'h6c2f 	:	val_out <= 16'hbbe7;
         16'h6c30, 16'h6c31, 16'h6c32, 16'h6c33, 16'h6c34, 16'h6c35, 16'h6c36, 16'h6c37 	:	val_out <= 16'hbbd1;
         16'h6c38, 16'h6c39, 16'h6c3a, 16'h6c3b, 16'h6c3c, 16'h6c3d, 16'h6c3e, 16'h6c3f 	:	val_out <= 16'hbbbb;
         16'h6c40, 16'h6c41, 16'h6c42, 16'h6c43, 16'h6c44, 16'h6c45, 16'h6c46, 16'h6c47 	:	val_out <= 16'hbba5;
         16'h6c48, 16'h6c49, 16'h6c4a, 16'h6c4b, 16'h6c4c, 16'h6c4d, 16'h6c4e, 16'h6c4f 	:	val_out <= 16'hbb8e;
         16'h6c50, 16'h6c51, 16'h6c52, 16'h6c53, 16'h6c54, 16'h6c55, 16'h6c56, 16'h6c57 	:	val_out <= 16'hbb78;
         16'h6c58, 16'h6c59, 16'h6c5a, 16'h6c5b, 16'h6c5c, 16'h6c5d, 16'h6c5e, 16'h6c5f 	:	val_out <= 16'hbb62;
         16'h6c60, 16'h6c61, 16'h6c62, 16'h6c63, 16'h6c64, 16'h6c65, 16'h6c66, 16'h6c67 	:	val_out <= 16'hbb4c;
         16'h6c68, 16'h6c69, 16'h6c6a, 16'h6c6b, 16'h6c6c, 16'h6c6d, 16'h6c6e, 16'h6c6f 	:	val_out <= 16'hbb35;
         16'h6c70, 16'h6c71, 16'h6c72, 16'h6c73, 16'h6c74, 16'h6c75, 16'h6c76, 16'h6c77 	:	val_out <= 16'hbb1f;
         16'h6c78, 16'h6c79, 16'h6c7a, 16'h6c7b, 16'h6c7c, 16'h6c7d, 16'h6c7e, 16'h6c7f 	:	val_out <= 16'hbb09;
         16'h6c80, 16'h6c81, 16'h6c82, 16'h6c83, 16'h6c84, 16'h6c85, 16'h6c86, 16'h6c87 	:	val_out <= 16'hbaf2;
         16'h6c88, 16'h6c89, 16'h6c8a, 16'h6c8b, 16'h6c8c, 16'h6c8d, 16'h6c8e, 16'h6c8f 	:	val_out <= 16'hbadc;
         16'h6c90, 16'h6c91, 16'h6c92, 16'h6c93, 16'h6c94, 16'h6c95, 16'h6c96, 16'h6c97 	:	val_out <= 16'hbac6;
         16'h6c98, 16'h6c99, 16'h6c9a, 16'h6c9b, 16'h6c9c, 16'h6c9d, 16'h6c9e, 16'h6c9f 	:	val_out <= 16'hbaaf;
         16'h6ca0, 16'h6ca1, 16'h6ca2, 16'h6ca3, 16'h6ca4, 16'h6ca5, 16'h6ca6, 16'h6ca7 	:	val_out <= 16'hba99;
         16'h6ca8, 16'h6ca9, 16'h6caa, 16'h6cab, 16'h6cac, 16'h6cad, 16'h6cae, 16'h6caf 	:	val_out <= 16'hba83;
         16'h6cb0, 16'h6cb1, 16'h6cb2, 16'h6cb3, 16'h6cb4, 16'h6cb5, 16'h6cb6, 16'h6cb7 	:	val_out <= 16'hba6c;
         16'h6cb8, 16'h6cb9, 16'h6cba, 16'h6cbb, 16'h6cbc, 16'h6cbd, 16'h6cbe, 16'h6cbf 	:	val_out <= 16'hba56;
         16'h6cc0, 16'h6cc1, 16'h6cc2, 16'h6cc3, 16'h6cc4, 16'h6cc5, 16'h6cc6, 16'h6cc7 	:	val_out <= 16'hba40;
         16'h6cc8, 16'h6cc9, 16'h6cca, 16'h6ccb, 16'h6ccc, 16'h6ccd, 16'h6cce, 16'h6ccf 	:	val_out <= 16'hba29;
         16'h6cd0, 16'h6cd1, 16'h6cd2, 16'h6cd3, 16'h6cd4, 16'h6cd5, 16'h6cd6, 16'h6cd7 	:	val_out <= 16'hba13;
         16'h6cd8, 16'h6cd9, 16'h6cda, 16'h6cdb, 16'h6cdc, 16'h6cdd, 16'h6cde, 16'h6cdf 	:	val_out <= 16'hb9fd;
         16'h6ce0, 16'h6ce1, 16'h6ce2, 16'h6ce3, 16'h6ce4, 16'h6ce5, 16'h6ce6, 16'h6ce7 	:	val_out <= 16'hb9e6;
         16'h6ce8, 16'h6ce9, 16'h6cea, 16'h6ceb, 16'h6cec, 16'h6ced, 16'h6cee, 16'h6cef 	:	val_out <= 16'hb9d0;
         16'h6cf0, 16'h6cf1, 16'h6cf2, 16'h6cf3, 16'h6cf4, 16'h6cf5, 16'h6cf6, 16'h6cf7 	:	val_out <= 16'hb9b9;
         16'h6cf8, 16'h6cf9, 16'h6cfa, 16'h6cfb, 16'h6cfc, 16'h6cfd, 16'h6cfe, 16'h6cff 	:	val_out <= 16'hb9a3;
         16'h6d00, 16'h6d01, 16'h6d02, 16'h6d03, 16'h6d04, 16'h6d05, 16'h6d06, 16'h6d07 	:	val_out <= 16'hb98c;
         16'h6d08, 16'h6d09, 16'h6d0a, 16'h6d0b, 16'h6d0c, 16'h6d0d, 16'h6d0e, 16'h6d0f 	:	val_out <= 16'hb976;
         16'h6d10, 16'h6d11, 16'h6d12, 16'h6d13, 16'h6d14, 16'h6d15, 16'h6d16, 16'h6d17 	:	val_out <= 16'hb95f;
         16'h6d18, 16'h6d19, 16'h6d1a, 16'h6d1b, 16'h6d1c, 16'h6d1d, 16'h6d1e, 16'h6d1f 	:	val_out <= 16'hb949;
         16'h6d20, 16'h6d21, 16'h6d22, 16'h6d23, 16'h6d24, 16'h6d25, 16'h6d26, 16'h6d27 	:	val_out <= 16'hb932;
         16'h6d28, 16'h6d29, 16'h6d2a, 16'h6d2b, 16'h6d2c, 16'h6d2d, 16'h6d2e, 16'h6d2f 	:	val_out <= 16'hb91c;
         16'h6d30, 16'h6d31, 16'h6d32, 16'h6d33, 16'h6d34, 16'h6d35, 16'h6d36, 16'h6d37 	:	val_out <= 16'hb906;
         16'h6d38, 16'h6d39, 16'h6d3a, 16'h6d3b, 16'h6d3c, 16'h6d3d, 16'h6d3e, 16'h6d3f 	:	val_out <= 16'hb8ef;
         16'h6d40, 16'h6d41, 16'h6d42, 16'h6d43, 16'h6d44, 16'h6d45, 16'h6d46, 16'h6d47 	:	val_out <= 16'hb8d8;
         16'h6d48, 16'h6d49, 16'h6d4a, 16'h6d4b, 16'h6d4c, 16'h6d4d, 16'h6d4e, 16'h6d4f 	:	val_out <= 16'hb8c2;
         16'h6d50, 16'h6d51, 16'h6d52, 16'h6d53, 16'h6d54, 16'h6d55, 16'h6d56, 16'h6d57 	:	val_out <= 16'hb8ab;
         16'h6d58, 16'h6d59, 16'h6d5a, 16'h6d5b, 16'h6d5c, 16'h6d5d, 16'h6d5e, 16'h6d5f 	:	val_out <= 16'hb895;
         16'h6d60, 16'h6d61, 16'h6d62, 16'h6d63, 16'h6d64, 16'h6d65, 16'h6d66, 16'h6d67 	:	val_out <= 16'hb87e;
         16'h6d68, 16'h6d69, 16'h6d6a, 16'h6d6b, 16'h6d6c, 16'h6d6d, 16'h6d6e, 16'h6d6f 	:	val_out <= 16'hb868;
         16'h6d70, 16'h6d71, 16'h6d72, 16'h6d73, 16'h6d74, 16'h6d75, 16'h6d76, 16'h6d77 	:	val_out <= 16'hb851;
         16'h6d78, 16'h6d79, 16'h6d7a, 16'h6d7b, 16'h6d7c, 16'h6d7d, 16'h6d7e, 16'h6d7f 	:	val_out <= 16'hb83b;
         16'h6d80, 16'h6d81, 16'h6d82, 16'h6d83, 16'h6d84, 16'h6d85, 16'h6d86, 16'h6d87 	:	val_out <= 16'hb824;
         16'h6d88, 16'h6d89, 16'h6d8a, 16'h6d8b, 16'h6d8c, 16'h6d8d, 16'h6d8e, 16'h6d8f 	:	val_out <= 16'hb80d;
         16'h6d90, 16'h6d91, 16'h6d92, 16'h6d93, 16'h6d94, 16'h6d95, 16'h6d96, 16'h6d97 	:	val_out <= 16'hb7f7;
         16'h6d98, 16'h6d99, 16'h6d9a, 16'h6d9b, 16'h6d9c, 16'h6d9d, 16'h6d9e, 16'h6d9f 	:	val_out <= 16'hb7e0;
         16'h6da0, 16'h6da1, 16'h6da2, 16'h6da3, 16'h6da4, 16'h6da5, 16'h6da6, 16'h6da7 	:	val_out <= 16'hb7ca;
         16'h6da8, 16'h6da9, 16'h6daa, 16'h6dab, 16'h6dac, 16'h6dad, 16'h6dae, 16'h6daf 	:	val_out <= 16'hb7b3;
         16'h6db0, 16'h6db1, 16'h6db2, 16'h6db3, 16'h6db4, 16'h6db5, 16'h6db6, 16'h6db7 	:	val_out <= 16'hb79c;
         16'h6db8, 16'h6db9, 16'h6dba, 16'h6dbb, 16'h6dbc, 16'h6dbd, 16'h6dbe, 16'h6dbf 	:	val_out <= 16'hb786;
         16'h6dc0, 16'h6dc1, 16'h6dc2, 16'h6dc3, 16'h6dc4, 16'h6dc5, 16'h6dc6, 16'h6dc7 	:	val_out <= 16'hb76f;
         16'h6dc8, 16'h6dc9, 16'h6dca, 16'h6dcb, 16'h6dcc, 16'h6dcd, 16'h6dce, 16'h6dcf 	:	val_out <= 16'hb758;
         16'h6dd0, 16'h6dd1, 16'h6dd2, 16'h6dd3, 16'h6dd4, 16'h6dd5, 16'h6dd6, 16'h6dd7 	:	val_out <= 16'hb742;
         16'h6dd8, 16'h6dd9, 16'h6dda, 16'h6ddb, 16'h6ddc, 16'h6ddd, 16'h6dde, 16'h6ddf 	:	val_out <= 16'hb72b;
         16'h6de0, 16'h6de1, 16'h6de2, 16'h6de3, 16'h6de4, 16'h6de5, 16'h6de6, 16'h6de7 	:	val_out <= 16'hb714;
         16'h6de8, 16'h6de9, 16'h6dea, 16'h6deb, 16'h6dec, 16'h6ded, 16'h6dee, 16'h6def 	:	val_out <= 16'hb6fe;
         16'h6df0, 16'h6df1, 16'h6df2, 16'h6df3, 16'h6df4, 16'h6df5, 16'h6df6, 16'h6df7 	:	val_out <= 16'hb6e7;
         16'h6df8, 16'h6df9, 16'h6dfa, 16'h6dfb, 16'h6dfc, 16'h6dfd, 16'h6dfe, 16'h6dff 	:	val_out <= 16'hb6d0;
         16'h6e00, 16'h6e01, 16'h6e02, 16'h6e03, 16'h6e04, 16'h6e05, 16'h6e06, 16'h6e07 	:	val_out <= 16'hb6ba;
         16'h6e08, 16'h6e09, 16'h6e0a, 16'h6e0b, 16'h6e0c, 16'h6e0d, 16'h6e0e, 16'h6e0f 	:	val_out <= 16'hb6a3;
         16'h6e10, 16'h6e11, 16'h6e12, 16'h6e13, 16'h6e14, 16'h6e15, 16'h6e16, 16'h6e17 	:	val_out <= 16'hb68c;
         16'h6e18, 16'h6e19, 16'h6e1a, 16'h6e1b, 16'h6e1c, 16'h6e1d, 16'h6e1e, 16'h6e1f 	:	val_out <= 16'hb675;
         16'h6e20, 16'h6e21, 16'h6e22, 16'h6e23, 16'h6e24, 16'h6e25, 16'h6e26, 16'h6e27 	:	val_out <= 16'hb65f;
         16'h6e28, 16'h6e29, 16'h6e2a, 16'h6e2b, 16'h6e2c, 16'h6e2d, 16'h6e2e, 16'h6e2f 	:	val_out <= 16'hb648;
         16'h6e30, 16'h6e31, 16'h6e32, 16'h6e33, 16'h6e34, 16'h6e35, 16'h6e36, 16'h6e37 	:	val_out <= 16'hb631;
         16'h6e38, 16'h6e39, 16'h6e3a, 16'h6e3b, 16'h6e3c, 16'h6e3d, 16'h6e3e, 16'h6e3f 	:	val_out <= 16'hb61a;
         16'h6e40, 16'h6e41, 16'h6e42, 16'h6e43, 16'h6e44, 16'h6e45, 16'h6e46, 16'h6e47 	:	val_out <= 16'hb604;
         16'h6e48, 16'h6e49, 16'h6e4a, 16'h6e4b, 16'h6e4c, 16'h6e4d, 16'h6e4e, 16'h6e4f 	:	val_out <= 16'hb5ed;
         16'h6e50, 16'h6e51, 16'h6e52, 16'h6e53, 16'h6e54, 16'h6e55, 16'h6e56, 16'h6e57 	:	val_out <= 16'hb5d6;
         16'h6e58, 16'h6e59, 16'h6e5a, 16'h6e5b, 16'h6e5c, 16'h6e5d, 16'h6e5e, 16'h6e5f 	:	val_out <= 16'hb5bf;
         16'h6e60, 16'h6e61, 16'h6e62, 16'h6e63, 16'h6e64, 16'h6e65, 16'h6e66, 16'h6e67 	:	val_out <= 16'hb5a8;
         16'h6e68, 16'h6e69, 16'h6e6a, 16'h6e6b, 16'h6e6c, 16'h6e6d, 16'h6e6e, 16'h6e6f 	:	val_out <= 16'hb592;
         16'h6e70, 16'h6e71, 16'h6e72, 16'h6e73, 16'h6e74, 16'h6e75, 16'h6e76, 16'h6e77 	:	val_out <= 16'hb57b;
         16'h6e78, 16'h6e79, 16'h6e7a, 16'h6e7b, 16'h6e7c, 16'h6e7d, 16'h6e7e, 16'h6e7f 	:	val_out <= 16'hb564;
         16'h6e80, 16'h6e81, 16'h6e82, 16'h6e83, 16'h6e84, 16'h6e85, 16'h6e86, 16'h6e87 	:	val_out <= 16'hb54d;
         16'h6e88, 16'h6e89, 16'h6e8a, 16'h6e8b, 16'h6e8c, 16'h6e8d, 16'h6e8e, 16'h6e8f 	:	val_out <= 16'hb536;
         16'h6e90, 16'h6e91, 16'h6e92, 16'h6e93, 16'h6e94, 16'h6e95, 16'h6e96, 16'h6e97 	:	val_out <= 16'hb51f;
         16'h6e98, 16'h6e99, 16'h6e9a, 16'h6e9b, 16'h6e9c, 16'h6e9d, 16'h6e9e, 16'h6e9f 	:	val_out <= 16'hb508;
         16'h6ea0, 16'h6ea1, 16'h6ea2, 16'h6ea3, 16'h6ea4, 16'h6ea5, 16'h6ea6, 16'h6ea7 	:	val_out <= 16'hb4f2;
         16'h6ea8, 16'h6ea9, 16'h6eaa, 16'h6eab, 16'h6eac, 16'h6ead, 16'h6eae, 16'h6eaf 	:	val_out <= 16'hb4db;
         16'h6eb0, 16'h6eb1, 16'h6eb2, 16'h6eb3, 16'h6eb4, 16'h6eb5, 16'h6eb6, 16'h6eb7 	:	val_out <= 16'hb4c4;
         16'h6eb8, 16'h6eb9, 16'h6eba, 16'h6ebb, 16'h6ebc, 16'h6ebd, 16'h6ebe, 16'h6ebf 	:	val_out <= 16'hb4ad;
         16'h6ec0, 16'h6ec1, 16'h6ec2, 16'h6ec3, 16'h6ec4, 16'h6ec5, 16'h6ec6, 16'h6ec7 	:	val_out <= 16'hb496;
         16'h6ec8, 16'h6ec9, 16'h6eca, 16'h6ecb, 16'h6ecc, 16'h6ecd, 16'h6ece, 16'h6ecf 	:	val_out <= 16'hb47f;
         16'h6ed0, 16'h6ed1, 16'h6ed2, 16'h6ed3, 16'h6ed4, 16'h6ed5, 16'h6ed6, 16'h6ed7 	:	val_out <= 16'hb468;
         16'h6ed8, 16'h6ed9, 16'h6eda, 16'h6edb, 16'h6edc, 16'h6edd, 16'h6ede, 16'h6edf 	:	val_out <= 16'hb451;
         16'h6ee0, 16'h6ee1, 16'h6ee2, 16'h6ee3, 16'h6ee4, 16'h6ee5, 16'h6ee6, 16'h6ee7 	:	val_out <= 16'hb43a;
         16'h6ee8, 16'h6ee9, 16'h6eea, 16'h6eeb, 16'h6eec, 16'h6eed, 16'h6eee, 16'h6eef 	:	val_out <= 16'hb423;
         16'h6ef0, 16'h6ef1, 16'h6ef2, 16'h6ef3, 16'h6ef4, 16'h6ef5, 16'h6ef6, 16'h6ef7 	:	val_out <= 16'hb40c;
         16'h6ef8, 16'h6ef9, 16'h6efa, 16'h6efb, 16'h6efc, 16'h6efd, 16'h6efe, 16'h6eff 	:	val_out <= 16'hb3f5;
         16'h6f00, 16'h6f01, 16'h6f02, 16'h6f03, 16'h6f04, 16'h6f05, 16'h6f06, 16'h6f07 	:	val_out <= 16'hb3de;
         16'h6f08, 16'h6f09, 16'h6f0a, 16'h6f0b, 16'h6f0c, 16'h6f0d, 16'h6f0e, 16'h6f0f 	:	val_out <= 16'hb3c7;
         16'h6f10, 16'h6f11, 16'h6f12, 16'h6f13, 16'h6f14, 16'h6f15, 16'h6f16, 16'h6f17 	:	val_out <= 16'hb3b0;
         16'h6f18, 16'h6f19, 16'h6f1a, 16'h6f1b, 16'h6f1c, 16'h6f1d, 16'h6f1e, 16'h6f1f 	:	val_out <= 16'hb399;
         16'h6f20, 16'h6f21, 16'h6f22, 16'h6f23, 16'h6f24, 16'h6f25, 16'h6f26, 16'h6f27 	:	val_out <= 16'hb382;
         16'h6f28, 16'h6f29, 16'h6f2a, 16'h6f2b, 16'h6f2c, 16'h6f2d, 16'h6f2e, 16'h6f2f 	:	val_out <= 16'hb36b;
         16'h6f30, 16'h6f31, 16'h6f32, 16'h6f33, 16'h6f34, 16'h6f35, 16'h6f36, 16'h6f37 	:	val_out <= 16'hb354;
         16'h6f38, 16'h6f39, 16'h6f3a, 16'h6f3b, 16'h6f3c, 16'h6f3d, 16'h6f3e, 16'h6f3f 	:	val_out <= 16'hb33d;
         16'h6f40, 16'h6f41, 16'h6f42, 16'h6f43, 16'h6f44, 16'h6f45, 16'h6f46, 16'h6f47 	:	val_out <= 16'hb326;
         16'h6f48, 16'h6f49, 16'h6f4a, 16'h6f4b, 16'h6f4c, 16'h6f4d, 16'h6f4e, 16'h6f4f 	:	val_out <= 16'hb30f;
         16'h6f50, 16'h6f51, 16'h6f52, 16'h6f53, 16'h6f54, 16'h6f55, 16'h6f56, 16'h6f57 	:	val_out <= 16'hb2f8;
         16'h6f58, 16'h6f59, 16'h6f5a, 16'h6f5b, 16'h6f5c, 16'h6f5d, 16'h6f5e, 16'h6f5f 	:	val_out <= 16'hb2e1;
         16'h6f60, 16'h6f61, 16'h6f62, 16'h6f63, 16'h6f64, 16'h6f65, 16'h6f66, 16'h6f67 	:	val_out <= 16'hb2ca;
         16'h6f68, 16'h6f69, 16'h6f6a, 16'h6f6b, 16'h6f6c, 16'h6f6d, 16'h6f6e, 16'h6f6f 	:	val_out <= 16'hb2b3;
         16'h6f70, 16'h6f71, 16'h6f72, 16'h6f73, 16'h6f74, 16'h6f75, 16'h6f76, 16'h6f77 	:	val_out <= 16'hb29c;
         16'h6f78, 16'h6f79, 16'h6f7a, 16'h6f7b, 16'h6f7c, 16'h6f7d, 16'h6f7e, 16'h6f7f 	:	val_out <= 16'hb285;
         16'h6f80, 16'h6f81, 16'h6f82, 16'h6f83, 16'h6f84, 16'h6f85, 16'h6f86, 16'h6f87 	:	val_out <= 16'hb26e;
         16'h6f88, 16'h6f89, 16'h6f8a, 16'h6f8b, 16'h6f8c, 16'h6f8d, 16'h6f8e, 16'h6f8f 	:	val_out <= 16'hb257;
         16'h6f90, 16'h6f91, 16'h6f92, 16'h6f93, 16'h6f94, 16'h6f95, 16'h6f96, 16'h6f97 	:	val_out <= 16'hb240;
         16'h6f98, 16'h6f99, 16'h6f9a, 16'h6f9b, 16'h6f9c, 16'h6f9d, 16'h6f9e, 16'h6f9f 	:	val_out <= 16'hb228;
         16'h6fa0, 16'h6fa1, 16'h6fa2, 16'h6fa3, 16'h6fa4, 16'h6fa5, 16'h6fa6, 16'h6fa7 	:	val_out <= 16'hb211;
         16'h6fa8, 16'h6fa9, 16'h6faa, 16'h6fab, 16'h6fac, 16'h6fad, 16'h6fae, 16'h6faf 	:	val_out <= 16'hb1fa;
         16'h6fb0, 16'h6fb1, 16'h6fb2, 16'h6fb3, 16'h6fb4, 16'h6fb5, 16'h6fb6, 16'h6fb7 	:	val_out <= 16'hb1e3;
         16'h6fb8, 16'h6fb9, 16'h6fba, 16'h6fbb, 16'h6fbc, 16'h6fbd, 16'h6fbe, 16'h6fbf 	:	val_out <= 16'hb1cc;
         16'h6fc0, 16'h6fc1, 16'h6fc2, 16'h6fc3, 16'h6fc4, 16'h6fc5, 16'h6fc6, 16'h6fc7 	:	val_out <= 16'hb1b5;
         16'h6fc8, 16'h6fc9, 16'h6fca, 16'h6fcb, 16'h6fcc, 16'h6fcd, 16'h6fce, 16'h6fcf 	:	val_out <= 16'hb19e;
         16'h6fd0, 16'h6fd1, 16'h6fd2, 16'h6fd3, 16'h6fd4, 16'h6fd5, 16'h6fd6, 16'h6fd7 	:	val_out <= 16'hb186;
         16'h6fd8, 16'h6fd9, 16'h6fda, 16'h6fdb, 16'h6fdc, 16'h6fdd, 16'h6fde, 16'h6fdf 	:	val_out <= 16'hb16f;
         16'h6fe0, 16'h6fe1, 16'h6fe2, 16'h6fe3, 16'h6fe4, 16'h6fe5, 16'h6fe6, 16'h6fe7 	:	val_out <= 16'hb158;
         16'h6fe8, 16'h6fe9, 16'h6fea, 16'h6feb, 16'h6fec, 16'h6fed, 16'h6fee, 16'h6fef 	:	val_out <= 16'hb141;
         16'h6ff0, 16'h6ff1, 16'h6ff2, 16'h6ff3, 16'h6ff4, 16'h6ff5, 16'h6ff6, 16'h6ff7 	:	val_out <= 16'hb12a;
         16'h6ff8, 16'h6ff9, 16'h6ffa, 16'h6ffb, 16'h6ffc, 16'h6ffd, 16'h6ffe, 16'h6fff 	:	val_out <= 16'hb112;
         16'h7000, 16'h7001, 16'h7002, 16'h7003, 16'h7004, 16'h7005, 16'h7006, 16'h7007 	:	val_out <= 16'hb0fb;
         16'h7008, 16'h7009, 16'h700a, 16'h700b, 16'h700c, 16'h700d, 16'h700e, 16'h700f 	:	val_out <= 16'hb0e4;
         16'h7010, 16'h7011, 16'h7012, 16'h7013, 16'h7014, 16'h7015, 16'h7016, 16'h7017 	:	val_out <= 16'hb0cd;
         16'h7018, 16'h7019, 16'h701a, 16'h701b, 16'h701c, 16'h701d, 16'h701e, 16'h701f 	:	val_out <= 16'hb0b6;
         16'h7020, 16'h7021, 16'h7022, 16'h7023, 16'h7024, 16'h7025, 16'h7026, 16'h7027 	:	val_out <= 16'hb09e;
         16'h7028, 16'h7029, 16'h702a, 16'h702b, 16'h702c, 16'h702d, 16'h702e, 16'h702f 	:	val_out <= 16'hb087;
         16'h7030, 16'h7031, 16'h7032, 16'h7033, 16'h7034, 16'h7035, 16'h7036, 16'h7037 	:	val_out <= 16'hb070;
         16'h7038, 16'h7039, 16'h703a, 16'h703b, 16'h703c, 16'h703d, 16'h703e, 16'h703f 	:	val_out <= 16'hb059;
         16'h7040, 16'h7041, 16'h7042, 16'h7043, 16'h7044, 16'h7045, 16'h7046, 16'h7047 	:	val_out <= 16'hb041;
         16'h7048, 16'h7049, 16'h704a, 16'h704b, 16'h704c, 16'h704d, 16'h704e, 16'h704f 	:	val_out <= 16'hb02a;
         16'h7050, 16'h7051, 16'h7052, 16'h7053, 16'h7054, 16'h7055, 16'h7056, 16'h7057 	:	val_out <= 16'hb013;
         16'h7058, 16'h7059, 16'h705a, 16'h705b, 16'h705c, 16'h705d, 16'h705e, 16'h705f 	:	val_out <= 16'haffb;
         16'h7060, 16'h7061, 16'h7062, 16'h7063, 16'h7064, 16'h7065, 16'h7066, 16'h7067 	:	val_out <= 16'hafe4;
         16'h7068, 16'h7069, 16'h706a, 16'h706b, 16'h706c, 16'h706d, 16'h706e, 16'h706f 	:	val_out <= 16'hafcd;
         16'h7070, 16'h7071, 16'h7072, 16'h7073, 16'h7074, 16'h7075, 16'h7076, 16'h7077 	:	val_out <= 16'hafb5;
         16'h7078, 16'h7079, 16'h707a, 16'h707b, 16'h707c, 16'h707d, 16'h707e, 16'h707f 	:	val_out <= 16'haf9e;
         16'h7080, 16'h7081, 16'h7082, 16'h7083, 16'h7084, 16'h7085, 16'h7086, 16'h7087 	:	val_out <= 16'haf87;
         16'h7088, 16'h7089, 16'h708a, 16'h708b, 16'h708c, 16'h708d, 16'h708e, 16'h708f 	:	val_out <= 16'haf6f;
         16'h7090, 16'h7091, 16'h7092, 16'h7093, 16'h7094, 16'h7095, 16'h7096, 16'h7097 	:	val_out <= 16'haf58;
         16'h7098, 16'h7099, 16'h709a, 16'h709b, 16'h709c, 16'h709d, 16'h709e, 16'h709f 	:	val_out <= 16'haf41;
         16'h70a0, 16'h70a1, 16'h70a2, 16'h70a3, 16'h70a4, 16'h70a5, 16'h70a6, 16'h70a7 	:	val_out <= 16'haf29;
         16'h70a8, 16'h70a9, 16'h70aa, 16'h70ab, 16'h70ac, 16'h70ad, 16'h70ae, 16'h70af 	:	val_out <= 16'haf12;
         16'h70b0, 16'h70b1, 16'h70b2, 16'h70b3, 16'h70b4, 16'h70b5, 16'h70b6, 16'h70b7 	:	val_out <= 16'haefb;
         16'h70b8, 16'h70b9, 16'h70ba, 16'h70bb, 16'h70bc, 16'h70bd, 16'h70be, 16'h70bf 	:	val_out <= 16'haee3;
         16'h70c0, 16'h70c1, 16'h70c2, 16'h70c3, 16'h70c4, 16'h70c5, 16'h70c6, 16'h70c7 	:	val_out <= 16'haecc;
         16'h70c8, 16'h70c9, 16'h70ca, 16'h70cb, 16'h70cc, 16'h70cd, 16'h70ce, 16'h70cf 	:	val_out <= 16'haeb5;
         16'h70d0, 16'h70d1, 16'h70d2, 16'h70d3, 16'h70d4, 16'h70d5, 16'h70d6, 16'h70d7 	:	val_out <= 16'hae9d;
         16'h70d8, 16'h70d9, 16'h70da, 16'h70db, 16'h70dc, 16'h70dd, 16'h70de, 16'h70df 	:	val_out <= 16'hae86;
         16'h70e0, 16'h70e1, 16'h70e2, 16'h70e3, 16'h70e4, 16'h70e5, 16'h70e6, 16'h70e7 	:	val_out <= 16'hae6e;
         16'h70e8, 16'h70e9, 16'h70ea, 16'h70eb, 16'h70ec, 16'h70ed, 16'h70ee, 16'h70ef 	:	val_out <= 16'hae57;
         16'h70f0, 16'h70f1, 16'h70f2, 16'h70f3, 16'h70f4, 16'h70f5, 16'h70f6, 16'h70f7 	:	val_out <= 16'hae3f;
         16'h70f8, 16'h70f9, 16'h70fa, 16'h70fb, 16'h70fc, 16'h70fd, 16'h70fe, 16'h70ff 	:	val_out <= 16'hae28;
         16'h7100, 16'h7101, 16'h7102, 16'h7103, 16'h7104, 16'h7105, 16'h7106, 16'h7107 	:	val_out <= 16'hae11;
         16'h7108, 16'h7109, 16'h710a, 16'h710b, 16'h710c, 16'h710d, 16'h710e, 16'h710f 	:	val_out <= 16'hadf9;
         16'h7110, 16'h7111, 16'h7112, 16'h7113, 16'h7114, 16'h7115, 16'h7116, 16'h7117 	:	val_out <= 16'hade2;
         16'h7118, 16'h7119, 16'h711a, 16'h711b, 16'h711c, 16'h711d, 16'h711e, 16'h711f 	:	val_out <= 16'hadca;
         16'h7120, 16'h7121, 16'h7122, 16'h7123, 16'h7124, 16'h7125, 16'h7126, 16'h7127 	:	val_out <= 16'hadb3;
         16'h7128, 16'h7129, 16'h712a, 16'h712b, 16'h712c, 16'h712d, 16'h712e, 16'h712f 	:	val_out <= 16'had9b;
         16'h7130, 16'h7131, 16'h7132, 16'h7133, 16'h7134, 16'h7135, 16'h7136, 16'h7137 	:	val_out <= 16'had84;
         16'h7138, 16'h7139, 16'h713a, 16'h713b, 16'h713c, 16'h713d, 16'h713e, 16'h713f 	:	val_out <= 16'had6c;
         16'h7140, 16'h7141, 16'h7142, 16'h7143, 16'h7144, 16'h7145, 16'h7146, 16'h7147 	:	val_out <= 16'had55;
         16'h7148, 16'h7149, 16'h714a, 16'h714b, 16'h714c, 16'h714d, 16'h714e, 16'h714f 	:	val_out <= 16'had3d;
         16'h7150, 16'h7151, 16'h7152, 16'h7153, 16'h7154, 16'h7155, 16'h7156, 16'h7157 	:	val_out <= 16'had26;
         16'h7158, 16'h7159, 16'h715a, 16'h715b, 16'h715c, 16'h715d, 16'h715e, 16'h715f 	:	val_out <= 16'had0e;
         16'h7160, 16'h7161, 16'h7162, 16'h7163, 16'h7164, 16'h7165, 16'h7166, 16'h7167 	:	val_out <= 16'hacf7;
         16'h7168, 16'h7169, 16'h716a, 16'h716b, 16'h716c, 16'h716d, 16'h716e, 16'h716f 	:	val_out <= 16'hacdf;
         16'h7170, 16'h7171, 16'h7172, 16'h7173, 16'h7174, 16'h7175, 16'h7176, 16'h7177 	:	val_out <= 16'hacc8;
         16'h7178, 16'h7179, 16'h717a, 16'h717b, 16'h717c, 16'h717d, 16'h717e, 16'h717f 	:	val_out <= 16'hacb0;
         16'h7180, 16'h7181, 16'h7182, 16'h7183, 16'h7184, 16'h7185, 16'h7186, 16'h7187 	:	val_out <= 16'hac98;
         16'h7188, 16'h7189, 16'h718a, 16'h718b, 16'h718c, 16'h718d, 16'h718e, 16'h718f 	:	val_out <= 16'hac81;
         16'h7190, 16'h7191, 16'h7192, 16'h7193, 16'h7194, 16'h7195, 16'h7196, 16'h7197 	:	val_out <= 16'hac69;
         16'h7198, 16'h7199, 16'h719a, 16'h719b, 16'h719c, 16'h719d, 16'h719e, 16'h719f 	:	val_out <= 16'hac52;
         16'h71a0, 16'h71a1, 16'h71a2, 16'h71a3, 16'h71a4, 16'h71a5, 16'h71a6, 16'h71a7 	:	val_out <= 16'hac3a;
         16'h71a8, 16'h71a9, 16'h71aa, 16'h71ab, 16'h71ac, 16'h71ad, 16'h71ae, 16'h71af 	:	val_out <= 16'hac23;
         16'h71b0, 16'h71b1, 16'h71b2, 16'h71b3, 16'h71b4, 16'h71b5, 16'h71b6, 16'h71b7 	:	val_out <= 16'hac0b;
         16'h71b8, 16'h71b9, 16'h71ba, 16'h71bb, 16'h71bc, 16'h71bd, 16'h71be, 16'h71bf 	:	val_out <= 16'habf3;
         16'h71c0, 16'h71c1, 16'h71c2, 16'h71c3, 16'h71c4, 16'h71c5, 16'h71c6, 16'h71c7 	:	val_out <= 16'habdc;
         16'h71c8, 16'h71c9, 16'h71ca, 16'h71cb, 16'h71cc, 16'h71cd, 16'h71ce, 16'h71cf 	:	val_out <= 16'habc4;
         16'h71d0, 16'h71d1, 16'h71d2, 16'h71d3, 16'h71d4, 16'h71d5, 16'h71d6, 16'h71d7 	:	val_out <= 16'habad;
         16'h71d8, 16'h71d9, 16'h71da, 16'h71db, 16'h71dc, 16'h71dd, 16'h71de, 16'h71df 	:	val_out <= 16'hab95;
         16'h71e0, 16'h71e1, 16'h71e2, 16'h71e3, 16'h71e4, 16'h71e5, 16'h71e6, 16'h71e7 	:	val_out <= 16'hab7d;
         16'h71e8, 16'h71e9, 16'h71ea, 16'h71eb, 16'h71ec, 16'h71ed, 16'h71ee, 16'h71ef 	:	val_out <= 16'hab66;
         16'h71f0, 16'h71f1, 16'h71f2, 16'h71f3, 16'h71f4, 16'h71f5, 16'h71f6, 16'h71f7 	:	val_out <= 16'hab4e;
         16'h71f8, 16'h71f9, 16'h71fa, 16'h71fb, 16'h71fc, 16'h71fd, 16'h71fe, 16'h71ff 	:	val_out <= 16'hab36;
         16'h7200, 16'h7201, 16'h7202, 16'h7203, 16'h7204, 16'h7205, 16'h7206, 16'h7207 	:	val_out <= 16'hab1f;
         16'h7208, 16'h7209, 16'h720a, 16'h720b, 16'h720c, 16'h720d, 16'h720e, 16'h720f 	:	val_out <= 16'hab07;
         16'h7210, 16'h7211, 16'h7212, 16'h7213, 16'h7214, 16'h7215, 16'h7216, 16'h7217 	:	val_out <= 16'haaef;
         16'h7218, 16'h7219, 16'h721a, 16'h721b, 16'h721c, 16'h721d, 16'h721e, 16'h721f 	:	val_out <= 16'haad8;
         16'h7220, 16'h7221, 16'h7222, 16'h7223, 16'h7224, 16'h7225, 16'h7226, 16'h7227 	:	val_out <= 16'haac0;
         16'h7228, 16'h7229, 16'h722a, 16'h722b, 16'h722c, 16'h722d, 16'h722e, 16'h722f 	:	val_out <= 16'haaa8;
         16'h7230, 16'h7231, 16'h7232, 16'h7233, 16'h7234, 16'h7235, 16'h7236, 16'h7237 	:	val_out <= 16'haa91;
         16'h7238, 16'h7239, 16'h723a, 16'h723b, 16'h723c, 16'h723d, 16'h723e, 16'h723f 	:	val_out <= 16'haa79;
         16'h7240, 16'h7241, 16'h7242, 16'h7243, 16'h7244, 16'h7245, 16'h7246, 16'h7247 	:	val_out <= 16'haa61;
         16'h7248, 16'h7249, 16'h724a, 16'h724b, 16'h724c, 16'h724d, 16'h724e, 16'h724f 	:	val_out <= 16'haa49;
         16'h7250, 16'h7251, 16'h7252, 16'h7253, 16'h7254, 16'h7255, 16'h7256, 16'h7257 	:	val_out <= 16'haa32;
         16'h7258, 16'h7259, 16'h725a, 16'h725b, 16'h725c, 16'h725d, 16'h725e, 16'h725f 	:	val_out <= 16'haa1a;
         16'h7260, 16'h7261, 16'h7262, 16'h7263, 16'h7264, 16'h7265, 16'h7266, 16'h7267 	:	val_out <= 16'haa02;
         16'h7268, 16'h7269, 16'h726a, 16'h726b, 16'h726c, 16'h726d, 16'h726e, 16'h726f 	:	val_out <= 16'ha9eb;
         16'h7270, 16'h7271, 16'h7272, 16'h7273, 16'h7274, 16'h7275, 16'h7276, 16'h7277 	:	val_out <= 16'ha9d3;
         16'h7278, 16'h7279, 16'h727a, 16'h727b, 16'h727c, 16'h727d, 16'h727e, 16'h727f 	:	val_out <= 16'ha9bb;
         16'h7280, 16'h7281, 16'h7282, 16'h7283, 16'h7284, 16'h7285, 16'h7286, 16'h7287 	:	val_out <= 16'ha9a3;
         16'h7288, 16'h7289, 16'h728a, 16'h728b, 16'h728c, 16'h728d, 16'h728e, 16'h728f 	:	val_out <= 16'ha98b;
         16'h7290, 16'h7291, 16'h7292, 16'h7293, 16'h7294, 16'h7295, 16'h7296, 16'h7297 	:	val_out <= 16'ha974;
         16'h7298, 16'h7299, 16'h729a, 16'h729b, 16'h729c, 16'h729d, 16'h729e, 16'h729f 	:	val_out <= 16'ha95c;
         16'h72a0, 16'h72a1, 16'h72a2, 16'h72a3, 16'h72a4, 16'h72a5, 16'h72a6, 16'h72a7 	:	val_out <= 16'ha944;
         16'h72a8, 16'h72a9, 16'h72aa, 16'h72ab, 16'h72ac, 16'h72ad, 16'h72ae, 16'h72af 	:	val_out <= 16'ha92c;
         16'h72b0, 16'h72b1, 16'h72b2, 16'h72b3, 16'h72b4, 16'h72b5, 16'h72b6, 16'h72b7 	:	val_out <= 16'ha915;
         16'h72b8, 16'h72b9, 16'h72ba, 16'h72bb, 16'h72bc, 16'h72bd, 16'h72be, 16'h72bf 	:	val_out <= 16'ha8fd;
         16'h72c0, 16'h72c1, 16'h72c2, 16'h72c3, 16'h72c4, 16'h72c5, 16'h72c6, 16'h72c7 	:	val_out <= 16'ha8e5;
         16'h72c8, 16'h72c9, 16'h72ca, 16'h72cb, 16'h72cc, 16'h72cd, 16'h72ce, 16'h72cf 	:	val_out <= 16'ha8cd;
         16'h72d0, 16'h72d1, 16'h72d2, 16'h72d3, 16'h72d4, 16'h72d5, 16'h72d6, 16'h72d7 	:	val_out <= 16'ha8b5;
         16'h72d8, 16'h72d9, 16'h72da, 16'h72db, 16'h72dc, 16'h72dd, 16'h72de, 16'h72df 	:	val_out <= 16'ha89d;
         16'h72e0, 16'h72e1, 16'h72e2, 16'h72e3, 16'h72e4, 16'h72e5, 16'h72e6, 16'h72e7 	:	val_out <= 16'ha886;
         16'h72e8, 16'h72e9, 16'h72ea, 16'h72eb, 16'h72ec, 16'h72ed, 16'h72ee, 16'h72ef 	:	val_out <= 16'ha86e;
         16'h72f0, 16'h72f1, 16'h72f2, 16'h72f3, 16'h72f4, 16'h72f5, 16'h72f6, 16'h72f7 	:	val_out <= 16'ha856;
         16'h72f8, 16'h72f9, 16'h72fa, 16'h72fb, 16'h72fc, 16'h72fd, 16'h72fe, 16'h72ff 	:	val_out <= 16'ha83e;
         16'h7300, 16'h7301, 16'h7302, 16'h7303, 16'h7304, 16'h7305, 16'h7306, 16'h7307 	:	val_out <= 16'ha826;
         16'h7308, 16'h7309, 16'h730a, 16'h730b, 16'h730c, 16'h730d, 16'h730e, 16'h730f 	:	val_out <= 16'ha80e;
         16'h7310, 16'h7311, 16'h7312, 16'h7313, 16'h7314, 16'h7315, 16'h7316, 16'h7317 	:	val_out <= 16'ha7f6;
         16'h7318, 16'h7319, 16'h731a, 16'h731b, 16'h731c, 16'h731d, 16'h731e, 16'h731f 	:	val_out <= 16'ha7df;
         16'h7320, 16'h7321, 16'h7322, 16'h7323, 16'h7324, 16'h7325, 16'h7326, 16'h7327 	:	val_out <= 16'ha7c7;
         16'h7328, 16'h7329, 16'h732a, 16'h732b, 16'h732c, 16'h732d, 16'h732e, 16'h732f 	:	val_out <= 16'ha7af;
         16'h7330, 16'h7331, 16'h7332, 16'h7333, 16'h7334, 16'h7335, 16'h7336, 16'h7337 	:	val_out <= 16'ha797;
         16'h7338, 16'h7339, 16'h733a, 16'h733b, 16'h733c, 16'h733d, 16'h733e, 16'h733f 	:	val_out <= 16'ha77f;
         16'h7340, 16'h7341, 16'h7342, 16'h7343, 16'h7344, 16'h7345, 16'h7346, 16'h7347 	:	val_out <= 16'ha767;
         16'h7348, 16'h7349, 16'h734a, 16'h734b, 16'h734c, 16'h734d, 16'h734e, 16'h734f 	:	val_out <= 16'ha74f;
         16'h7350, 16'h7351, 16'h7352, 16'h7353, 16'h7354, 16'h7355, 16'h7356, 16'h7357 	:	val_out <= 16'ha737;
         16'h7358, 16'h7359, 16'h735a, 16'h735b, 16'h735c, 16'h735d, 16'h735e, 16'h735f 	:	val_out <= 16'ha71f;
         16'h7360, 16'h7361, 16'h7362, 16'h7363, 16'h7364, 16'h7365, 16'h7366, 16'h7367 	:	val_out <= 16'ha707;
         16'h7368, 16'h7369, 16'h736a, 16'h736b, 16'h736c, 16'h736d, 16'h736e, 16'h736f 	:	val_out <= 16'ha6ef;
         16'h7370, 16'h7371, 16'h7372, 16'h7373, 16'h7374, 16'h7375, 16'h7376, 16'h7377 	:	val_out <= 16'ha6d8;
         16'h7378, 16'h7379, 16'h737a, 16'h737b, 16'h737c, 16'h737d, 16'h737e, 16'h737f 	:	val_out <= 16'ha6c0;
         16'h7380, 16'h7381, 16'h7382, 16'h7383, 16'h7384, 16'h7385, 16'h7386, 16'h7387 	:	val_out <= 16'ha6a8;
         16'h7388, 16'h7389, 16'h738a, 16'h738b, 16'h738c, 16'h738d, 16'h738e, 16'h738f 	:	val_out <= 16'ha690;
         16'h7390, 16'h7391, 16'h7392, 16'h7393, 16'h7394, 16'h7395, 16'h7396, 16'h7397 	:	val_out <= 16'ha678;
         16'h7398, 16'h7399, 16'h739a, 16'h739b, 16'h739c, 16'h739d, 16'h739e, 16'h739f 	:	val_out <= 16'ha660;
         16'h73a0, 16'h73a1, 16'h73a2, 16'h73a3, 16'h73a4, 16'h73a5, 16'h73a6, 16'h73a7 	:	val_out <= 16'ha648;
         16'h73a8, 16'h73a9, 16'h73aa, 16'h73ab, 16'h73ac, 16'h73ad, 16'h73ae, 16'h73af 	:	val_out <= 16'ha630;
         16'h73b0, 16'h73b1, 16'h73b2, 16'h73b3, 16'h73b4, 16'h73b5, 16'h73b6, 16'h73b7 	:	val_out <= 16'ha618;
         16'h73b8, 16'h73b9, 16'h73ba, 16'h73bb, 16'h73bc, 16'h73bd, 16'h73be, 16'h73bf 	:	val_out <= 16'ha600;
         16'h73c0, 16'h73c1, 16'h73c2, 16'h73c3, 16'h73c4, 16'h73c5, 16'h73c6, 16'h73c7 	:	val_out <= 16'ha5e8;
         16'h73c8, 16'h73c9, 16'h73ca, 16'h73cb, 16'h73cc, 16'h73cd, 16'h73ce, 16'h73cf 	:	val_out <= 16'ha5d0;
         16'h73d0, 16'h73d1, 16'h73d2, 16'h73d3, 16'h73d4, 16'h73d5, 16'h73d6, 16'h73d7 	:	val_out <= 16'ha5b8;
         16'h73d8, 16'h73d9, 16'h73da, 16'h73db, 16'h73dc, 16'h73dd, 16'h73de, 16'h73df 	:	val_out <= 16'ha5a0;
         16'h73e0, 16'h73e1, 16'h73e2, 16'h73e3, 16'h73e4, 16'h73e5, 16'h73e6, 16'h73e7 	:	val_out <= 16'ha588;
         16'h73e8, 16'h73e9, 16'h73ea, 16'h73eb, 16'h73ec, 16'h73ed, 16'h73ee, 16'h73ef 	:	val_out <= 16'ha570;
         16'h73f0, 16'h73f1, 16'h73f2, 16'h73f3, 16'h73f4, 16'h73f5, 16'h73f6, 16'h73f7 	:	val_out <= 16'ha558;
         16'h73f8, 16'h73f9, 16'h73fa, 16'h73fb, 16'h73fc, 16'h73fd, 16'h73fe, 16'h73ff 	:	val_out <= 16'ha540;
         16'h7400, 16'h7401, 16'h7402, 16'h7403, 16'h7404, 16'h7405, 16'h7406, 16'h7407 	:	val_out <= 16'ha528;
         16'h7408, 16'h7409, 16'h740a, 16'h740b, 16'h740c, 16'h740d, 16'h740e, 16'h740f 	:	val_out <= 16'ha50f;
         16'h7410, 16'h7411, 16'h7412, 16'h7413, 16'h7414, 16'h7415, 16'h7416, 16'h7417 	:	val_out <= 16'ha4f7;
         16'h7418, 16'h7419, 16'h741a, 16'h741b, 16'h741c, 16'h741d, 16'h741e, 16'h741f 	:	val_out <= 16'ha4df;
         16'h7420, 16'h7421, 16'h7422, 16'h7423, 16'h7424, 16'h7425, 16'h7426, 16'h7427 	:	val_out <= 16'ha4c7;
         16'h7428, 16'h7429, 16'h742a, 16'h742b, 16'h742c, 16'h742d, 16'h742e, 16'h742f 	:	val_out <= 16'ha4af;
         16'h7430, 16'h7431, 16'h7432, 16'h7433, 16'h7434, 16'h7435, 16'h7436, 16'h7437 	:	val_out <= 16'ha497;
         16'h7438, 16'h7439, 16'h743a, 16'h743b, 16'h743c, 16'h743d, 16'h743e, 16'h743f 	:	val_out <= 16'ha47f;
         16'h7440, 16'h7441, 16'h7442, 16'h7443, 16'h7444, 16'h7445, 16'h7446, 16'h7447 	:	val_out <= 16'ha467;
         16'h7448, 16'h7449, 16'h744a, 16'h744b, 16'h744c, 16'h744d, 16'h744e, 16'h744f 	:	val_out <= 16'ha44f;
         16'h7450, 16'h7451, 16'h7452, 16'h7453, 16'h7454, 16'h7455, 16'h7456, 16'h7457 	:	val_out <= 16'ha437;
         16'h7458, 16'h7459, 16'h745a, 16'h745b, 16'h745c, 16'h745d, 16'h745e, 16'h745f 	:	val_out <= 16'ha41f;
         16'h7460, 16'h7461, 16'h7462, 16'h7463, 16'h7464, 16'h7465, 16'h7466, 16'h7467 	:	val_out <= 16'ha407;
         16'h7468, 16'h7469, 16'h746a, 16'h746b, 16'h746c, 16'h746d, 16'h746e, 16'h746f 	:	val_out <= 16'ha3ee;
         16'h7470, 16'h7471, 16'h7472, 16'h7473, 16'h7474, 16'h7475, 16'h7476, 16'h7477 	:	val_out <= 16'ha3d6;
         16'h7478, 16'h7479, 16'h747a, 16'h747b, 16'h747c, 16'h747d, 16'h747e, 16'h747f 	:	val_out <= 16'ha3be;
         16'h7480, 16'h7481, 16'h7482, 16'h7483, 16'h7484, 16'h7485, 16'h7486, 16'h7487 	:	val_out <= 16'ha3a6;
         16'h7488, 16'h7489, 16'h748a, 16'h748b, 16'h748c, 16'h748d, 16'h748e, 16'h748f 	:	val_out <= 16'ha38e;
         16'h7490, 16'h7491, 16'h7492, 16'h7493, 16'h7494, 16'h7495, 16'h7496, 16'h7497 	:	val_out <= 16'ha376;
         16'h7498, 16'h7499, 16'h749a, 16'h749b, 16'h749c, 16'h749d, 16'h749e, 16'h749f 	:	val_out <= 16'ha35e;
         16'h74a0, 16'h74a1, 16'h74a2, 16'h74a3, 16'h74a4, 16'h74a5, 16'h74a6, 16'h74a7 	:	val_out <= 16'ha345;
         16'h74a8, 16'h74a9, 16'h74aa, 16'h74ab, 16'h74ac, 16'h74ad, 16'h74ae, 16'h74af 	:	val_out <= 16'ha32d;
         16'h74b0, 16'h74b1, 16'h74b2, 16'h74b3, 16'h74b4, 16'h74b5, 16'h74b6, 16'h74b7 	:	val_out <= 16'ha315;
         16'h74b8, 16'h74b9, 16'h74ba, 16'h74bb, 16'h74bc, 16'h74bd, 16'h74be, 16'h74bf 	:	val_out <= 16'ha2fd;
         16'h74c0, 16'h74c1, 16'h74c2, 16'h74c3, 16'h74c4, 16'h74c5, 16'h74c6, 16'h74c7 	:	val_out <= 16'ha2e5;
         16'h74c8, 16'h74c9, 16'h74ca, 16'h74cb, 16'h74cc, 16'h74cd, 16'h74ce, 16'h74cf 	:	val_out <= 16'ha2cd;
         16'h74d0, 16'h74d1, 16'h74d2, 16'h74d3, 16'h74d4, 16'h74d5, 16'h74d6, 16'h74d7 	:	val_out <= 16'ha2b4;
         16'h74d8, 16'h74d9, 16'h74da, 16'h74db, 16'h74dc, 16'h74dd, 16'h74de, 16'h74df 	:	val_out <= 16'ha29c;
         16'h74e0, 16'h74e1, 16'h74e2, 16'h74e3, 16'h74e4, 16'h74e5, 16'h74e6, 16'h74e7 	:	val_out <= 16'ha284;
         16'h74e8, 16'h74e9, 16'h74ea, 16'h74eb, 16'h74ec, 16'h74ed, 16'h74ee, 16'h74ef 	:	val_out <= 16'ha26c;
         16'h74f0, 16'h74f1, 16'h74f2, 16'h74f3, 16'h74f4, 16'h74f5, 16'h74f6, 16'h74f7 	:	val_out <= 16'ha254;
         16'h74f8, 16'h74f9, 16'h74fa, 16'h74fb, 16'h74fc, 16'h74fd, 16'h74fe, 16'h74ff 	:	val_out <= 16'ha23b;
         16'h7500, 16'h7501, 16'h7502, 16'h7503, 16'h7504, 16'h7505, 16'h7506, 16'h7507 	:	val_out <= 16'ha223;
         16'h7508, 16'h7509, 16'h750a, 16'h750b, 16'h750c, 16'h750d, 16'h750e, 16'h750f 	:	val_out <= 16'ha20b;
         16'h7510, 16'h7511, 16'h7512, 16'h7513, 16'h7514, 16'h7515, 16'h7516, 16'h7517 	:	val_out <= 16'ha1f3;
         16'h7518, 16'h7519, 16'h751a, 16'h751b, 16'h751c, 16'h751d, 16'h751e, 16'h751f 	:	val_out <= 16'ha1da;
         16'h7520, 16'h7521, 16'h7522, 16'h7523, 16'h7524, 16'h7525, 16'h7526, 16'h7527 	:	val_out <= 16'ha1c2;
         16'h7528, 16'h7529, 16'h752a, 16'h752b, 16'h752c, 16'h752d, 16'h752e, 16'h752f 	:	val_out <= 16'ha1aa;
         16'h7530, 16'h7531, 16'h7532, 16'h7533, 16'h7534, 16'h7535, 16'h7536, 16'h7537 	:	val_out <= 16'ha192;
         16'h7538, 16'h7539, 16'h753a, 16'h753b, 16'h753c, 16'h753d, 16'h753e, 16'h753f 	:	val_out <= 16'ha179;
         16'h7540, 16'h7541, 16'h7542, 16'h7543, 16'h7544, 16'h7545, 16'h7546, 16'h7547 	:	val_out <= 16'ha161;
         16'h7548, 16'h7549, 16'h754a, 16'h754b, 16'h754c, 16'h754d, 16'h754e, 16'h754f 	:	val_out <= 16'ha149;
         16'h7550, 16'h7551, 16'h7552, 16'h7553, 16'h7554, 16'h7555, 16'h7556, 16'h7557 	:	val_out <= 16'ha131;
         16'h7558, 16'h7559, 16'h755a, 16'h755b, 16'h755c, 16'h755d, 16'h755e, 16'h755f 	:	val_out <= 16'ha118;
         16'h7560, 16'h7561, 16'h7562, 16'h7563, 16'h7564, 16'h7565, 16'h7566, 16'h7567 	:	val_out <= 16'ha100;
         16'h7568, 16'h7569, 16'h756a, 16'h756b, 16'h756c, 16'h756d, 16'h756e, 16'h756f 	:	val_out <= 16'ha0e8;
         16'h7570, 16'h7571, 16'h7572, 16'h7573, 16'h7574, 16'h7575, 16'h7576, 16'h7577 	:	val_out <= 16'ha0d0;
         16'h7578, 16'h7579, 16'h757a, 16'h757b, 16'h757c, 16'h757d, 16'h757e, 16'h757f 	:	val_out <= 16'ha0b7;
         16'h7580, 16'h7581, 16'h7582, 16'h7583, 16'h7584, 16'h7585, 16'h7586, 16'h7587 	:	val_out <= 16'ha09f;
         16'h7588, 16'h7589, 16'h758a, 16'h758b, 16'h758c, 16'h758d, 16'h758e, 16'h758f 	:	val_out <= 16'ha087;
         16'h7590, 16'h7591, 16'h7592, 16'h7593, 16'h7594, 16'h7595, 16'h7596, 16'h7597 	:	val_out <= 16'ha06e;
         16'h7598, 16'h7599, 16'h759a, 16'h759b, 16'h759c, 16'h759d, 16'h759e, 16'h759f 	:	val_out <= 16'ha056;
         16'h75a0, 16'h75a1, 16'h75a2, 16'h75a3, 16'h75a4, 16'h75a5, 16'h75a6, 16'h75a7 	:	val_out <= 16'ha03e;
         16'h75a8, 16'h75a9, 16'h75aa, 16'h75ab, 16'h75ac, 16'h75ad, 16'h75ae, 16'h75af 	:	val_out <= 16'ha025;
         16'h75b0, 16'h75b1, 16'h75b2, 16'h75b3, 16'h75b4, 16'h75b5, 16'h75b6, 16'h75b7 	:	val_out <= 16'ha00d;
         16'h75b8, 16'h75b9, 16'h75ba, 16'h75bb, 16'h75bc, 16'h75bd, 16'h75be, 16'h75bf 	:	val_out <= 16'h9ff5;
         16'h75c0, 16'h75c1, 16'h75c2, 16'h75c3, 16'h75c4, 16'h75c5, 16'h75c6, 16'h75c7 	:	val_out <= 16'h9fdc;
         16'h75c8, 16'h75c9, 16'h75ca, 16'h75cb, 16'h75cc, 16'h75cd, 16'h75ce, 16'h75cf 	:	val_out <= 16'h9fc4;
         16'h75d0, 16'h75d1, 16'h75d2, 16'h75d3, 16'h75d4, 16'h75d5, 16'h75d6, 16'h75d7 	:	val_out <= 16'h9fac;
         16'h75d8, 16'h75d9, 16'h75da, 16'h75db, 16'h75dc, 16'h75dd, 16'h75de, 16'h75df 	:	val_out <= 16'h9f93;
         16'h75e0, 16'h75e1, 16'h75e2, 16'h75e3, 16'h75e4, 16'h75e5, 16'h75e6, 16'h75e7 	:	val_out <= 16'h9f7b;
         16'h75e8, 16'h75e9, 16'h75ea, 16'h75eb, 16'h75ec, 16'h75ed, 16'h75ee, 16'h75ef 	:	val_out <= 16'h9f63;
         16'h75f0, 16'h75f1, 16'h75f2, 16'h75f3, 16'h75f4, 16'h75f5, 16'h75f6, 16'h75f7 	:	val_out <= 16'h9f4a;
         16'h75f8, 16'h75f9, 16'h75fa, 16'h75fb, 16'h75fc, 16'h75fd, 16'h75fe, 16'h75ff 	:	val_out <= 16'h9f32;
         16'h7600, 16'h7601, 16'h7602, 16'h7603, 16'h7604, 16'h7605, 16'h7606, 16'h7607 	:	val_out <= 16'h9f19;
         16'h7608, 16'h7609, 16'h760a, 16'h760b, 16'h760c, 16'h760d, 16'h760e, 16'h760f 	:	val_out <= 16'h9f01;
         16'h7610, 16'h7611, 16'h7612, 16'h7613, 16'h7614, 16'h7615, 16'h7616, 16'h7617 	:	val_out <= 16'h9ee9;
         16'h7618, 16'h7619, 16'h761a, 16'h761b, 16'h761c, 16'h761d, 16'h761e, 16'h761f 	:	val_out <= 16'h9ed0;
         16'h7620, 16'h7621, 16'h7622, 16'h7623, 16'h7624, 16'h7625, 16'h7626, 16'h7627 	:	val_out <= 16'h9eb8;
         16'h7628, 16'h7629, 16'h762a, 16'h762b, 16'h762c, 16'h762d, 16'h762e, 16'h762f 	:	val_out <= 16'h9ea0;
         16'h7630, 16'h7631, 16'h7632, 16'h7633, 16'h7634, 16'h7635, 16'h7636, 16'h7637 	:	val_out <= 16'h9e87;
         16'h7638, 16'h7639, 16'h763a, 16'h763b, 16'h763c, 16'h763d, 16'h763e, 16'h763f 	:	val_out <= 16'h9e6f;
         16'h7640, 16'h7641, 16'h7642, 16'h7643, 16'h7644, 16'h7645, 16'h7646, 16'h7647 	:	val_out <= 16'h9e56;
         16'h7648, 16'h7649, 16'h764a, 16'h764b, 16'h764c, 16'h764d, 16'h764e, 16'h764f 	:	val_out <= 16'h9e3e;
         16'h7650, 16'h7651, 16'h7652, 16'h7653, 16'h7654, 16'h7655, 16'h7656, 16'h7657 	:	val_out <= 16'h9e25;
         16'h7658, 16'h7659, 16'h765a, 16'h765b, 16'h765c, 16'h765d, 16'h765e, 16'h765f 	:	val_out <= 16'h9e0d;
         16'h7660, 16'h7661, 16'h7662, 16'h7663, 16'h7664, 16'h7665, 16'h7666, 16'h7667 	:	val_out <= 16'h9df5;
         16'h7668, 16'h7669, 16'h766a, 16'h766b, 16'h766c, 16'h766d, 16'h766e, 16'h766f 	:	val_out <= 16'h9ddc;
         16'h7670, 16'h7671, 16'h7672, 16'h7673, 16'h7674, 16'h7675, 16'h7676, 16'h7677 	:	val_out <= 16'h9dc4;
         16'h7678, 16'h7679, 16'h767a, 16'h767b, 16'h767c, 16'h767d, 16'h767e, 16'h767f 	:	val_out <= 16'h9dab;
         16'h7680, 16'h7681, 16'h7682, 16'h7683, 16'h7684, 16'h7685, 16'h7686, 16'h7687 	:	val_out <= 16'h9d93;
         16'h7688, 16'h7689, 16'h768a, 16'h768b, 16'h768c, 16'h768d, 16'h768e, 16'h768f 	:	val_out <= 16'h9d7a;
         16'h7690, 16'h7691, 16'h7692, 16'h7693, 16'h7694, 16'h7695, 16'h7696, 16'h7697 	:	val_out <= 16'h9d62;
         16'h7698, 16'h7699, 16'h769a, 16'h769b, 16'h769c, 16'h769d, 16'h769e, 16'h769f 	:	val_out <= 16'h9d49;
         16'h76a0, 16'h76a1, 16'h76a2, 16'h76a3, 16'h76a4, 16'h76a5, 16'h76a6, 16'h76a7 	:	val_out <= 16'h9d31;
         16'h76a8, 16'h76a9, 16'h76aa, 16'h76ab, 16'h76ac, 16'h76ad, 16'h76ae, 16'h76af 	:	val_out <= 16'h9d18;
         16'h76b0, 16'h76b1, 16'h76b2, 16'h76b3, 16'h76b4, 16'h76b5, 16'h76b6, 16'h76b7 	:	val_out <= 16'h9d00;
         16'h76b8, 16'h76b9, 16'h76ba, 16'h76bb, 16'h76bc, 16'h76bd, 16'h76be, 16'h76bf 	:	val_out <= 16'h9ce8;
         16'h76c0, 16'h76c1, 16'h76c2, 16'h76c3, 16'h76c4, 16'h76c5, 16'h76c6, 16'h76c7 	:	val_out <= 16'h9ccf;
         16'h76c8, 16'h76c9, 16'h76ca, 16'h76cb, 16'h76cc, 16'h76cd, 16'h76ce, 16'h76cf 	:	val_out <= 16'h9cb7;
         16'h76d0, 16'h76d1, 16'h76d2, 16'h76d3, 16'h76d4, 16'h76d5, 16'h76d6, 16'h76d7 	:	val_out <= 16'h9c9e;
         16'h76d8, 16'h76d9, 16'h76da, 16'h76db, 16'h76dc, 16'h76dd, 16'h76de, 16'h76df 	:	val_out <= 16'h9c86;
         16'h76e0, 16'h76e1, 16'h76e2, 16'h76e3, 16'h76e4, 16'h76e5, 16'h76e6, 16'h76e7 	:	val_out <= 16'h9c6d;
         16'h76e8, 16'h76e9, 16'h76ea, 16'h76eb, 16'h76ec, 16'h76ed, 16'h76ee, 16'h76ef 	:	val_out <= 16'h9c55;
         16'h76f0, 16'h76f1, 16'h76f2, 16'h76f3, 16'h76f4, 16'h76f5, 16'h76f6, 16'h76f7 	:	val_out <= 16'h9c3c;
         16'h76f8, 16'h76f9, 16'h76fa, 16'h76fb, 16'h76fc, 16'h76fd, 16'h76fe, 16'h76ff 	:	val_out <= 16'h9c24;
         16'h7700, 16'h7701, 16'h7702, 16'h7703, 16'h7704, 16'h7705, 16'h7706, 16'h7707 	:	val_out <= 16'h9c0b;
         16'h7708, 16'h7709, 16'h770a, 16'h770b, 16'h770c, 16'h770d, 16'h770e, 16'h770f 	:	val_out <= 16'h9bf2;
         16'h7710, 16'h7711, 16'h7712, 16'h7713, 16'h7714, 16'h7715, 16'h7716, 16'h7717 	:	val_out <= 16'h9bda;
         16'h7718, 16'h7719, 16'h771a, 16'h771b, 16'h771c, 16'h771d, 16'h771e, 16'h771f 	:	val_out <= 16'h9bc1;
         16'h7720, 16'h7721, 16'h7722, 16'h7723, 16'h7724, 16'h7725, 16'h7726, 16'h7727 	:	val_out <= 16'h9ba9;
         16'h7728, 16'h7729, 16'h772a, 16'h772b, 16'h772c, 16'h772d, 16'h772e, 16'h772f 	:	val_out <= 16'h9b90;
         16'h7730, 16'h7731, 16'h7732, 16'h7733, 16'h7734, 16'h7735, 16'h7736, 16'h7737 	:	val_out <= 16'h9b78;
         16'h7738, 16'h7739, 16'h773a, 16'h773b, 16'h773c, 16'h773d, 16'h773e, 16'h773f 	:	val_out <= 16'h9b5f;
         16'h7740, 16'h7741, 16'h7742, 16'h7743, 16'h7744, 16'h7745, 16'h7746, 16'h7747 	:	val_out <= 16'h9b47;
         16'h7748, 16'h7749, 16'h774a, 16'h774b, 16'h774c, 16'h774d, 16'h774e, 16'h774f 	:	val_out <= 16'h9b2e;
         16'h7750, 16'h7751, 16'h7752, 16'h7753, 16'h7754, 16'h7755, 16'h7756, 16'h7757 	:	val_out <= 16'h9b16;
         16'h7758, 16'h7759, 16'h775a, 16'h775b, 16'h775c, 16'h775d, 16'h775e, 16'h775f 	:	val_out <= 16'h9afd;
         16'h7760, 16'h7761, 16'h7762, 16'h7763, 16'h7764, 16'h7765, 16'h7766, 16'h7767 	:	val_out <= 16'h9ae4;
         16'h7768, 16'h7769, 16'h776a, 16'h776b, 16'h776c, 16'h776d, 16'h776e, 16'h776f 	:	val_out <= 16'h9acc;
         16'h7770, 16'h7771, 16'h7772, 16'h7773, 16'h7774, 16'h7775, 16'h7776, 16'h7777 	:	val_out <= 16'h9ab3;
         16'h7778, 16'h7779, 16'h777a, 16'h777b, 16'h777c, 16'h777d, 16'h777e, 16'h777f 	:	val_out <= 16'h9a9b;
         16'h7780, 16'h7781, 16'h7782, 16'h7783, 16'h7784, 16'h7785, 16'h7786, 16'h7787 	:	val_out <= 16'h9a82;
         16'h7788, 16'h7789, 16'h778a, 16'h778b, 16'h778c, 16'h778d, 16'h778e, 16'h778f 	:	val_out <= 16'h9a6a;
         16'h7790, 16'h7791, 16'h7792, 16'h7793, 16'h7794, 16'h7795, 16'h7796, 16'h7797 	:	val_out <= 16'h9a51;
         16'h7798, 16'h7799, 16'h779a, 16'h779b, 16'h779c, 16'h779d, 16'h779e, 16'h779f 	:	val_out <= 16'h9a38;
         16'h77a0, 16'h77a1, 16'h77a2, 16'h77a3, 16'h77a4, 16'h77a5, 16'h77a6, 16'h77a7 	:	val_out <= 16'h9a20;
         16'h77a8, 16'h77a9, 16'h77aa, 16'h77ab, 16'h77ac, 16'h77ad, 16'h77ae, 16'h77af 	:	val_out <= 16'h9a07;
         16'h77b0, 16'h77b1, 16'h77b2, 16'h77b3, 16'h77b4, 16'h77b5, 16'h77b6, 16'h77b7 	:	val_out <= 16'h99ef;
         16'h77b8, 16'h77b9, 16'h77ba, 16'h77bb, 16'h77bc, 16'h77bd, 16'h77be, 16'h77bf 	:	val_out <= 16'h99d6;
         16'h77c0, 16'h77c1, 16'h77c2, 16'h77c3, 16'h77c4, 16'h77c5, 16'h77c6, 16'h77c7 	:	val_out <= 16'h99bd;
         16'h77c8, 16'h77c9, 16'h77ca, 16'h77cb, 16'h77cc, 16'h77cd, 16'h77ce, 16'h77cf 	:	val_out <= 16'h99a5;
         16'h77d0, 16'h77d1, 16'h77d2, 16'h77d3, 16'h77d4, 16'h77d5, 16'h77d6, 16'h77d7 	:	val_out <= 16'h998c;
         16'h77d8, 16'h77d9, 16'h77da, 16'h77db, 16'h77dc, 16'h77dd, 16'h77de, 16'h77df 	:	val_out <= 16'h9973;
         16'h77e0, 16'h77e1, 16'h77e2, 16'h77e3, 16'h77e4, 16'h77e5, 16'h77e6, 16'h77e7 	:	val_out <= 16'h995b;
         16'h77e8, 16'h77e9, 16'h77ea, 16'h77eb, 16'h77ec, 16'h77ed, 16'h77ee, 16'h77ef 	:	val_out <= 16'h9942;
         16'h77f0, 16'h77f1, 16'h77f2, 16'h77f3, 16'h77f4, 16'h77f5, 16'h77f6, 16'h77f7 	:	val_out <= 16'h992a;
         16'h77f8, 16'h77f9, 16'h77fa, 16'h77fb, 16'h77fc, 16'h77fd, 16'h77fe, 16'h77ff 	:	val_out <= 16'h9911;
         16'h7800, 16'h7801, 16'h7802, 16'h7803, 16'h7804, 16'h7805, 16'h7806, 16'h7807 	:	val_out <= 16'h98f8;
         16'h7808, 16'h7809, 16'h780a, 16'h780b, 16'h780c, 16'h780d, 16'h780e, 16'h780f 	:	val_out <= 16'h98e0;
         16'h7810, 16'h7811, 16'h7812, 16'h7813, 16'h7814, 16'h7815, 16'h7816, 16'h7817 	:	val_out <= 16'h98c7;
         16'h7818, 16'h7819, 16'h781a, 16'h781b, 16'h781c, 16'h781d, 16'h781e, 16'h781f 	:	val_out <= 16'h98ae;
         16'h7820, 16'h7821, 16'h7822, 16'h7823, 16'h7824, 16'h7825, 16'h7826, 16'h7827 	:	val_out <= 16'h9896;
         16'h7828, 16'h7829, 16'h782a, 16'h782b, 16'h782c, 16'h782d, 16'h782e, 16'h782f 	:	val_out <= 16'h987d;
         16'h7830, 16'h7831, 16'h7832, 16'h7833, 16'h7834, 16'h7835, 16'h7836, 16'h7837 	:	val_out <= 16'h9864;
         16'h7838, 16'h7839, 16'h783a, 16'h783b, 16'h783c, 16'h783d, 16'h783e, 16'h783f 	:	val_out <= 16'h984c;
         16'h7840, 16'h7841, 16'h7842, 16'h7843, 16'h7844, 16'h7845, 16'h7846, 16'h7847 	:	val_out <= 16'h9833;
         16'h7848, 16'h7849, 16'h784a, 16'h784b, 16'h784c, 16'h784d, 16'h784e, 16'h784f 	:	val_out <= 16'h981a;
         16'h7850, 16'h7851, 16'h7852, 16'h7853, 16'h7854, 16'h7855, 16'h7856, 16'h7857 	:	val_out <= 16'h9802;
         16'h7858, 16'h7859, 16'h785a, 16'h785b, 16'h785c, 16'h785d, 16'h785e, 16'h785f 	:	val_out <= 16'h97e9;
         16'h7860, 16'h7861, 16'h7862, 16'h7863, 16'h7864, 16'h7865, 16'h7866, 16'h7867 	:	val_out <= 16'h97d0;
         16'h7868, 16'h7869, 16'h786a, 16'h786b, 16'h786c, 16'h786d, 16'h786e, 16'h786f 	:	val_out <= 16'h97b7;
         16'h7870, 16'h7871, 16'h7872, 16'h7873, 16'h7874, 16'h7875, 16'h7876, 16'h7877 	:	val_out <= 16'h979f;
         16'h7878, 16'h7879, 16'h787a, 16'h787b, 16'h787c, 16'h787d, 16'h787e, 16'h787f 	:	val_out <= 16'h9786;
         16'h7880, 16'h7881, 16'h7882, 16'h7883, 16'h7884, 16'h7885, 16'h7886, 16'h7887 	:	val_out <= 16'h976d;
         16'h7888, 16'h7889, 16'h788a, 16'h788b, 16'h788c, 16'h788d, 16'h788e, 16'h788f 	:	val_out <= 16'h9755;
         16'h7890, 16'h7891, 16'h7892, 16'h7893, 16'h7894, 16'h7895, 16'h7896, 16'h7897 	:	val_out <= 16'h973c;
         16'h7898, 16'h7899, 16'h789a, 16'h789b, 16'h789c, 16'h789d, 16'h789e, 16'h789f 	:	val_out <= 16'h9723;
         16'h78a0, 16'h78a1, 16'h78a2, 16'h78a3, 16'h78a4, 16'h78a5, 16'h78a6, 16'h78a7 	:	val_out <= 16'h970a;
         16'h78a8, 16'h78a9, 16'h78aa, 16'h78ab, 16'h78ac, 16'h78ad, 16'h78ae, 16'h78af 	:	val_out <= 16'h96f2;
         16'h78b0, 16'h78b1, 16'h78b2, 16'h78b3, 16'h78b4, 16'h78b5, 16'h78b6, 16'h78b7 	:	val_out <= 16'h96d9;
         16'h78b8, 16'h78b9, 16'h78ba, 16'h78bb, 16'h78bc, 16'h78bd, 16'h78be, 16'h78bf 	:	val_out <= 16'h96c0;
         16'h78c0, 16'h78c1, 16'h78c2, 16'h78c3, 16'h78c4, 16'h78c5, 16'h78c6, 16'h78c7 	:	val_out <= 16'h96a8;
         16'h78c8, 16'h78c9, 16'h78ca, 16'h78cb, 16'h78cc, 16'h78cd, 16'h78ce, 16'h78cf 	:	val_out <= 16'h968f;
         16'h78d0, 16'h78d1, 16'h78d2, 16'h78d3, 16'h78d4, 16'h78d5, 16'h78d6, 16'h78d7 	:	val_out <= 16'h9676;
         16'h78d8, 16'h78d9, 16'h78da, 16'h78db, 16'h78dc, 16'h78dd, 16'h78de, 16'h78df 	:	val_out <= 16'h965d;
         16'h78e0, 16'h78e1, 16'h78e2, 16'h78e3, 16'h78e4, 16'h78e5, 16'h78e6, 16'h78e7 	:	val_out <= 16'h9645;
         16'h78e8, 16'h78e9, 16'h78ea, 16'h78eb, 16'h78ec, 16'h78ed, 16'h78ee, 16'h78ef 	:	val_out <= 16'h962c;
         16'h78f0, 16'h78f1, 16'h78f2, 16'h78f3, 16'h78f4, 16'h78f5, 16'h78f6, 16'h78f7 	:	val_out <= 16'h9613;
         16'h78f8, 16'h78f9, 16'h78fa, 16'h78fb, 16'h78fc, 16'h78fd, 16'h78fe, 16'h78ff 	:	val_out <= 16'h95fa;
         16'h7900, 16'h7901, 16'h7902, 16'h7903, 16'h7904, 16'h7905, 16'h7906, 16'h7907 	:	val_out <= 16'h95e2;
         16'h7908, 16'h7909, 16'h790a, 16'h790b, 16'h790c, 16'h790d, 16'h790e, 16'h790f 	:	val_out <= 16'h95c9;
         16'h7910, 16'h7911, 16'h7912, 16'h7913, 16'h7914, 16'h7915, 16'h7916, 16'h7917 	:	val_out <= 16'h95b0;
         16'h7918, 16'h7919, 16'h791a, 16'h791b, 16'h791c, 16'h791d, 16'h791e, 16'h791f 	:	val_out <= 16'h9597;
         16'h7920, 16'h7921, 16'h7922, 16'h7923, 16'h7924, 16'h7925, 16'h7926, 16'h7927 	:	val_out <= 16'h957f;
         16'h7928, 16'h7929, 16'h792a, 16'h792b, 16'h792c, 16'h792d, 16'h792e, 16'h792f 	:	val_out <= 16'h9566;
         16'h7930, 16'h7931, 16'h7932, 16'h7933, 16'h7934, 16'h7935, 16'h7936, 16'h7937 	:	val_out <= 16'h954d;
         16'h7938, 16'h7939, 16'h793a, 16'h793b, 16'h793c, 16'h793d, 16'h793e, 16'h793f 	:	val_out <= 16'h9534;
         16'h7940, 16'h7941, 16'h7942, 16'h7943, 16'h7944, 16'h7945, 16'h7946, 16'h7947 	:	val_out <= 16'h951b;
         16'h7948, 16'h7949, 16'h794a, 16'h794b, 16'h794c, 16'h794d, 16'h794e, 16'h794f 	:	val_out <= 16'h9503;
         16'h7950, 16'h7951, 16'h7952, 16'h7953, 16'h7954, 16'h7955, 16'h7956, 16'h7957 	:	val_out <= 16'h94ea;
         16'h7958, 16'h7959, 16'h795a, 16'h795b, 16'h795c, 16'h795d, 16'h795e, 16'h795f 	:	val_out <= 16'h94d1;
         16'h7960, 16'h7961, 16'h7962, 16'h7963, 16'h7964, 16'h7965, 16'h7966, 16'h7967 	:	val_out <= 16'h94b8;
         16'h7968, 16'h7969, 16'h796a, 16'h796b, 16'h796c, 16'h796d, 16'h796e, 16'h796f 	:	val_out <= 16'h949f;
         16'h7970, 16'h7971, 16'h7972, 16'h7973, 16'h7974, 16'h7975, 16'h7976, 16'h7977 	:	val_out <= 16'h9487;
         16'h7978, 16'h7979, 16'h797a, 16'h797b, 16'h797c, 16'h797d, 16'h797e, 16'h797f 	:	val_out <= 16'h946e;
         16'h7980, 16'h7981, 16'h7982, 16'h7983, 16'h7984, 16'h7985, 16'h7986, 16'h7987 	:	val_out <= 16'h9455;
         16'h7988, 16'h7989, 16'h798a, 16'h798b, 16'h798c, 16'h798d, 16'h798e, 16'h798f 	:	val_out <= 16'h943c;
         16'h7990, 16'h7991, 16'h7992, 16'h7993, 16'h7994, 16'h7995, 16'h7996, 16'h7997 	:	val_out <= 16'h9423;
         16'h7998, 16'h7999, 16'h799a, 16'h799b, 16'h799c, 16'h799d, 16'h799e, 16'h799f 	:	val_out <= 16'h940b;
         16'h79a0, 16'h79a1, 16'h79a2, 16'h79a3, 16'h79a4, 16'h79a5, 16'h79a6, 16'h79a7 	:	val_out <= 16'h93f2;
         16'h79a8, 16'h79a9, 16'h79aa, 16'h79ab, 16'h79ac, 16'h79ad, 16'h79ae, 16'h79af 	:	val_out <= 16'h93d9;
         16'h79b0, 16'h79b1, 16'h79b2, 16'h79b3, 16'h79b4, 16'h79b5, 16'h79b6, 16'h79b7 	:	val_out <= 16'h93c0;
         16'h79b8, 16'h79b9, 16'h79ba, 16'h79bb, 16'h79bc, 16'h79bd, 16'h79be, 16'h79bf 	:	val_out <= 16'h93a7;
         16'h79c0, 16'h79c1, 16'h79c2, 16'h79c3, 16'h79c4, 16'h79c5, 16'h79c6, 16'h79c7 	:	val_out <= 16'h938e;
         16'h79c8, 16'h79c9, 16'h79ca, 16'h79cb, 16'h79cc, 16'h79cd, 16'h79ce, 16'h79cf 	:	val_out <= 16'h9376;
         16'h79d0, 16'h79d1, 16'h79d2, 16'h79d3, 16'h79d4, 16'h79d5, 16'h79d6, 16'h79d7 	:	val_out <= 16'h935d;
         16'h79d8, 16'h79d9, 16'h79da, 16'h79db, 16'h79dc, 16'h79dd, 16'h79de, 16'h79df 	:	val_out <= 16'h9344;
         16'h79e0, 16'h79e1, 16'h79e2, 16'h79e3, 16'h79e4, 16'h79e5, 16'h79e6, 16'h79e7 	:	val_out <= 16'h932b;
         16'h79e8, 16'h79e9, 16'h79ea, 16'h79eb, 16'h79ec, 16'h79ed, 16'h79ee, 16'h79ef 	:	val_out <= 16'h9312;
         16'h79f0, 16'h79f1, 16'h79f2, 16'h79f3, 16'h79f4, 16'h79f5, 16'h79f6, 16'h79f7 	:	val_out <= 16'h92f9;
         16'h79f8, 16'h79f9, 16'h79fa, 16'h79fb, 16'h79fc, 16'h79fd, 16'h79fe, 16'h79ff 	:	val_out <= 16'h92e0;
         16'h7a00, 16'h7a01, 16'h7a02, 16'h7a03, 16'h7a04, 16'h7a05, 16'h7a06, 16'h7a07 	:	val_out <= 16'h92c8;
         16'h7a08, 16'h7a09, 16'h7a0a, 16'h7a0b, 16'h7a0c, 16'h7a0d, 16'h7a0e, 16'h7a0f 	:	val_out <= 16'h92af;
         16'h7a10, 16'h7a11, 16'h7a12, 16'h7a13, 16'h7a14, 16'h7a15, 16'h7a16, 16'h7a17 	:	val_out <= 16'h9296;
         16'h7a18, 16'h7a19, 16'h7a1a, 16'h7a1b, 16'h7a1c, 16'h7a1d, 16'h7a1e, 16'h7a1f 	:	val_out <= 16'h927d;
         16'h7a20, 16'h7a21, 16'h7a22, 16'h7a23, 16'h7a24, 16'h7a25, 16'h7a26, 16'h7a27 	:	val_out <= 16'h9264;
         16'h7a28, 16'h7a29, 16'h7a2a, 16'h7a2b, 16'h7a2c, 16'h7a2d, 16'h7a2e, 16'h7a2f 	:	val_out <= 16'h924b;
         16'h7a30, 16'h7a31, 16'h7a32, 16'h7a33, 16'h7a34, 16'h7a35, 16'h7a36, 16'h7a37 	:	val_out <= 16'h9232;
         16'h7a38, 16'h7a39, 16'h7a3a, 16'h7a3b, 16'h7a3c, 16'h7a3d, 16'h7a3e, 16'h7a3f 	:	val_out <= 16'h9219;
         16'h7a40, 16'h7a41, 16'h7a42, 16'h7a43, 16'h7a44, 16'h7a45, 16'h7a46, 16'h7a47 	:	val_out <= 16'h9201;
         16'h7a48, 16'h7a49, 16'h7a4a, 16'h7a4b, 16'h7a4c, 16'h7a4d, 16'h7a4e, 16'h7a4f 	:	val_out <= 16'h91e8;
         16'h7a50, 16'h7a51, 16'h7a52, 16'h7a53, 16'h7a54, 16'h7a55, 16'h7a56, 16'h7a57 	:	val_out <= 16'h91cf;
         16'h7a58, 16'h7a59, 16'h7a5a, 16'h7a5b, 16'h7a5c, 16'h7a5d, 16'h7a5e, 16'h7a5f 	:	val_out <= 16'h91b6;
         16'h7a60, 16'h7a61, 16'h7a62, 16'h7a63, 16'h7a64, 16'h7a65, 16'h7a66, 16'h7a67 	:	val_out <= 16'h919d;
         16'h7a68, 16'h7a69, 16'h7a6a, 16'h7a6b, 16'h7a6c, 16'h7a6d, 16'h7a6e, 16'h7a6f 	:	val_out <= 16'h9184;
         16'h7a70, 16'h7a71, 16'h7a72, 16'h7a73, 16'h7a74, 16'h7a75, 16'h7a76, 16'h7a77 	:	val_out <= 16'h916b;
         16'h7a78, 16'h7a79, 16'h7a7a, 16'h7a7b, 16'h7a7c, 16'h7a7d, 16'h7a7e, 16'h7a7f 	:	val_out <= 16'h9152;
         16'h7a80, 16'h7a81, 16'h7a82, 16'h7a83, 16'h7a84, 16'h7a85, 16'h7a86, 16'h7a87 	:	val_out <= 16'h9139;
         16'h7a88, 16'h7a89, 16'h7a8a, 16'h7a8b, 16'h7a8c, 16'h7a8d, 16'h7a8e, 16'h7a8f 	:	val_out <= 16'h9121;
         16'h7a90, 16'h7a91, 16'h7a92, 16'h7a93, 16'h7a94, 16'h7a95, 16'h7a96, 16'h7a97 	:	val_out <= 16'h9108;
         16'h7a98, 16'h7a99, 16'h7a9a, 16'h7a9b, 16'h7a9c, 16'h7a9d, 16'h7a9e, 16'h7a9f 	:	val_out <= 16'h90ef;
         16'h7aa0, 16'h7aa1, 16'h7aa2, 16'h7aa3, 16'h7aa4, 16'h7aa5, 16'h7aa6, 16'h7aa7 	:	val_out <= 16'h90d6;
         16'h7aa8, 16'h7aa9, 16'h7aaa, 16'h7aab, 16'h7aac, 16'h7aad, 16'h7aae, 16'h7aaf 	:	val_out <= 16'h90bd;
         16'h7ab0, 16'h7ab1, 16'h7ab2, 16'h7ab3, 16'h7ab4, 16'h7ab5, 16'h7ab6, 16'h7ab7 	:	val_out <= 16'h90a4;
         16'h7ab8, 16'h7ab9, 16'h7aba, 16'h7abb, 16'h7abc, 16'h7abd, 16'h7abe, 16'h7abf 	:	val_out <= 16'h908b;
         16'h7ac0, 16'h7ac1, 16'h7ac2, 16'h7ac3, 16'h7ac4, 16'h7ac5, 16'h7ac6, 16'h7ac7 	:	val_out <= 16'h9072;
         16'h7ac8, 16'h7ac9, 16'h7aca, 16'h7acb, 16'h7acc, 16'h7acd, 16'h7ace, 16'h7acf 	:	val_out <= 16'h9059;
         16'h7ad0, 16'h7ad1, 16'h7ad2, 16'h7ad3, 16'h7ad4, 16'h7ad5, 16'h7ad6, 16'h7ad7 	:	val_out <= 16'h9040;
         16'h7ad8, 16'h7ad9, 16'h7ada, 16'h7adb, 16'h7adc, 16'h7add, 16'h7ade, 16'h7adf 	:	val_out <= 16'h9027;
         16'h7ae0, 16'h7ae1, 16'h7ae2, 16'h7ae3, 16'h7ae4, 16'h7ae5, 16'h7ae6, 16'h7ae7 	:	val_out <= 16'h900e;
         16'h7ae8, 16'h7ae9, 16'h7aea, 16'h7aeb, 16'h7aec, 16'h7aed, 16'h7aee, 16'h7aef 	:	val_out <= 16'h8ff5;
         16'h7af0, 16'h7af1, 16'h7af2, 16'h7af3, 16'h7af4, 16'h7af5, 16'h7af6, 16'h7af7 	:	val_out <= 16'h8fdd;
         16'h7af8, 16'h7af9, 16'h7afa, 16'h7afb, 16'h7afc, 16'h7afd, 16'h7afe, 16'h7aff 	:	val_out <= 16'h8fc4;
         16'h7b00, 16'h7b01, 16'h7b02, 16'h7b03, 16'h7b04, 16'h7b05, 16'h7b06, 16'h7b07 	:	val_out <= 16'h8fab;
         16'h7b08, 16'h7b09, 16'h7b0a, 16'h7b0b, 16'h7b0c, 16'h7b0d, 16'h7b0e, 16'h7b0f 	:	val_out <= 16'h8f92;
         16'h7b10, 16'h7b11, 16'h7b12, 16'h7b13, 16'h7b14, 16'h7b15, 16'h7b16, 16'h7b17 	:	val_out <= 16'h8f79;
         16'h7b18, 16'h7b19, 16'h7b1a, 16'h7b1b, 16'h7b1c, 16'h7b1d, 16'h7b1e, 16'h7b1f 	:	val_out <= 16'h8f60;
         16'h7b20, 16'h7b21, 16'h7b22, 16'h7b23, 16'h7b24, 16'h7b25, 16'h7b26, 16'h7b27 	:	val_out <= 16'h8f47;
         16'h7b28, 16'h7b29, 16'h7b2a, 16'h7b2b, 16'h7b2c, 16'h7b2d, 16'h7b2e, 16'h7b2f 	:	val_out <= 16'h8f2e;
         16'h7b30, 16'h7b31, 16'h7b32, 16'h7b33, 16'h7b34, 16'h7b35, 16'h7b36, 16'h7b37 	:	val_out <= 16'h8f15;
         16'h7b38, 16'h7b39, 16'h7b3a, 16'h7b3b, 16'h7b3c, 16'h7b3d, 16'h7b3e, 16'h7b3f 	:	val_out <= 16'h8efc;
         16'h7b40, 16'h7b41, 16'h7b42, 16'h7b43, 16'h7b44, 16'h7b45, 16'h7b46, 16'h7b47 	:	val_out <= 16'h8ee3;
         16'h7b48, 16'h7b49, 16'h7b4a, 16'h7b4b, 16'h7b4c, 16'h7b4d, 16'h7b4e, 16'h7b4f 	:	val_out <= 16'h8eca;
         16'h7b50, 16'h7b51, 16'h7b52, 16'h7b53, 16'h7b54, 16'h7b55, 16'h7b56, 16'h7b57 	:	val_out <= 16'h8eb1;
         16'h7b58, 16'h7b59, 16'h7b5a, 16'h7b5b, 16'h7b5c, 16'h7b5d, 16'h7b5e, 16'h7b5f 	:	val_out <= 16'h8e98;
         16'h7b60, 16'h7b61, 16'h7b62, 16'h7b63, 16'h7b64, 16'h7b65, 16'h7b66, 16'h7b67 	:	val_out <= 16'h8e7f;
         16'h7b68, 16'h7b69, 16'h7b6a, 16'h7b6b, 16'h7b6c, 16'h7b6d, 16'h7b6e, 16'h7b6f 	:	val_out <= 16'h8e66;
         16'h7b70, 16'h7b71, 16'h7b72, 16'h7b73, 16'h7b74, 16'h7b75, 16'h7b76, 16'h7b77 	:	val_out <= 16'h8e4d;
         16'h7b78, 16'h7b79, 16'h7b7a, 16'h7b7b, 16'h7b7c, 16'h7b7d, 16'h7b7e, 16'h7b7f 	:	val_out <= 16'h8e34;
         16'h7b80, 16'h7b81, 16'h7b82, 16'h7b83, 16'h7b84, 16'h7b85, 16'h7b86, 16'h7b87 	:	val_out <= 16'h8e1b;
         16'h7b88, 16'h7b89, 16'h7b8a, 16'h7b8b, 16'h7b8c, 16'h7b8d, 16'h7b8e, 16'h7b8f 	:	val_out <= 16'h8e02;
         16'h7b90, 16'h7b91, 16'h7b92, 16'h7b93, 16'h7b94, 16'h7b95, 16'h7b96, 16'h7b97 	:	val_out <= 16'h8de9;
         16'h7b98, 16'h7b99, 16'h7b9a, 16'h7b9b, 16'h7b9c, 16'h7b9d, 16'h7b9e, 16'h7b9f 	:	val_out <= 16'h8dd0;
         16'h7ba0, 16'h7ba1, 16'h7ba2, 16'h7ba3, 16'h7ba4, 16'h7ba5, 16'h7ba6, 16'h7ba7 	:	val_out <= 16'h8db7;
         16'h7ba8, 16'h7ba9, 16'h7baa, 16'h7bab, 16'h7bac, 16'h7bad, 16'h7bae, 16'h7baf 	:	val_out <= 16'h8d9e;
         16'h7bb0, 16'h7bb1, 16'h7bb2, 16'h7bb3, 16'h7bb4, 16'h7bb5, 16'h7bb6, 16'h7bb7 	:	val_out <= 16'h8d85;
         16'h7bb8, 16'h7bb9, 16'h7bba, 16'h7bbb, 16'h7bbc, 16'h7bbd, 16'h7bbe, 16'h7bbf 	:	val_out <= 16'h8d6c;
         16'h7bc0, 16'h7bc1, 16'h7bc2, 16'h7bc3, 16'h7bc4, 16'h7bc5, 16'h7bc6, 16'h7bc7 	:	val_out <= 16'h8d53;
         16'h7bc8, 16'h7bc9, 16'h7bca, 16'h7bcb, 16'h7bcc, 16'h7bcd, 16'h7bce, 16'h7bcf 	:	val_out <= 16'h8d3a;
         16'h7bd0, 16'h7bd1, 16'h7bd2, 16'h7bd3, 16'h7bd4, 16'h7bd5, 16'h7bd6, 16'h7bd7 	:	val_out <= 16'h8d21;
         16'h7bd8, 16'h7bd9, 16'h7bda, 16'h7bdb, 16'h7bdc, 16'h7bdd, 16'h7bde, 16'h7bdf 	:	val_out <= 16'h8d08;
         16'h7be0, 16'h7be1, 16'h7be2, 16'h7be3, 16'h7be4, 16'h7be5, 16'h7be6, 16'h7be7 	:	val_out <= 16'h8cef;
         16'h7be8, 16'h7be9, 16'h7bea, 16'h7beb, 16'h7bec, 16'h7bed, 16'h7bee, 16'h7bef 	:	val_out <= 16'h8cd6;
         16'h7bf0, 16'h7bf1, 16'h7bf2, 16'h7bf3, 16'h7bf4, 16'h7bf5, 16'h7bf6, 16'h7bf7 	:	val_out <= 16'h8cbd;
         16'h7bf8, 16'h7bf9, 16'h7bfa, 16'h7bfb, 16'h7bfc, 16'h7bfd, 16'h7bfe, 16'h7bff 	:	val_out <= 16'h8ca4;
         16'h7c00, 16'h7c01, 16'h7c02, 16'h7c03, 16'h7c04, 16'h7c05, 16'h7c06, 16'h7c07 	:	val_out <= 16'h8c8b;
         16'h7c08, 16'h7c09, 16'h7c0a, 16'h7c0b, 16'h7c0c, 16'h7c0d, 16'h7c0e, 16'h7c0f 	:	val_out <= 16'h8c72;
         16'h7c10, 16'h7c11, 16'h7c12, 16'h7c13, 16'h7c14, 16'h7c15, 16'h7c16, 16'h7c17 	:	val_out <= 16'h8c59;
         16'h7c18, 16'h7c19, 16'h7c1a, 16'h7c1b, 16'h7c1c, 16'h7c1d, 16'h7c1e, 16'h7c1f 	:	val_out <= 16'h8c40;
         16'h7c20, 16'h7c21, 16'h7c22, 16'h7c23, 16'h7c24, 16'h7c25, 16'h7c26, 16'h7c27 	:	val_out <= 16'h8c27;
         16'h7c28, 16'h7c29, 16'h7c2a, 16'h7c2b, 16'h7c2c, 16'h7c2d, 16'h7c2e, 16'h7c2f 	:	val_out <= 16'h8c0e;
         16'h7c30, 16'h7c31, 16'h7c32, 16'h7c33, 16'h7c34, 16'h7c35, 16'h7c36, 16'h7c37 	:	val_out <= 16'h8bf5;
         16'h7c38, 16'h7c39, 16'h7c3a, 16'h7c3b, 16'h7c3c, 16'h7c3d, 16'h7c3e, 16'h7c3f 	:	val_out <= 16'h8bdc;
         16'h7c40, 16'h7c41, 16'h7c42, 16'h7c43, 16'h7c44, 16'h7c45, 16'h7c46, 16'h7c47 	:	val_out <= 16'h8bc3;
         16'h7c48, 16'h7c49, 16'h7c4a, 16'h7c4b, 16'h7c4c, 16'h7c4d, 16'h7c4e, 16'h7c4f 	:	val_out <= 16'h8baa;
         16'h7c50, 16'h7c51, 16'h7c52, 16'h7c53, 16'h7c54, 16'h7c55, 16'h7c56, 16'h7c57 	:	val_out <= 16'h8b91;
         16'h7c58, 16'h7c59, 16'h7c5a, 16'h7c5b, 16'h7c5c, 16'h7c5d, 16'h7c5e, 16'h7c5f 	:	val_out <= 16'h8b78;
         16'h7c60, 16'h7c61, 16'h7c62, 16'h7c63, 16'h7c64, 16'h7c65, 16'h7c66, 16'h7c67 	:	val_out <= 16'h8b5f;
         16'h7c68, 16'h7c69, 16'h7c6a, 16'h7c6b, 16'h7c6c, 16'h7c6d, 16'h7c6e, 16'h7c6f 	:	val_out <= 16'h8b46;
         16'h7c70, 16'h7c71, 16'h7c72, 16'h7c73, 16'h7c74, 16'h7c75, 16'h7c76, 16'h7c77 	:	val_out <= 16'h8b2d;
         16'h7c78, 16'h7c79, 16'h7c7a, 16'h7c7b, 16'h7c7c, 16'h7c7d, 16'h7c7e, 16'h7c7f 	:	val_out <= 16'h8b14;
         16'h7c80, 16'h7c81, 16'h7c82, 16'h7c83, 16'h7c84, 16'h7c85, 16'h7c86, 16'h7c87 	:	val_out <= 16'h8afb;
         16'h7c88, 16'h7c89, 16'h7c8a, 16'h7c8b, 16'h7c8c, 16'h7c8d, 16'h7c8e, 16'h7c8f 	:	val_out <= 16'h8ae2;
         16'h7c90, 16'h7c91, 16'h7c92, 16'h7c93, 16'h7c94, 16'h7c95, 16'h7c96, 16'h7c97 	:	val_out <= 16'h8ac9;
         16'h7c98, 16'h7c99, 16'h7c9a, 16'h7c9b, 16'h7c9c, 16'h7c9d, 16'h7c9e, 16'h7c9f 	:	val_out <= 16'h8ab0;
         16'h7ca0, 16'h7ca1, 16'h7ca2, 16'h7ca3, 16'h7ca4, 16'h7ca5, 16'h7ca6, 16'h7ca7 	:	val_out <= 16'h8a97;
         16'h7ca8, 16'h7ca9, 16'h7caa, 16'h7cab, 16'h7cac, 16'h7cad, 16'h7cae, 16'h7caf 	:	val_out <= 16'h8a7e;
         16'h7cb0, 16'h7cb1, 16'h7cb2, 16'h7cb3, 16'h7cb4, 16'h7cb5, 16'h7cb6, 16'h7cb7 	:	val_out <= 16'h8a65;
         16'h7cb8, 16'h7cb9, 16'h7cba, 16'h7cbb, 16'h7cbc, 16'h7cbd, 16'h7cbe, 16'h7cbf 	:	val_out <= 16'h8a4c;
         16'h7cc0, 16'h7cc1, 16'h7cc2, 16'h7cc3, 16'h7cc4, 16'h7cc5, 16'h7cc6, 16'h7cc7 	:	val_out <= 16'h8a33;
         16'h7cc8, 16'h7cc9, 16'h7cca, 16'h7ccb, 16'h7ccc, 16'h7ccd, 16'h7cce, 16'h7ccf 	:	val_out <= 16'h8a19;
         16'h7cd0, 16'h7cd1, 16'h7cd2, 16'h7cd3, 16'h7cd4, 16'h7cd5, 16'h7cd6, 16'h7cd7 	:	val_out <= 16'h8a00;
         16'h7cd8, 16'h7cd9, 16'h7cda, 16'h7cdb, 16'h7cdc, 16'h7cdd, 16'h7cde, 16'h7cdf 	:	val_out <= 16'h89e7;
         16'h7ce0, 16'h7ce1, 16'h7ce2, 16'h7ce3, 16'h7ce4, 16'h7ce5, 16'h7ce6, 16'h7ce7 	:	val_out <= 16'h89ce;
         16'h7ce8, 16'h7ce9, 16'h7cea, 16'h7ceb, 16'h7cec, 16'h7ced, 16'h7cee, 16'h7cef 	:	val_out <= 16'h89b5;
         16'h7cf0, 16'h7cf1, 16'h7cf2, 16'h7cf3, 16'h7cf4, 16'h7cf5, 16'h7cf6, 16'h7cf7 	:	val_out <= 16'h899c;
         16'h7cf8, 16'h7cf9, 16'h7cfa, 16'h7cfb, 16'h7cfc, 16'h7cfd, 16'h7cfe, 16'h7cff 	:	val_out <= 16'h8983;
         16'h7d00, 16'h7d01, 16'h7d02, 16'h7d03, 16'h7d04, 16'h7d05, 16'h7d06, 16'h7d07 	:	val_out <= 16'h896a;
         16'h7d08, 16'h7d09, 16'h7d0a, 16'h7d0b, 16'h7d0c, 16'h7d0d, 16'h7d0e, 16'h7d0f 	:	val_out <= 16'h8951;
         16'h7d10, 16'h7d11, 16'h7d12, 16'h7d13, 16'h7d14, 16'h7d15, 16'h7d16, 16'h7d17 	:	val_out <= 16'h8938;
         16'h7d18, 16'h7d19, 16'h7d1a, 16'h7d1b, 16'h7d1c, 16'h7d1d, 16'h7d1e, 16'h7d1f 	:	val_out <= 16'h891f;
         16'h7d20, 16'h7d21, 16'h7d22, 16'h7d23, 16'h7d24, 16'h7d25, 16'h7d26, 16'h7d27 	:	val_out <= 16'h8906;
         16'h7d28, 16'h7d29, 16'h7d2a, 16'h7d2b, 16'h7d2c, 16'h7d2d, 16'h7d2e, 16'h7d2f 	:	val_out <= 16'h88ed;
         16'h7d30, 16'h7d31, 16'h7d32, 16'h7d33, 16'h7d34, 16'h7d35, 16'h7d36, 16'h7d37 	:	val_out <= 16'h88d4;
         16'h7d38, 16'h7d39, 16'h7d3a, 16'h7d3b, 16'h7d3c, 16'h7d3d, 16'h7d3e, 16'h7d3f 	:	val_out <= 16'h88bb;
         16'h7d40, 16'h7d41, 16'h7d42, 16'h7d43, 16'h7d44, 16'h7d45, 16'h7d46, 16'h7d47 	:	val_out <= 16'h88a2;
         16'h7d48, 16'h7d49, 16'h7d4a, 16'h7d4b, 16'h7d4c, 16'h7d4d, 16'h7d4e, 16'h7d4f 	:	val_out <= 16'h8888;
         16'h7d50, 16'h7d51, 16'h7d52, 16'h7d53, 16'h7d54, 16'h7d55, 16'h7d56, 16'h7d57 	:	val_out <= 16'h886f;
         16'h7d58, 16'h7d59, 16'h7d5a, 16'h7d5b, 16'h7d5c, 16'h7d5d, 16'h7d5e, 16'h7d5f 	:	val_out <= 16'h8856;
         16'h7d60, 16'h7d61, 16'h7d62, 16'h7d63, 16'h7d64, 16'h7d65, 16'h7d66, 16'h7d67 	:	val_out <= 16'h883d;
         16'h7d68, 16'h7d69, 16'h7d6a, 16'h7d6b, 16'h7d6c, 16'h7d6d, 16'h7d6e, 16'h7d6f 	:	val_out <= 16'h8824;
         16'h7d70, 16'h7d71, 16'h7d72, 16'h7d73, 16'h7d74, 16'h7d75, 16'h7d76, 16'h7d77 	:	val_out <= 16'h880b;
         16'h7d78, 16'h7d79, 16'h7d7a, 16'h7d7b, 16'h7d7c, 16'h7d7d, 16'h7d7e, 16'h7d7f 	:	val_out <= 16'h87f2;
         16'h7d80, 16'h7d81, 16'h7d82, 16'h7d83, 16'h7d84, 16'h7d85, 16'h7d86, 16'h7d87 	:	val_out <= 16'h87d9;
         16'h7d88, 16'h7d89, 16'h7d8a, 16'h7d8b, 16'h7d8c, 16'h7d8d, 16'h7d8e, 16'h7d8f 	:	val_out <= 16'h87c0;
         16'h7d90, 16'h7d91, 16'h7d92, 16'h7d93, 16'h7d94, 16'h7d95, 16'h7d96, 16'h7d97 	:	val_out <= 16'h87a7;
         16'h7d98, 16'h7d99, 16'h7d9a, 16'h7d9b, 16'h7d9c, 16'h7d9d, 16'h7d9e, 16'h7d9f 	:	val_out <= 16'h878e;
         16'h7da0, 16'h7da1, 16'h7da2, 16'h7da3, 16'h7da4, 16'h7da5, 16'h7da6, 16'h7da7 	:	val_out <= 16'h8775;
         16'h7da8, 16'h7da9, 16'h7daa, 16'h7dab, 16'h7dac, 16'h7dad, 16'h7dae, 16'h7daf 	:	val_out <= 16'h875b;
         16'h7db0, 16'h7db1, 16'h7db2, 16'h7db3, 16'h7db4, 16'h7db5, 16'h7db6, 16'h7db7 	:	val_out <= 16'h8742;
         16'h7db8, 16'h7db9, 16'h7dba, 16'h7dbb, 16'h7dbc, 16'h7dbd, 16'h7dbe, 16'h7dbf 	:	val_out <= 16'h8729;
         16'h7dc0, 16'h7dc1, 16'h7dc2, 16'h7dc3, 16'h7dc4, 16'h7dc5, 16'h7dc6, 16'h7dc7 	:	val_out <= 16'h8710;
         16'h7dc8, 16'h7dc9, 16'h7dca, 16'h7dcb, 16'h7dcc, 16'h7dcd, 16'h7dce, 16'h7dcf 	:	val_out <= 16'h86f7;
         16'h7dd0, 16'h7dd1, 16'h7dd2, 16'h7dd3, 16'h7dd4, 16'h7dd5, 16'h7dd6, 16'h7dd7 	:	val_out <= 16'h86de;
         16'h7dd8, 16'h7dd9, 16'h7dda, 16'h7ddb, 16'h7ddc, 16'h7ddd, 16'h7dde, 16'h7ddf 	:	val_out <= 16'h86c5;
         16'h7de0, 16'h7de1, 16'h7de2, 16'h7de3, 16'h7de4, 16'h7de5, 16'h7de6, 16'h7de7 	:	val_out <= 16'h86ac;
         16'h7de8, 16'h7de9, 16'h7dea, 16'h7deb, 16'h7dec, 16'h7ded, 16'h7dee, 16'h7def 	:	val_out <= 16'h8693;
         16'h7df0, 16'h7df1, 16'h7df2, 16'h7df3, 16'h7df4, 16'h7df5, 16'h7df6, 16'h7df7 	:	val_out <= 16'h867a;
         16'h7df8, 16'h7df9, 16'h7dfa, 16'h7dfb, 16'h7dfc, 16'h7dfd, 16'h7dfe, 16'h7dff 	:	val_out <= 16'h8660;
         16'h7e00, 16'h7e01, 16'h7e02, 16'h7e03, 16'h7e04, 16'h7e05, 16'h7e06, 16'h7e07 	:	val_out <= 16'h8647;
         16'h7e08, 16'h7e09, 16'h7e0a, 16'h7e0b, 16'h7e0c, 16'h7e0d, 16'h7e0e, 16'h7e0f 	:	val_out <= 16'h862e;
         16'h7e10, 16'h7e11, 16'h7e12, 16'h7e13, 16'h7e14, 16'h7e15, 16'h7e16, 16'h7e17 	:	val_out <= 16'h8615;
         16'h7e18, 16'h7e19, 16'h7e1a, 16'h7e1b, 16'h7e1c, 16'h7e1d, 16'h7e1e, 16'h7e1f 	:	val_out <= 16'h85fc;
         16'h7e20, 16'h7e21, 16'h7e22, 16'h7e23, 16'h7e24, 16'h7e25, 16'h7e26, 16'h7e27 	:	val_out <= 16'h85e3;
         16'h7e28, 16'h7e29, 16'h7e2a, 16'h7e2b, 16'h7e2c, 16'h7e2d, 16'h7e2e, 16'h7e2f 	:	val_out <= 16'h85ca;
         16'h7e30, 16'h7e31, 16'h7e32, 16'h7e33, 16'h7e34, 16'h7e35, 16'h7e36, 16'h7e37 	:	val_out <= 16'h85b1;
         16'h7e38, 16'h7e39, 16'h7e3a, 16'h7e3b, 16'h7e3c, 16'h7e3d, 16'h7e3e, 16'h7e3f 	:	val_out <= 16'h8598;
         16'h7e40, 16'h7e41, 16'h7e42, 16'h7e43, 16'h7e44, 16'h7e45, 16'h7e46, 16'h7e47 	:	val_out <= 16'h857f;
         16'h7e48, 16'h7e49, 16'h7e4a, 16'h7e4b, 16'h7e4c, 16'h7e4d, 16'h7e4e, 16'h7e4f 	:	val_out <= 16'h8565;
         16'h7e50, 16'h7e51, 16'h7e52, 16'h7e53, 16'h7e54, 16'h7e55, 16'h7e56, 16'h7e57 	:	val_out <= 16'h854c;
         16'h7e58, 16'h7e59, 16'h7e5a, 16'h7e5b, 16'h7e5c, 16'h7e5d, 16'h7e5e, 16'h7e5f 	:	val_out <= 16'h8533;
         16'h7e60, 16'h7e61, 16'h7e62, 16'h7e63, 16'h7e64, 16'h7e65, 16'h7e66, 16'h7e67 	:	val_out <= 16'h851a;
         16'h7e68, 16'h7e69, 16'h7e6a, 16'h7e6b, 16'h7e6c, 16'h7e6d, 16'h7e6e, 16'h7e6f 	:	val_out <= 16'h8501;
         16'h7e70, 16'h7e71, 16'h7e72, 16'h7e73, 16'h7e74, 16'h7e75, 16'h7e76, 16'h7e77 	:	val_out <= 16'h84e8;
         16'h7e78, 16'h7e79, 16'h7e7a, 16'h7e7b, 16'h7e7c, 16'h7e7d, 16'h7e7e, 16'h7e7f 	:	val_out <= 16'h84cf;
         16'h7e80, 16'h7e81, 16'h7e82, 16'h7e83, 16'h7e84, 16'h7e85, 16'h7e86, 16'h7e87 	:	val_out <= 16'h84b6;
         16'h7e88, 16'h7e89, 16'h7e8a, 16'h7e8b, 16'h7e8c, 16'h7e8d, 16'h7e8e, 16'h7e8f 	:	val_out <= 16'h849c;
         16'h7e90, 16'h7e91, 16'h7e92, 16'h7e93, 16'h7e94, 16'h7e95, 16'h7e96, 16'h7e97 	:	val_out <= 16'h8483;
         16'h7e98, 16'h7e99, 16'h7e9a, 16'h7e9b, 16'h7e9c, 16'h7e9d, 16'h7e9e, 16'h7e9f 	:	val_out <= 16'h846a;
         16'h7ea0, 16'h7ea1, 16'h7ea2, 16'h7ea3, 16'h7ea4, 16'h7ea5, 16'h7ea6, 16'h7ea7 	:	val_out <= 16'h8451;
         16'h7ea8, 16'h7ea9, 16'h7eaa, 16'h7eab, 16'h7eac, 16'h7ead, 16'h7eae, 16'h7eaf 	:	val_out <= 16'h8438;
         16'h7eb0, 16'h7eb1, 16'h7eb2, 16'h7eb3, 16'h7eb4, 16'h7eb5, 16'h7eb6, 16'h7eb7 	:	val_out <= 16'h841f;
         16'h7eb8, 16'h7eb9, 16'h7eba, 16'h7ebb, 16'h7ebc, 16'h7ebd, 16'h7ebe, 16'h7ebf 	:	val_out <= 16'h8406;
         16'h7ec0, 16'h7ec1, 16'h7ec2, 16'h7ec3, 16'h7ec4, 16'h7ec5, 16'h7ec6, 16'h7ec7 	:	val_out <= 16'h83ed;
         16'h7ec8, 16'h7ec9, 16'h7eca, 16'h7ecb, 16'h7ecc, 16'h7ecd, 16'h7ece, 16'h7ecf 	:	val_out <= 16'h83d4;
         16'h7ed0, 16'h7ed1, 16'h7ed2, 16'h7ed3, 16'h7ed4, 16'h7ed5, 16'h7ed6, 16'h7ed7 	:	val_out <= 16'h83ba;
         16'h7ed8, 16'h7ed9, 16'h7eda, 16'h7edb, 16'h7edc, 16'h7edd, 16'h7ede, 16'h7edf 	:	val_out <= 16'h83a1;
         16'h7ee0, 16'h7ee1, 16'h7ee2, 16'h7ee3, 16'h7ee4, 16'h7ee5, 16'h7ee6, 16'h7ee7 	:	val_out <= 16'h8388;
         16'h7ee8, 16'h7ee9, 16'h7eea, 16'h7eeb, 16'h7eec, 16'h7eed, 16'h7eee, 16'h7eef 	:	val_out <= 16'h836f;
         16'h7ef0, 16'h7ef1, 16'h7ef2, 16'h7ef3, 16'h7ef4, 16'h7ef5, 16'h7ef6, 16'h7ef7 	:	val_out <= 16'h8356;
         16'h7ef8, 16'h7ef9, 16'h7efa, 16'h7efb, 16'h7efc, 16'h7efd, 16'h7efe, 16'h7eff 	:	val_out <= 16'h833d;
         16'h7f00, 16'h7f01, 16'h7f02, 16'h7f03, 16'h7f04, 16'h7f05, 16'h7f06, 16'h7f07 	:	val_out <= 16'h8324;
         16'h7f08, 16'h7f09, 16'h7f0a, 16'h7f0b, 16'h7f0c, 16'h7f0d, 16'h7f0e, 16'h7f0f 	:	val_out <= 16'h830b;
         16'h7f10, 16'h7f11, 16'h7f12, 16'h7f13, 16'h7f14, 16'h7f15, 16'h7f16, 16'h7f17 	:	val_out <= 16'h82f1;
         16'h7f18, 16'h7f19, 16'h7f1a, 16'h7f1b, 16'h7f1c, 16'h7f1d, 16'h7f1e, 16'h7f1f 	:	val_out <= 16'h82d8;
         16'h7f20, 16'h7f21, 16'h7f22, 16'h7f23, 16'h7f24, 16'h7f25, 16'h7f26, 16'h7f27 	:	val_out <= 16'h82bf;
         16'h7f28, 16'h7f29, 16'h7f2a, 16'h7f2b, 16'h7f2c, 16'h7f2d, 16'h7f2e, 16'h7f2f 	:	val_out <= 16'h82a6;
         16'h7f30, 16'h7f31, 16'h7f32, 16'h7f33, 16'h7f34, 16'h7f35, 16'h7f36, 16'h7f37 	:	val_out <= 16'h828d;
         16'h7f38, 16'h7f39, 16'h7f3a, 16'h7f3b, 16'h7f3c, 16'h7f3d, 16'h7f3e, 16'h7f3f 	:	val_out <= 16'h8274;
         16'h7f40, 16'h7f41, 16'h7f42, 16'h7f43, 16'h7f44, 16'h7f45, 16'h7f46, 16'h7f47 	:	val_out <= 16'h825b;
         16'h7f48, 16'h7f49, 16'h7f4a, 16'h7f4b, 16'h7f4c, 16'h7f4d, 16'h7f4e, 16'h7f4f 	:	val_out <= 16'h8242;
         16'h7f50, 16'h7f51, 16'h7f52, 16'h7f53, 16'h7f54, 16'h7f55, 16'h7f56, 16'h7f57 	:	val_out <= 16'h8228;
         16'h7f58, 16'h7f59, 16'h7f5a, 16'h7f5b, 16'h7f5c, 16'h7f5d, 16'h7f5e, 16'h7f5f 	:	val_out <= 16'h820f;
         16'h7f60, 16'h7f61, 16'h7f62, 16'h7f63, 16'h7f64, 16'h7f65, 16'h7f66, 16'h7f67 	:	val_out <= 16'h81f6;
         16'h7f68, 16'h7f69, 16'h7f6a, 16'h7f6b, 16'h7f6c, 16'h7f6d, 16'h7f6e, 16'h7f6f 	:	val_out <= 16'h81dd;
         16'h7f70, 16'h7f71, 16'h7f72, 16'h7f73, 16'h7f74, 16'h7f75, 16'h7f76, 16'h7f77 	:	val_out <= 16'h81c4;
         16'h7f78, 16'h7f79, 16'h7f7a, 16'h7f7b, 16'h7f7c, 16'h7f7d, 16'h7f7e, 16'h7f7f 	:	val_out <= 16'h81ab;
         16'h7f80, 16'h7f81, 16'h7f82, 16'h7f83, 16'h7f84, 16'h7f85, 16'h7f86, 16'h7f87 	:	val_out <= 16'h8192;
         16'h7f88, 16'h7f89, 16'h7f8a, 16'h7f8b, 16'h7f8c, 16'h7f8d, 16'h7f8e, 16'h7f8f 	:	val_out <= 16'h8178;
         16'h7f90, 16'h7f91, 16'h7f92, 16'h7f93, 16'h7f94, 16'h7f95, 16'h7f96, 16'h7f97 	:	val_out <= 16'h815f;
         16'h7f98, 16'h7f99, 16'h7f9a, 16'h7f9b, 16'h7f9c, 16'h7f9d, 16'h7f9e, 16'h7f9f 	:	val_out <= 16'h8146;
         16'h7fa0, 16'h7fa1, 16'h7fa2, 16'h7fa3, 16'h7fa4, 16'h7fa5, 16'h7fa6, 16'h7fa7 	:	val_out <= 16'h812d;
         16'h7fa8, 16'h7fa9, 16'h7faa, 16'h7fab, 16'h7fac, 16'h7fad, 16'h7fae, 16'h7faf 	:	val_out <= 16'h8114;
         16'h7fb0, 16'h7fb1, 16'h7fb2, 16'h7fb3, 16'h7fb4, 16'h7fb5, 16'h7fb6, 16'h7fb7 	:	val_out <= 16'h80fb;
         16'h7fb8, 16'h7fb9, 16'h7fba, 16'h7fbb, 16'h7fbc, 16'h7fbd, 16'h7fbe, 16'h7fbf 	:	val_out <= 16'h80e2;
         16'h7fc0, 16'h7fc1, 16'h7fc2, 16'h7fc3, 16'h7fc4, 16'h7fc5, 16'h7fc6, 16'h7fc7 	:	val_out <= 16'h80c9;
         16'h7fc8, 16'h7fc9, 16'h7fca, 16'h7fcb, 16'h7fcc, 16'h7fcd, 16'h7fce, 16'h7fcf 	:	val_out <= 16'h80af;
         16'h7fd0, 16'h7fd1, 16'h7fd2, 16'h7fd3, 16'h7fd4, 16'h7fd5, 16'h7fd6, 16'h7fd7 	:	val_out <= 16'h8096;
         16'h7fd8, 16'h7fd9, 16'h7fda, 16'h7fdb, 16'h7fdc, 16'h7fdd, 16'h7fde, 16'h7fdf 	:	val_out <= 16'h807d;
         16'h7fe0, 16'h7fe1, 16'h7fe2, 16'h7fe3, 16'h7fe4, 16'h7fe5, 16'h7fe6, 16'h7fe7 	:	val_out <= 16'h8064;
         16'h7fe8, 16'h7fe9, 16'h7fea, 16'h7feb, 16'h7fec, 16'h7fed, 16'h7fee, 16'h7fef 	:	val_out <= 16'h804b;
         16'h7ff0, 16'h7ff1, 16'h7ff2, 16'h7ff3, 16'h7ff4, 16'h7ff5, 16'h7ff6, 16'h7ff7 	:	val_out <= 16'h8032;
         16'h7ff8, 16'h7ff9, 16'h7ffa, 16'h7ffb, 16'h7ffc, 16'h7ffd, 16'h7ffe, 16'h7fff 	:	val_out <= 16'h8019;
         16'h8000, 16'h8001, 16'h8002, 16'h8003, 16'h8004, 16'h8005, 16'h8006, 16'h8007 	:	val_out <= 16'h8000;
         16'h8008, 16'h8009, 16'h800a, 16'h800b, 16'h800c, 16'h800d, 16'h800e, 16'h800f 	:	val_out <= 16'h7fe6;
         16'h8010, 16'h8011, 16'h8012, 16'h8013, 16'h8014, 16'h8015, 16'h8016, 16'h8017 	:	val_out <= 16'h7fcd;
         16'h8018, 16'h8019, 16'h801a, 16'h801b, 16'h801c, 16'h801d, 16'h801e, 16'h801f 	:	val_out <= 16'h7fb4;
         16'h8020, 16'h8021, 16'h8022, 16'h8023, 16'h8024, 16'h8025, 16'h8026, 16'h8027 	:	val_out <= 16'h7f9b;
         16'h8028, 16'h8029, 16'h802a, 16'h802b, 16'h802c, 16'h802d, 16'h802e, 16'h802f 	:	val_out <= 16'h7f82;
         16'h8030, 16'h8031, 16'h8032, 16'h8033, 16'h8034, 16'h8035, 16'h8036, 16'h8037 	:	val_out <= 16'h7f69;
         16'h8038, 16'h8039, 16'h803a, 16'h803b, 16'h803c, 16'h803d, 16'h803e, 16'h803f 	:	val_out <= 16'h7f50;
         16'h8040, 16'h8041, 16'h8042, 16'h8043, 16'h8044, 16'h8045, 16'h8046, 16'h8047 	:	val_out <= 16'h7f36;
         16'h8048, 16'h8049, 16'h804a, 16'h804b, 16'h804c, 16'h804d, 16'h804e, 16'h804f 	:	val_out <= 16'h7f1d;
         16'h8050, 16'h8051, 16'h8052, 16'h8053, 16'h8054, 16'h8055, 16'h8056, 16'h8057 	:	val_out <= 16'h7f04;
         16'h8058, 16'h8059, 16'h805a, 16'h805b, 16'h805c, 16'h805d, 16'h805e, 16'h805f 	:	val_out <= 16'h7eeb;
         16'h8060, 16'h8061, 16'h8062, 16'h8063, 16'h8064, 16'h8065, 16'h8066, 16'h8067 	:	val_out <= 16'h7ed2;
         16'h8068, 16'h8069, 16'h806a, 16'h806b, 16'h806c, 16'h806d, 16'h806e, 16'h806f 	:	val_out <= 16'h7eb9;
         16'h8070, 16'h8071, 16'h8072, 16'h8073, 16'h8074, 16'h8075, 16'h8076, 16'h8077 	:	val_out <= 16'h7ea0;
         16'h8078, 16'h8079, 16'h807a, 16'h807b, 16'h807c, 16'h807d, 16'h807e, 16'h807f 	:	val_out <= 16'h7e87;
         16'h8080, 16'h8081, 16'h8082, 16'h8083, 16'h8084, 16'h8085, 16'h8086, 16'h8087 	:	val_out <= 16'h7e6d;
         16'h8088, 16'h8089, 16'h808a, 16'h808b, 16'h808c, 16'h808d, 16'h808e, 16'h808f 	:	val_out <= 16'h7e54;
         16'h8090, 16'h8091, 16'h8092, 16'h8093, 16'h8094, 16'h8095, 16'h8096, 16'h8097 	:	val_out <= 16'h7e3b;
         16'h8098, 16'h8099, 16'h809a, 16'h809b, 16'h809c, 16'h809d, 16'h809e, 16'h809f 	:	val_out <= 16'h7e22;
         16'h80a0, 16'h80a1, 16'h80a2, 16'h80a3, 16'h80a4, 16'h80a5, 16'h80a6, 16'h80a7 	:	val_out <= 16'h7e09;
         16'h80a8, 16'h80a9, 16'h80aa, 16'h80ab, 16'h80ac, 16'h80ad, 16'h80ae, 16'h80af 	:	val_out <= 16'h7df0;
         16'h80b0, 16'h80b1, 16'h80b2, 16'h80b3, 16'h80b4, 16'h80b5, 16'h80b6, 16'h80b7 	:	val_out <= 16'h7dd7;
         16'h80b8, 16'h80b9, 16'h80ba, 16'h80bb, 16'h80bc, 16'h80bd, 16'h80be, 16'h80bf 	:	val_out <= 16'h7dbd;
         16'h80c0, 16'h80c1, 16'h80c2, 16'h80c3, 16'h80c4, 16'h80c5, 16'h80c6, 16'h80c7 	:	val_out <= 16'h7da4;
         16'h80c8, 16'h80c9, 16'h80ca, 16'h80cb, 16'h80cc, 16'h80cd, 16'h80ce, 16'h80cf 	:	val_out <= 16'h7d8b;
         16'h80d0, 16'h80d1, 16'h80d2, 16'h80d3, 16'h80d4, 16'h80d5, 16'h80d6, 16'h80d7 	:	val_out <= 16'h7d72;
         16'h80d8, 16'h80d9, 16'h80da, 16'h80db, 16'h80dc, 16'h80dd, 16'h80de, 16'h80df 	:	val_out <= 16'h7d59;
         16'h80e0, 16'h80e1, 16'h80e2, 16'h80e3, 16'h80e4, 16'h80e5, 16'h80e6, 16'h80e7 	:	val_out <= 16'h7d40;
         16'h80e8, 16'h80e9, 16'h80ea, 16'h80eb, 16'h80ec, 16'h80ed, 16'h80ee, 16'h80ef 	:	val_out <= 16'h7d27;
         16'h80f0, 16'h80f1, 16'h80f2, 16'h80f3, 16'h80f4, 16'h80f5, 16'h80f6, 16'h80f7 	:	val_out <= 16'h7d0e;
         16'h80f8, 16'h80f9, 16'h80fa, 16'h80fb, 16'h80fc, 16'h80fd, 16'h80fe, 16'h80ff 	:	val_out <= 16'h7cf4;
         16'h8100, 16'h8101, 16'h8102, 16'h8103, 16'h8104, 16'h8105, 16'h8106, 16'h8107 	:	val_out <= 16'h7cdb;
         16'h8108, 16'h8109, 16'h810a, 16'h810b, 16'h810c, 16'h810d, 16'h810e, 16'h810f 	:	val_out <= 16'h7cc2;
         16'h8110, 16'h8111, 16'h8112, 16'h8113, 16'h8114, 16'h8115, 16'h8116, 16'h8117 	:	val_out <= 16'h7ca9;
         16'h8118, 16'h8119, 16'h811a, 16'h811b, 16'h811c, 16'h811d, 16'h811e, 16'h811f 	:	val_out <= 16'h7c90;
         16'h8120, 16'h8121, 16'h8122, 16'h8123, 16'h8124, 16'h8125, 16'h8126, 16'h8127 	:	val_out <= 16'h7c77;
         16'h8128, 16'h8129, 16'h812a, 16'h812b, 16'h812c, 16'h812d, 16'h812e, 16'h812f 	:	val_out <= 16'h7c5e;
         16'h8130, 16'h8131, 16'h8132, 16'h8133, 16'h8134, 16'h8135, 16'h8136, 16'h8137 	:	val_out <= 16'h7c45;
         16'h8138, 16'h8139, 16'h813a, 16'h813b, 16'h813c, 16'h813d, 16'h813e, 16'h813f 	:	val_out <= 16'h7c2b;
         16'h8140, 16'h8141, 16'h8142, 16'h8143, 16'h8144, 16'h8145, 16'h8146, 16'h8147 	:	val_out <= 16'h7c12;
         16'h8148, 16'h8149, 16'h814a, 16'h814b, 16'h814c, 16'h814d, 16'h814e, 16'h814f 	:	val_out <= 16'h7bf9;
         16'h8150, 16'h8151, 16'h8152, 16'h8153, 16'h8154, 16'h8155, 16'h8156, 16'h8157 	:	val_out <= 16'h7be0;
         16'h8158, 16'h8159, 16'h815a, 16'h815b, 16'h815c, 16'h815d, 16'h815e, 16'h815f 	:	val_out <= 16'h7bc7;
         16'h8160, 16'h8161, 16'h8162, 16'h8163, 16'h8164, 16'h8165, 16'h8166, 16'h8167 	:	val_out <= 16'h7bae;
         16'h8168, 16'h8169, 16'h816a, 16'h816b, 16'h816c, 16'h816d, 16'h816e, 16'h816f 	:	val_out <= 16'h7b95;
         16'h8170, 16'h8171, 16'h8172, 16'h8173, 16'h8174, 16'h8175, 16'h8176, 16'h8177 	:	val_out <= 16'h7b7c;
         16'h8178, 16'h8179, 16'h817a, 16'h817b, 16'h817c, 16'h817d, 16'h817e, 16'h817f 	:	val_out <= 16'h7b63;
         16'h8180, 16'h8181, 16'h8182, 16'h8183, 16'h8184, 16'h8185, 16'h8186, 16'h8187 	:	val_out <= 16'h7b49;
         16'h8188, 16'h8189, 16'h818a, 16'h818b, 16'h818c, 16'h818d, 16'h818e, 16'h818f 	:	val_out <= 16'h7b30;
         16'h8190, 16'h8191, 16'h8192, 16'h8193, 16'h8194, 16'h8195, 16'h8196, 16'h8197 	:	val_out <= 16'h7b17;
         16'h8198, 16'h8199, 16'h819a, 16'h819b, 16'h819c, 16'h819d, 16'h819e, 16'h819f 	:	val_out <= 16'h7afe;
         16'h81a0, 16'h81a1, 16'h81a2, 16'h81a3, 16'h81a4, 16'h81a5, 16'h81a6, 16'h81a7 	:	val_out <= 16'h7ae5;
         16'h81a8, 16'h81a9, 16'h81aa, 16'h81ab, 16'h81ac, 16'h81ad, 16'h81ae, 16'h81af 	:	val_out <= 16'h7acc;
         16'h81b0, 16'h81b1, 16'h81b2, 16'h81b3, 16'h81b4, 16'h81b5, 16'h81b6, 16'h81b7 	:	val_out <= 16'h7ab3;
         16'h81b8, 16'h81b9, 16'h81ba, 16'h81bb, 16'h81bc, 16'h81bd, 16'h81be, 16'h81bf 	:	val_out <= 16'h7a9a;
         16'h81c0, 16'h81c1, 16'h81c2, 16'h81c3, 16'h81c4, 16'h81c5, 16'h81c6, 16'h81c7 	:	val_out <= 16'h7a80;
         16'h81c8, 16'h81c9, 16'h81ca, 16'h81cb, 16'h81cc, 16'h81cd, 16'h81ce, 16'h81cf 	:	val_out <= 16'h7a67;
         16'h81d0, 16'h81d1, 16'h81d2, 16'h81d3, 16'h81d4, 16'h81d5, 16'h81d6, 16'h81d7 	:	val_out <= 16'h7a4e;
         16'h81d8, 16'h81d9, 16'h81da, 16'h81db, 16'h81dc, 16'h81dd, 16'h81de, 16'h81df 	:	val_out <= 16'h7a35;
         16'h81e0, 16'h81e1, 16'h81e2, 16'h81e3, 16'h81e4, 16'h81e5, 16'h81e6, 16'h81e7 	:	val_out <= 16'h7a1c;
         16'h81e8, 16'h81e9, 16'h81ea, 16'h81eb, 16'h81ec, 16'h81ed, 16'h81ee, 16'h81ef 	:	val_out <= 16'h7a03;
         16'h81f0, 16'h81f1, 16'h81f2, 16'h81f3, 16'h81f4, 16'h81f5, 16'h81f6, 16'h81f7 	:	val_out <= 16'h79ea;
         16'h81f8, 16'h81f9, 16'h81fa, 16'h81fb, 16'h81fc, 16'h81fd, 16'h81fe, 16'h81ff 	:	val_out <= 16'h79d1;
         16'h8200, 16'h8201, 16'h8202, 16'h8203, 16'h8204, 16'h8205, 16'h8206, 16'h8207 	:	val_out <= 16'h79b8;
         16'h8208, 16'h8209, 16'h820a, 16'h820b, 16'h820c, 16'h820d, 16'h820e, 16'h820f 	:	val_out <= 16'h799f;
         16'h8210, 16'h8211, 16'h8212, 16'h8213, 16'h8214, 16'h8215, 16'h8216, 16'h8217 	:	val_out <= 16'h7985;
         16'h8218, 16'h8219, 16'h821a, 16'h821b, 16'h821c, 16'h821d, 16'h821e, 16'h821f 	:	val_out <= 16'h796c;
         16'h8220, 16'h8221, 16'h8222, 16'h8223, 16'h8224, 16'h8225, 16'h8226, 16'h8227 	:	val_out <= 16'h7953;
         16'h8228, 16'h8229, 16'h822a, 16'h822b, 16'h822c, 16'h822d, 16'h822e, 16'h822f 	:	val_out <= 16'h793a;
         16'h8230, 16'h8231, 16'h8232, 16'h8233, 16'h8234, 16'h8235, 16'h8236, 16'h8237 	:	val_out <= 16'h7921;
         16'h8238, 16'h8239, 16'h823a, 16'h823b, 16'h823c, 16'h823d, 16'h823e, 16'h823f 	:	val_out <= 16'h7908;
         16'h8240, 16'h8241, 16'h8242, 16'h8243, 16'h8244, 16'h8245, 16'h8246, 16'h8247 	:	val_out <= 16'h78ef;
         16'h8248, 16'h8249, 16'h824a, 16'h824b, 16'h824c, 16'h824d, 16'h824e, 16'h824f 	:	val_out <= 16'h78d6;
         16'h8250, 16'h8251, 16'h8252, 16'h8253, 16'h8254, 16'h8255, 16'h8256, 16'h8257 	:	val_out <= 16'h78bd;
         16'h8258, 16'h8259, 16'h825a, 16'h825b, 16'h825c, 16'h825d, 16'h825e, 16'h825f 	:	val_out <= 16'h78a4;
         16'h8260, 16'h8261, 16'h8262, 16'h8263, 16'h8264, 16'h8265, 16'h8266, 16'h8267 	:	val_out <= 16'h788a;
         16'h8268, 16'h8269, 16'h826a, 16'h826b, 16'h826c, 16'h826d, 16'h826e, 16'h826f 	:	val_out <= 16'h7871;
         16'h8270, 16'h8271, 16'h8272, 16'h8273, 16'h8274, 16'h8275, 16'h8276, 16'h8277 	:	val_out <= 16'h7858;
         16'h8278, 16'h8279, 16'h827a, 16'h827b, 16'h827c, 16'h827d, 16'h827e, 16'h827f 	:	val_out <= 16'h783f;
         16'h8280, 16'h8281, 16'h8282, 16'h8283, 16'h8284, 16'h8285, 16'h8286, 16'h8287 	:	val_out <= 16'h7826;
         16'h8288, 16'h8289, 16'h828a, 16'h828b, 16'h828c, 16'h828d, 16'h828e, 16'h828f 	:	val_out <= 16'h780d;
         16'h8290, 16'h8291, 16'h8292, 16'h8293, 16'h8294, 16'h8295, 16'h8296, 16'h8297 	:	val_out <= 16'h77f4;
         16'h8298, 16'h8299, 16'h829a, 16'h829b, 16'h829c, 16'h829d, 16'h829e, 16'h829f 	:	val_out <= 16'h77db;
         16'h82a0, 16'h82a1, 16'h82a2, 16'h82a3, 16'h82a4, 16'h82a5, 16'h82a6, 16'h82a7 	:	val_out <= 16'h77c2;
         16'h82a8, 16'h82a9, 16'h82aa, 16'h82ab, 16'h82ac, 16'h82ad, 16'h82ae, 16'h82af 	:	val_out <= 16'h77a9;
         16'h82b0, 16'h82b1, 16'h82b2, 16'h82b3, 16'h82b4, 16'h82b5, 16'h82b6, 16'h82b7 	:	val_out <= 16'h7790;
         16'h82b8, 16'h82b9, 16'h82ba, 16'h82bb, 16'h82bc, 16'h82bd, 16'h82be, 16'h82bf 	:	val_out <= 16'h7777;
         16'h82c0, 16'h82c1, 16'h82c2, 16'h82c3, 16'h82c4, 16'h82c5, 16'h82c6, 16'h82c7 	:	val_out <= 16'h775d;
         16'h82c8, 16'h82c9, 16'h82ca, 16'h82cb, 16'h82cc, 16'h82cd, 16'h82ce, 16'h82cf 	:	val_out <= 16'h7744;
         16'h82d0, 16'h82d1, 16'h82d2, 16'h82d3, 16'h82d4, 16'h82d5, 16'h82d6, 16'h82d7 	:	val_out <= 16'h772b;
         16'h82d8, 16'h82d9, 16'h82da, 16'h82db, 16'h82dc, 16'h82dd, 16'h82de, 16'h82df 	:	val_out <= 16'h7712;
         16'h82e0, 16'h82e1, 16'h82e2, 16'h82e3, 16'h82e4, 16'h82e5, 16'h82e6, 16'h82e7 	:	val_out <= 16'h76f9;
         16'h82e8, 16'h82e9, 16'h82ea, 16'h82eb, 16'h82ec, 16'h82ed, 16'h82ee, 16'h82ef 	:	val_out <= 16'h76e0;
         16'h82f0, 16'h82f1, 16'h82f2, 16'h82f3, 16'h82f4, 16'h82f5, 16'h82f6, 16'h82f7 	:	val_out <= 16'h76c7;
         16'h82f8, 16'h82f9, 16'h82fa, 16'h82fb, 16'h82fc, 16'h82fd, 16'h82fe, 16'h82ff 	:	val_out <= 16'h76ae;
         16'h8300, 16'h8301, 16'h8302, 16'h8303, 16'h8304, 16'h8305, 16'h8306, 16'h8307 	:	val_out <= 16'h7695;
         16'h8308, 16'h8309, 16'h830a, 16'h830b, 16'h830c, 16'h830d, 16'h830e, 16'h830f 	:	val_out <= 16'h767c;
         16'h8310, 16'h8311, 16'h8312, 16'h8313, 16'h8314, 16'h8315, 16'h8316, 16'h8317 	:	val_out <= 16'h7663;
         16'h8318, 16'h8319, 16'h831a, 16'h831b, 16'h831c, 16'h831d, 16'h831e, 16'h831f 	:	val_out <= 16'h764a;
         16'h8320, 16'h8321, 16'h8322, 16'h8323, 16'h8324, 16'h8325, 16'h8326, 16'h8327 	:	val_out <= 16'h7631;
         16'h8328, 16'h8329, 16'h832a, 16'h832b, 16'h832c, 16'h832d, 16'h832e, 16'h832f 	:	val_out <= 16'h7618;
         16'h8330, 16'h8331, 16'h8332, 16'h8333, 16'h8334, 16'h8335, 16'h8336, 16'h8337 	:	val_out <= 16'h75ff;
         16'h8338, 16'h8339, 16'h833a, 16'h833b, 16'h833c, 16'h833d, 16'h833e, 16'h833f 	:	val_out <= 16'h75e6;
         16'h8340, 16'h8341, 16'h8342, 16'h8343, 16'h8344, 16'h8345, 16'h8346, 16'h8347 	:	val_out <= 16'h75cc;
         16'h8348, 16'h8349, 16'h834a, 16'h834b, 16'h834c, 16'h834d, 16'h834e, 16'h834f 	:	val_out <= 16'h75b3;
         16'h8350, 16'h8351, 16'h8352, 16'h8353, 16'h8354, 16'h8355, 16'h8356, 16'h8357 	:	val_out <= 16'h759a;
         16'h8358, 16'h8359, 16'h835a, 16'h835b, 16'h835c, 16'h835d, 16'h835e, 16'h835f 	:	val_out <= 16'h7581;
         16'h8360, 16'h8361, 16'h8362, 16'h8363, 16'h8364, 16'h8365, 16'h8366, 16'h8367 	:	val_out <= 16'h7568;
         16'h8368, 16'h8369, 16'h836a, 16'h836b, 16'h836c, 16'h836d, 16'h836e, 16'h836f 	:	val_out <= 16'h754f;
         16'h8370, 16'h8371, 16'h8372, 16'h8373, 16'h8374, 16'h8375, 16'h8376, 16'h8377 	:	val_out <= 16'h7536;
         16'h8378, 16'h8379, 16'h837a, 16'h837b, 16'h837c, 16'h837d, 16'h837e, 16'h837f 	:	val_out <= 16'h751d;
         16'h8380, 16'h8381, 16'h8382, 16'h8383, 16'h8384, 16'h8385, 16'h8386, 16'h8387 	:	val_out <= 16'h7504;
         16'h8388, 16'h8389, 16'h838a, 16'h838b, 16'h838c, 16'h838d, 16'h838e, 16'h838f 	:	val_out <= 16'h74eb;
         16'h8390, 16'h8391, 16'h8392, 16'h8393, 16'h8394, 16'h8395, 16'h8396, 16'h8397 	:	val_out <= 16'h74d2;
         16'h8398, 16'h8399, 16'h839a, 16'h839b, 16'h839c, 16'h839d, 16'h839e, 16'h839f 	:	val_out <= 16'h74b9;
         16'h83a0, 16'h83a1, 16'h83a2, 16'h83a3, 16'h83a4, 16'h83a5, 16'h83a6, 16'h83a7 	:	val_out <= 16'h74a0;
         16'h83a8, 16'h83a9, 16'h83aa, 16'h83ab, 16'h83ac, 16'h83ad, 16'h83ae, 16'h83af 	:	val_out <= 16'h7487;
         16'h83b0, 16'h83b1, 16'h83b2, 16'h83b3, 16'h83b4, 16'h83b5, 16'h83b6, 16'h83b7 	:	val_out <= 16'h746e;
         16'h83b8, 16'h83b9, 16'h83ba, 16'h83bb, 16'h83bc, 16'h83bd, 16'h83be, 16'h83bf 	:	val_out <= 16'h7455;
         16'h83c0, 16'h83c1, 16'h83c2, 16'h83c3, 16'h83c4, 16'h83c5, 16'h83c6, 16'h83c7 	:	val_out <= 16'h743c;
         16'h83c8, 16'h83c9, 16'h83ca, 16'h83cb, 16'h83cc, 16'h83cd, 16'h83ce, 16'h83cf 	:	val_out <= 16'h7423;
         16'h83d0, 16'h83d1, 16'h83d2, 16'h83d3, 16'h83d4, 16'h83d5, 16'h83d6, 16'h83d7 	:	val_out <= 16'h740a;
         16'h83d8, 16'h83d9, 16'h83da, 16'h83db, 16'h83dc, 16'h83dd, 16'h83de, 16'h83df 	:	val_out <= 16'h73f1;
         16'h83e0, 16'h83e1, 16'h83e2, 16'h83e3, 16'h83e4, 16'h83e5, 16'h83e6, 16'h83e7 	:	val_out <= 16'h73d8;
         16'h83e8, 16'h83e9, 16'h83ea, 16'h83eb, 16'h83ec, 16'h83ed, 16'h83ee, 16'h83ef 	:	val_out <= 16'h73bf;
         16'h83f0, 16'h83f1, 16'h83f2, 16'h83f3, 16'h83f4, 16'h83f5, 16'h83f6, 16'h83f7 	:	val_out <= 16'h73a6;
         16'h83f8, 16'h83f9, 16'h83fa, 16'h83fb, 16'h83fc, 16'h83fd, 16'h83fe, 16'h83ff 	:	val_out <= 16'h738d;
         16'h8400, 16'h8401, 16'h8402, 16'h8403, 16'h8404, 16'h8405, 16'h8406, 16'h8407 	:	val_out <= 16'h7374;
         16'h8408, 16'h8409, 16'h840a, 16'h840b, 16'h840c, 16'h840d, 16'h840e, 16'h840f 	:	val_out <= 16'h735b;
         16'h8410, 16'h8411, 16'h8412, 16'h8413, 16'h8414, 16'h8415, 16'h8416, 16'h8417 	:	val_out <= 16'h7342;
         16'h8418, 16'h8419, 16'h841a, 16'h841b, 16'h841c, 16'h841d, 16'h841e, 16'h841f 	:	val_out <= 16'h7329;
         16'h8420, 16'h8421, 16'h8422, 16'h8423, 16'h8424, 16'h8425, 16'h8426, 16'h8427 	:	val_out <= 16'h7310;
         16'h8428, 16'h8429, 16'h842a, 16'h842b, 16'h842c, 16'h842d, 16'h842e, 16'h842f 	:	val_out <= 16'h72f7;
         16'h8430, 16'h8431, 16'h8432, 16'h8433, 16'h8434, 16'h8435, 16'h8436, 16'h8437 	:	val_out <= 16'h72de;
         16'h8438, 16'h8439, 16'h843a, 16'h843b, 16'h843c, 16'h843d, 16'h843e, 16'h843f 	:	val_out <= 16'h72c5;
         16'h8440, 16'h8441, 16'h8442, 16'h8443, 16'h8444, 16'h8445, 16'h8446, 16'h8447 	:	val_out <= 16'h72ac;
         16'h8448, 16'h8449, 16'h844a, 16'h844b, 16'h844c, 16'h844d, 16'h844e, 16'h844f 	:	val_out <= 16'h7293;
         16'h8450, 16'h8451, 16'h8452, 16'h8453, 16'h8454, 16'h8455, 16'h8456, 16'h8457 	:	val_out <= 16'h727a;
         16'h8458, 16'h8459, 16'h845a, 16'h845b, 16'h845c, 16'h845d, 16'h845e, 16'h845f 	:	val_out <= 16'h7261;
         16'h8460, 16'h8461, 16'h8462, 16'h8463, 16'h8464, 16'h8465, 16'h8466, 16'h8467 	:	val_out <= 16'h7248;
         16'h8468, 16'h8469, 16'h846a, 16'h846b, 16'h846c, 16'h846d, 16'h846e, 16'h846f 	:	val_out <= 16'h722f;
         16'h8470, 16'h8471, 16'h8472, 16'h8473, 16'h8474, 16'h8475, 16'h8476, 16'h8477 	:	val_out <= 16'h7216;
         16'h8478, 16'h8479, 16'h847a, 16'h847b, 16'h847c, 16'h847d, 16'h847e, 16'h847f 	:	val_out <= 16'h71fd;
         16'h8480, 16'h8481, 16'h8482, 16'h8483, 16'h8484, 16'h8485, 16'h8486, 16'h8487 	:	val_out <= 16'h71e4;
         16'h8488, 16'h8489, 16'h848a, 16'h848b, 16'h848c, 16'h848d, 16'h848e, 16'h848f 	:	val_out <= 16'h71cb;
         16'h8490, 16'h8491, 16'h8492, 16'h8493, 16'h8494, 16'h8495, 16'h8496, 16'h8497 	:	val_out <= 16'h71b2;
         16'h8498, 16'h8499, 16'h849a, 16'h849b, 16'h849c, 16'h849d, 16'h849e, 16'h849f 	:	val_out <= 16'h7199;
         16'h84a0, 16'h84a1, 16'h84a2, 16'h84a3, 16'h84a4, 16'h84a5, 16'h84a6, 16'h84a7 	:	val_out <= 16'h7180;
         16'h84a8, 16'h84a9, 16'h84aa, 16'h84ab, 16'h84ac, 16'h84ad, 16'h84ae, 16'h84af 	:	val_out <= 16'h7167;
         16'h84b0, 16'h84b1, 16'h84b2, 16'h84b3, 16'h84b4, 16'h84b5, 16'h84b6, 16'h84b7 	:	val_out <= 16'h714e;
         16'h84b8, 16'h84b9, 16'h84ba, 16'h84bb, 16'h84bc, 16'h84bd, 16'h84be, 16'h84bf 	:	val_out <= 16'h7135;
         16'h84c0, 16'h84c1, 16'h84c2, 16'h84c3, 16'h84c4, 16'h84c5, 16'h84c6, 16'h84c7 	:	val_out <= 16'h711c;
         16'h84c8, 16'h84c9, 16'h84ca, 16'h84cb, 16'h84cc, 16'h84cd, 16'h84ce, 16'h84cf 	:	val_out <= 16'h7103;
         16'h84d0, 16'h84d1, 16'h84d2, 16'h84d3, 16'h84d4, 16'h84d5, 16'h84d6, 16'h84d7 	:	val_out <= 16'h70ea;
         16'h84d8, 16'h84d9, 16'h84da, 16'h84db, 16'h84dc, 16'h84dd, 16'h84de, 16'h84df 	:	val_out <= 16'h70d1;
         16'h84e0, 16'h84e1, 16'h84e2, 16'h84e3, 16'h84e4, 16'h84e5, 16'h84e6, 16'h84e7 	:	val_out <= 16'h70b8;
         16'h84e8, 16'h84e9, 16'h84ea, 16'h84eb, 16'h84ec, 16'h84ed, 16'h84ee, 16'h84ef 	:	val_out <= 16'h709f;
         16'h84f0, 16'h84f1, 16'h84f2, 16'h84f3, 16'h84f4, 16'h84f5, 16'h84f6, 16'h84f7 	:	val_out <= 16'h7086;
         16'h84f8, 16'h84f9, 16'h84fa, 16'h84fb, 16'h84fc, 16'h84fd, 16'h84fe, 16'h84ff 	:	val_out <= 16'h706d;
         16'h8500, 16'h8501, 16'h8502, 16'h8503, 16'h8504, 16'h8505, 16'h8506, 16'h8507 	:	val_out <= 16'h7054;
         16'h8508, 16'h8509, 16'h850a, 16'h850b, 16'h850c, 16'h850d, 16'h850e, 16'h850f 	:	val_out <= 16'h703b;
         16'h8510, 16'h8511, 16'h8512, 16'h8513, 16'h8514, 16'h8515, 16'h8516, 16'h8517 	:	val_out <= 16'h7022;
         16'h8518, 16'h8519, 16'h851a, 16'h851b, 16'h851c, 16'h851d, 16'h851e, 16'h851f 	:	val_out <= 16'h700a;
         16'h8520, 16'h8521, 16'h8522, 16'h8523, 16'h8524, 16'h8525, 16'h8526, 16'h8527 	:	val_out <= 16'h6ff1;
         16'h8528, 16'h8529, 16'h852a, 16'h852b, 16'h852c, 16'h852d, 16'h852e, 16'h852f 	:	val_out <= 16'h6fd8;
         16'h8530, 16'h8531, 16'h8532, 16'h8533, 16'h8534, 16'h8535, 16'h8536, 16'h8537 	:	val_out <= 16'h6fbf;
         16'h8538, 16'h8539, 16'h853a, 16'h853b, 16'h853c, 16'h853d, 16'h853e, 16'h853f 	:	val_out <= 16'h6fa6;
         16'h8540, 16'h8541, 16'h8542, 16'h8543, 16'h8544, 16'h8545, 16'h8546, 16'h8547 	:	val_out <= 16'h6f8d;
         16'h8548, 16'h8549, 16'h854a, 16'h854b, 16'h854c, 16'h854d, 16'h854e, 16'h854f 	:	val_out <= 16'h6f74;
         16'h8550, 16'h8551, 16'h8552, 16'h8553, 16'h8554, 16'h8555, 16'h8556, 16'h8557 	:	val_out <= 16'h6f5b;
         16'h8558, 16'h8559, 16'h855a, 16'h855b, 16'h855c, 16'h855d, 16'h855e, 16'h855f 	:	val_out <= 16'h6f42;
         16'h8560, 16'h8561, 16'h8562, 16'h8563, 16'h8564, 16'h8565, 16'h8566, 16'h8567 	:	val_out <= 16'h6f29;
         16'h8568, 16'h8569, 16'h856a, 16'h856b, 16'h856c, 16'h856d, 16'h856e, 16'h856f 	:	val_out <= 16'h6f10;
         16'h8570, 16'h8571, 16'h8572, 16'h8573, 16'h8574, 16'h8575, 16'h8576, 16'h8577 	:	val_out <= 16'h6ef7;
         16'h8578, 16'h8579, 16'h857a, 16'h857b, 16'h857c, 16'h857d, 16'h857e, 16'h857f 	:	val_out <= 16'h6ede;
         16'h8580, 16'h8581, 16'h8582, 16'h8583, 16'h8584, 16'h8585, 16'h8586, 16'h8587 	:	val_out <= 16'h6ec6;
         16'h8588, 16'h8589, 16'h858a, 16'h858b, 16'h858c, 16'h858d, 16'h858e, 16'h858f 	:	val_out <= 16'h6ead;
         16'h8590, 16'h8591, 16'h8592, 16'h8593, 16'h8594, 16'h8595, 16'h8596, 16'h8597 	:	val_out <= 16'h6e94;
         16'h8598, 16'h8599, 16'h859a, 16'h859b, 16'h859c, 16'h859d, 16'h859e, 16'h859f 	:	val_out <= 16'h6e7b;
         16'h85a0, 16'h85a1, 16'h85a2, 16'h85a3, 16'h85a4, 16'h85a5, 16'h85a6, 16'h85a7 	:	val_out <= 16'h6e62;
         16'h85a8, 16'h85a9, 16'h85aa, 16'h85ab, 16'h85ac, 16'h85ad, 16'h85ae, 16'h85af 	:	val_out <= 16'h6e49;
         16'h85b0, 16'h85b1, 16'h85b2, 16'h85b3, 16'h85b4, 16'h85b5, 16'h85b6, 16'h85b7 	:	val_out <= 16'h6e30;
         16'h85b8, 16'h85b9, 16'h85ba, 16'h85bb, 16'h85bc, 16'h85bd, 16'h85be, 16'h85bf 	:	val_out <= 16'h6e17;
         16'h85c0, 16'h85c1, 16'h85c2, 16'h85c3, 16'h85c4, 16'h85c5, 16'h85c6, 16'h85c7 	:	val_out <= 16'h6dfe;
         16'h85c8, 16'h85c9, 16'h85ca, 16'h85cb, 16'h85cc, 16'h85cd, 16'h85ce, 16'h85cf 	:	val_out <= 16'h6de6;
         16'h85d0, 16'h85d1, 16'h85d2, 16'h85d3, 16'h85d4, 16'h85d5, 16'h85d6, 16'h85d7 	:	val_out <= 16'h6dcd;
         16'h85d8, 16'h85d9, 16'h85da, 16'h85db, 16'h85dc, 16'h85dd, 16'h85de, 16'h85df 	:	val_out <= 16'h6db4;
         16'h85e0, 16'h85e1, 16'h85e2, 16'h85e3, 16'h85e4, 16'h85e5, 16'h85e6, 16'h85e7 	:	val_out <= 16'h6d9b;
         16'h85e8, 16'h85e9, 16'h85ea, 16'h85eb, 16'h85ec, 16'h85ed, 16'h85ee, 16'h85ef 	:	val_out <= 16'h6d82;
         16'h85f0, 16'h85f1, 16'h85f2, 16'h85f3, 16'h85f4, 16'h85f5, 16'h85f6, 16'h85f7 	:	val_out <= 16'h6d69;
         16'h85f8, 16'h85f9, 16'h85fa, 16'h85fb, 16'h85fc, 16'h85fd, 16'h85fe, 16'h85ff 	:	val_out <= 16'h6d50;
         16'h8600, 16'h8601, 16'h8602, 16'h8603, 16'h8604, 16'h8605, 16'h8606, 16'h8607 	:	val_out <= 16'h6d37;
         16'h8608, 16'h8609, 16'h860a, 16'h860b, 16'h860c, 16'h860d, 16'h860e, 16'h860f 	:	val_out <= 16'h6d1f;
         16'h8610, 16'h8611, 16'h8612, 16'h8613, 16'h8614, 16'h8615, 16'h8616, 16'h8617 	:	val_out <= 16'h6d06;
         16'h8618, 16'h8619, 16'h861a, 16'h861b, 16'h861c, 16'h861d, 16'h861e, 16'h861f 	:	val_out <= 16'h6ced;
         16'h8620, 16'h8621, 16'h8622, 16'h8623, 16'h8624, 16'h8625, 16'h8626, 16'h8627 	:	val_out <= 16'h6cd4;
         16'h8628, 16'h8629, 16'h862a, 16'h862b, 16'h862c, 16'h862d, 16'h862e, 16'h862f 	:	val_out <= 16'h6cbb;
         16'h8630, 16'h8631, 16'h8632, 16'h8633, 16'h8634, 16'h8635, 16'h8636, 16'h8637 	:	val_out <= 16'h6ca2;
         16'h8638, 16'h8639, 16'h863a, 16'h863b, 16'h863c, 16'h863d, 16'h863e, 16'h863f 	:	val_out <= 16'h6c89;
         16'h8640, 16'h8641, 16'h8642, 16'h8643, 16'h8644, 16'h8645, 16'h8646, 16'h8647 	:	val_out <= 16'h6c71;
         16'h8648, 16'h8649, 16'h864a, 16'h864b, 16'h864c, 16'h864d, 16'h864e, 16'h864f 	:	val_out <= 16'h6c58;
         16'h8650, 16'h8651, 16'h8652, 16'h8653, 16'h8654, 16'h8655, 16'h8656, 16'h8657 	:	val_out <= 16'h6c3f;
         16'h8658, 16'h8659, 16'h865a, 16'h865b, 16'h865c, 16'h865d, 16'h865e, 16'h865f 	:	val_out <= 16'h6c26;
         16'h8660, 16'h8661, 16'h8662, 16'h8663, 16'h8664, 16'h8665, 16'h8666, 16'h8667 	:	val_out <= 16'h6c0d;
         16'h8668, 16'h8669, 16'h866a, 16'h866b, 16'h866c, 16'h866d, 16'h866e, 16'h866f 	:	val_out <= 16'h6bf4;
         16'h8670, 16'h8671, 16'h8672, 16'h8673, 16'h8674, 16'h8675, 16'h8676, 16'h8677 	:	val_out <= 16'h6bdc;
         16'h8678, 16'h8679, 16'h867a, 16'h867b, 16'h867c, 16'h867d, 16'h867e, 16'h867f 	:	val_out <= 16'h6bc3;
         16'h8680, 16'h8681, 16'h8682, 16'h8683, 16'h8684, 16'h8685, 16'h8686, 16'h8687 	:	val_out <= 16'h6baa;
         16'h8688, 16'h8689, 16'h868a, 16'h868b, 16'h868c, 16'h868d, 16'h868e, 16'h868f 	:	val_out <= 16'h6b91;
         16'h8690, 16'h8691, 16'h8692, 16'h8693, 16'h8694, 16'h8695, 16'h8696, 16'h8697 	:	val_out <= 16'h6b78;
         16'h8698, 16'h8699, 16'h869a, 16'h869b, 16'h869c, 16'h869d, 16'h869e, 16'h869f 	:	val_out <= 16'h6b60;
         16'h86a0, 16'h86a1, 16'h86a2, 16'h86a3, 16'h86a4, 16'h86a5, 16'h86a6, 16'h86a7 	:	val_out <= 16'h6b47;
         16'h86a8, 16'h86a9, 16'h86aa, 16'h86ab, 16'h86ac, 16'h86ad, 16'h86ae, 16'h86af 	:	val_out <= 16'h6b2e;
         16'h86b0, 16'h86b1, 16'h86b2, 16'h86b3, 16'h86b4, 16'h86b5, 16'h86b6, 16'h86b7 	:	val_out <= 16'h6b15;
         16'h86b8, 16'h86b9, 16'h86ba, 16'h86bb, 16'h86bc, 16'h86bd, 16'h86be, 16'h86bf 	:	val_out <= 16'h6afc;
         16'h86c0, 16'h86c1, 16'h86c2, 16'h86c3, 16'h86c4, 16'h86c5, 16'h86c6, 16'h86c7 	:	val_out <= 16'h6ae4;
         16'h86c8, 16'h86c9, 16'h86ca, 16'h86cb, 16'h86cc, 16'h86cd, 16'h86ce, 16'h86cf 	:	val_out <= 16'h6acb;
         16'h86d0, 16'h86d1, 16'h86d2, 16'h86d3, 16'h86d4, 16'h86d5, 16'h86d6, 16'h86d7 	:	val_out <= 16'h6ab2;
         16'h86d8, 16'h86d9, 16'h86da, 16'h86db, 16'h86dc, 16'h86dd, 16'h86de, 16'h86df 	:	val_out <= 16'h6a99;
         16'h86e0, 16'h86e1, 16'h86e2, 16'h86e3, 16'h86e4, 16'h86e5, 16'h86e6, 16'h86e7 	:	val_out <= 16'h6a80;
         16'h86e8, 16'h86e9, 16'h86ea, 16'h86eb, 16'h86ec, 16'h86ed, 16'h86ee, 16'h86ef 	:	val_out <= 16'h6a68;
         16'h86f0, 16'h86f1, 16'h86f2, 16'h86f3, 16'h86f4, 16'h86f5, 16'h86f6, 16'h86f7 	:	val_out <= 16'h6a4f;
         16'h86f8, 16'h86f9, 16'h86fa, 16'h86fb, 16'h86fc, 16'h86fd, 16'h86fe, 16'h86ff 	:	val_out <= 16'h6a36;
         16'h8700, 16'h8701, 16'h8702, 16'h8703, 16'h8704, 16'h8705, 16'h8706, 16'h8707 	:	val_out <= 16'h6a1d;
         16'h8708, 16'h8709, 16'h870a, 16'h870b, 16'h870c, 16'h870d, 16'h870e, 16'h870f 	:	val_out <= 16'h6a05;
         16'h8710, 16'h8711, 16'h8712, 16'h8713, 16'h8714, 16'h8715, 16'h8716, 16'h8717 	:	val_out <= 16'h69ec;
         16'h8718, 16'h8719, 16'h871a, 16'h871b, 16'h871c, 16'h871d, 16'h871e, 16'h871f 	:	val_out <= 16'h69d3;
         16'h8720, 16'h8721, 16'h8722, 16'h8723, 16'h8724, 16'h8725, 16'h8726, 16'h8727 	:	val_out <= 16'h69ba;
         16'h8728, 16'h8729, 16'h872a, 16'h872b, 16'h872c, 16'h872d, 16'h872e, 16'h872f 	:	val_out <= 16'h69a2;
         16'h8730, 16'h8731, 16'h8732, 16'h8733, 16'h8734, 16'h8735, 16'h8736, 16'h8737 	:	val_out <= 16'h6989;
         16'h8738, 16'h8739, 16'h873a, 16'h873b, 16'h873c, 16'h873d, 16'h873e, 16'h873f 	:	val_out <= 16'h6970;
         16'h8740, 16'h8741, 16'h8742, 16'h8743, 16'h8744, 16'h8745, 16'h8746, 16'h8747 	:	val_out <= 16'h6957;
         16'h8748, 16'h8749, 16'h874a, 16'h874b, 16'h874c, 16'h874d, 16'h874e, 16'h874f 	:	val_out <= 16'h693f;
         16'h8750, 16'h8751, 16'h8752, 16'h8753, 16'h8754, 16'h8755, 16'h8756, 16'h8757 	:	val_out <= 16'h6926;
         16'h8758, 16'h8759, 16'h875a, 16'h875b, 16'h875c, 16'h875d, 16'h875e, 16'h875f 	:	val_out <= 16'h690d;
         16'h8760, 16'h8761, 16'h8762, 16'h8763, 16'h8764, 16'h8765, 16'h8766, 16'h8767 	:	val_out <= 16'h68f5;
         16'h8768, 16'h8769, 16'h876a, 16'h876b, 16'h876c, 16'h876d, 16'h876e, 16'h876f 	:	val_out <= 16'h68dc;
         16'h8770, 16'h8771, 16'h8772, 16'h8773, 16'h8774, 16'h8775, 16'h8776, 16'h8777 	:	val_out <= 16'h68c3;
         16'h8778, 16'h8779, 16'h877a, 16'h877b, 16'h877c, 16'h877d, 16'h877e, 16'h877f 	:	val_out <= 16'h68aa;
         16'h8780, 16'h8781, 16'h8782, 16'h8783, 16'h8784, 16'h8785, 16'h8786, 16'h8787 	:	val_out <= 16'h6892;
         16'h8788, 16'h8789, 16'h878a, 16'h878b, 16'h878c, 16'h878d, 16'h878e, 16'h878f 	:	val_out <= 16'h6879;
         16'h8790, 16'h8791, 16'h8792, 16'h8793, 16'h8794, 16'h8795, 16'h8796, 16'h8797 	:	val_out <= 16'h6860;
         16'h8798, 16'h8799, 16'h879a, 16'h879b, 16'h879c, 16'h879d, 16'h879e, 16'h879f 	:	val_out <= 16'h6848;
         16'h87a0, 16'h87a1, 16'h87a2, 16'h87a3, 16'h87a4, 16'h87a5, 16'h87a6, 16'h87a7 	:	val_out <= 16'h682f;
         16'h87a8, 16'h87a9, 16'h87aa, 16'h87ab, 16'h87ac, 16'h87ad, 16'h87ae, 16'h87af 	:	val_out <= 16'h6816;
         16'h87b0, 16'h87b1, 16'h87b2, 16'h87b3, 16'h87b4, 16'h87b5, 16'h87b6, 16'h87b7 	:	val_out <= 16'h67fd;
         16'h87b8, 16'h87b9, 16'h87ba, 16'h87bb, 16'h87bc, 16'h87bd, 16'h87be, 16'h87bf 	:	val_out <= 16'h67e5;
         16'h87c0, 16'h87c1, 16'h87c2, 16'h87c3, 16'h87c4, 16'h87c5, 16'h87c6, 16'h87c7 	:	val_out <= 16'h67cc;
         16'h87c8, 16'h87c9, 16'h87ca, 16'h87cb, 16'h87cc, 16'h87cd, 16'h87ce, 16'h87cf 	:	val_out <= 16'h67b3;
         16'h87d0, 16'h87d1, 16'h87d2, 16'h87d3, 16'h87d4, 16'h87d5, 16'h87d6, 16'h87d7 	:	val_out <= 16'h679b;
         16'h87d8, 16'h87d9, 16'h87da, 16'h87db, 16'h87dc, 16'h87dd, 16'h87de, 16'h87df 	:	val_out <= 16'h6782;
         16'h87e0, 16'h87e1, 16'h87e2, 16'h87e3, 16'h87e4, 16'h87e5, 16'h87e6, 16'h87e7 	:	val_out <= 16'h6769;
         16'h87e8, 16'h87e9, 16'h87ea, 16'h87eb, 16'h87ec, 16'h87ed, 16'h87ee, 16'h87ef 	:	val_out <= 16'h6751;
         16'h87f0, 16'h87f1, 16'h87f2, 16'h87f3, 16'h87f4, 16'h87f5, 16'h87f6, 16'h87f7 	:	val_out <= 16'h6738;
         16'h87f8, 16'h87f9, 16'h87fa, 16'h87fb, 16'h87fc, 16'h87fd, 16'h87fe, 16'h87ff 	:	val_out <= 16'h671f;
         16'h8800, 16'h8801, 16'h8802, 16'h8803, 16'h8804, 16'h8805, 16'h8806, 16'h8807 	:	val_out <= 16'h6707;
         16'h8808, 16'h8809, 16'h880a, 16'h880b, 16'h880c, 16'h880d, 16'h880e, 16'h880f 	:	val_out <= 16'h66ee;
         16'h8810, 16'h8811, 16'h8812, 16'h8813, 16'h8814, 16'h8815, 16'h8816, 16'h8817 	:	val_out <= 16'h66d5;
         16'h8818, 16'h8819, 16'h881a, 16'h881b, 16'h881c, 16'h881d, 16'h881e, 16'h881f 	:	val_out <= 16'h66bd;
         16'h8820, 16'h8821, 16'h8822, 16'h8823, 16'h8824, 16'h8825, 16'h8826, 16'h8827 	:	val_out <= 16'h66a4;
         16'h8828, 16'h8829, 16'h882a, 16'h882b, 16'h882c, 16'h882d, 16'h882e, 16'h882f 	:	val_out <= 16'h668c;
         16'h8830, 16'h8831, 16'h8832, 16'h8833, 16'h8834, 16'h8835, 16'h8836, 16'h8837 	:	val_out <= 16'h6673;
         16'h8838, 16'h8839, 16'h883a, 16'h883b, 16'h883c, 16'h883d, 16'h883e, 16'h883f 	:	val_out <= 16'h665a;
         16'h8840, 16'h8841, 16'h8842, 16'h8843, 16'h8844, 16'h8845, 16'h8846, 16'h8847 	:	val_out <= 16'h6642;
         16'h8848, 16'h8849, 16'h884a, 16'h884b, 16'h884c, 16'h884d, 16'h884e, 16'h884f 	:	val_out <= 16'h6629;
         16'h8850, 16'h8851, 16'h8852, 16'h8853, 16'h8854, 16'h8855, 16'h8856, 16'h8857 	:	val_out <= 16'h6610;
         16'h8858, 16'h8859, 16'h885a, 16'h885b, 16'h885c, 16'h885d, 16'h885e, 16'h885f 	:	val_out <= 16'h65f8;
         16'h8860, 16'h8861, 16'h8862, 16'h8863, 16'h8864, 16'h8865, 16'h8866, 16'h8867 	:	val_out <= 16'h65df;
         16'h8868, 16'h8869, 16'h886a, 16'h886b, 16'h886c, 16'h886d, 16'h886e, 16'h886f 	:	val_out <= 16'h65c7;
         16'h8870, 16'h8871, 16'h8872, 16'h8873, 16'h8874, 16'h8875, 16'h8876, 16'h8877 	:	val_out <= 16'h65ae;
         16'h8878, 16'h8879, 16'h887a, 16'h887b, 16'h887c, 16'h887d, 16'h887e, 16'h887f 	:	val_out <= 16'h6595;
         16'h8880, 16'h8881, 16'h8882, 16'h8883, 16'h8884, 16'h8885, 16'h8886, 16'h8887 	:	val_out <= 16'h657d;
         16'h8888, 16'h8889, 16'h888a, 16'h888b, 16'h888c, 16'h888d, 16'h888e, 16'h888f 	:	val_out <= 16'h6564;
         16'h8890, 16'h8891, 16'h8892, 16'h8893, 16'h8894, 16'h8895, 16'h8896, 16'h8897 	:	val_out <= 16'h654c;
         16'h8898, 16'h8899, 16'h889a, 16'h889b, 16'h889c, 16'h889d, 16'h889e, 16'h889f 	:	val_out <= 16'h6533;
         16'h88a0, 16'h88a1, 16'h88a2, 16'h88a3, 16'h88a4, 16'h88a5, 16'h88a6, 16'h88a7 	:	val_out <= 16'h651b;
         16'h88a8, 16'h88a9, 16'h88aa, 16'h88ab, 16'h88ac, 16'h88ad, 16'h88ae, 16'h88af 	:	val_out <= 16'h6502;
         16'h88b0, 16'h88b1, 16'h88b2, 16'h88b3, 16'h88b4, 16'h88b5, 16'h88b6, 16'h88b7 	:	val_out <= 16'h64e9;
         16'h88b8, 16'h88b9, 16'h88ba, 16'h88bb, 16'h88bc, 16'h88bd, 16'h88be, 16'h88bf 	:	val_out <= 16'h64d1;
         16'h88c0, 16'h88c1, 16'h88c2, 16'h88c3, 16'h88c4, 16'h88c5, 16'h88c6, 16'h88c7 	:	val_out <= 16'h64b8;
         16'h88c8, 16'h88c9, 16'h88ca, 16'h88cb, 16'h88cc, 16'h88cd, 16'h88ce, 16'h88cf 	:	val_out <= 16'h64a0;
         16'h88d0, 16'h88d1, 16'h88d2, 16'h88d3, 16'h88d4, 16'h88d5, 16'h88d6, 16'h88d7 	:	val_out <= 16'h6487;
         16'h88d8, 16'h88d9, 16'h88da, 16'h88db, 16'h88dc, 16'h88dd, 16'h88de, 16'h88df 	:	val_out <= 16'h646f;
         16'h88e0, 16'h88e1, 16'h88e2, 16'h88e3, 16'h88e4, 16'h88e5, 16'h88e6, 16'h88e7 	:	val_out <= 16'h6456;
         16'h88e8, 16'h88e9, 16'h88ea, 16'h88eb, 16'h88ec, 16'h88ed, 16'h88ee, 16'h88ef 	:	val_out <= 16'h643e;
         16'h88f0, 16'h88f1, 16'h88f2, 16'h88f3, 16'h88f4, 16'h88f5, 16'h88f6, 16'h88f7 	:	val_out <= 16'h6425;
         16'h88f8, 16'h88f9, 16'h88fa, 16'h88fb, 16'h88fc, 16'h88fd, 16'h88fe, 16'h88ff 	:	val_out <= 16'h640d;
         16'h8900, 16'h8901, 16'h8902, 16'h8903, 16'h8904, 16'h8905, 16'h8906, 16'h8907 	:	val_out <= 16'h63f4;
         16'h8908, 16'h8909, 16'h890a, 16'h890b, 16'h890c, 16'h890d, 16'h890e, 16'h890f 	:	val_out <= 16'h63db;
         16'h8910, 16'h8911, 16'h8912, 16'h8913, 16'h8914, 16'h8915, 16'h8916, 16'h8917 	:	val_out <= 16'h63c3;
         16'h8918, 16'h8919, 16'h891a, 16'h891b, 16'h891c, 16'h891d, 16'h891e, 16'h891f 	:	val_out <= 16'h63aa;
         16'h8920, 16'h8921, 16'h8922, 16'h8923, 16'h8924, 16'h8925, 16'h8926, 16'h8927 	:	val_out <= 16'h6392;
         16'h8928, 16'h8929, 16'h892a, 16'h892b, 16'h892c, 16'h892d, 16'h892e, 16'h892f 	:	val_out <= 16'h6379;
         16'h8930, 16'h8931, 16'h8932, 16'h8933, 16'h8934, 16'h8935, 16'h8936, 16'h8937 	:	val_out <= 16'h6361;
         16'h8938, 16'h8939, 16'h893a, 16'h893b, 16'h893c, 16'h893d, 16'h893e, 16'h893f 	:	val_out <= 16'h6348;
         16'h8940, 16'h8941, 16'h8942, 16'h8943, 16'h8944, 16'h8945, 16'h8946, 16'h8947 	:	val_out <= 16'h6330;
         16'h8948, 16'h8949, 16'h894a, 16'h894b, 16'h894c, 16'h894d, 16'h894e, 16'h894f 	:	val_out <= 16'h6317;
         16'h8950, 16'h8951, 16'h8952, 16'h8953, 16'h8954, 16'h8955, 16'h8956, 16'h8957 	:	val_out <= 16'h62ff;
         16'h8958, 16'h8959, 16'h895a, 16'h895b, 16'h895c, 16'h895d, 16'h895e, 16'h895f 	:	val_out <= 16'h62e7;
         16'h8960, 16'h8961, 16'h8962, 16'h8963, 16'h8964, 16'h8965, 16'h8966, 16'h8967 	:	val_out <= 16'h62ce;
         16'h8968, 16'h8969, 16'h896a, 16'h896b, 16'h896c, 16'h896d, 16'h896e, 16'h896f 	:	val_out <= 16'h62b6;
         16'h8970, 16'h8971, 16'h8972, 16'h8973, 16'h8974, 16'h8975, 16'h8976, 16'h8977 	:	val_out <= 16'h629d;
         16'h8978, 16'h8979, 16'h897a, 16'h897b, 16'h897c, 16'h897d, 16'h897e, 16'h897f 	:	val_out <= 16'h6285;
         16'h8980, 16'h8981, 16'h8982, 16'h8983, 16'h8984, 16'h8985, 16'h8986, 16'h8987 	:	val_out <= 16'h626c;
         16'h8988, 16'h8989, 16'h898a, 16'h898b, 16'h898c, 16'h898d, 16'h898e, 16'h898f 	:	val_out <= 16'h6254;
         16'h8990, 16'h8991, 16'h8992, 16'h8993, 16'h8994, 16'h8995, 16'h8996, 16'h8997 	:	val_out <= 16'h623b;
         16'h8998, 16'h8999, 16'h899a, 16'h899b, 16'h899c, 16'h899d, 16'h899e, 16'h899f 	:	val_out <= 16'h6223;
         16'h89a0, 16'h89a1, 16'h89a2, 16'h89a3, 16'h89a4, 16'h89a5, 16'h89a6, 16'h89a7 	:	val_out <= 16'h620a;
         16'h89a8, 16'h89a9, 16'h89aa, 16'h89ab, 16'h89ac, 16'h89ad, 16'h89ae, 16'h89af 	:	val_out <= 16'h61f2;
         16'h89b0, 16'h89b1, 16'h89b2, 16'h89b3, 16'h89b4, 16'h89b5, 16'h89b6, 16'h89b7 	:	val_out <= 16'h61da;
         16'h89b8, 16'h89b9, 16'h89ba, 16'h89bb, 16'h89bc, 16'h89bd, 16'h89be, 16'h89bf 	:	val_out <= 16'h61c1;
         16'h89c0, 16'h89c1, 16'h89c2, 16'h89c3, 16'h89c4, 16'h89c5, 16'h89c6, 16'h89c7 	:	val_out <= 16'h61a9;
         16'h89c8, 16'h89c9, 16'h89ca, 16'h89cb, 16'h89cc, 16'h89cd, 16'h89ce, 16'h89cf 	:	val_out <= 16'h6190;
         16'h89d0, 16'h89d1, 16'h89d2, 16'h89d3, 16'h89d4, 16'h89d5, 16'h89d6, 16'h89d7 	:	val_out <= 16'h6178;
         16'h89d8, 16'h89d9, 16'h89da, 16'h89db, 16'h89dc, 16'h89dd, 16'h89de, 16'h89df 	:	val_out <= 16'h615f;
         16'h89e0, 16'h89e1, 16'h89e2, 16'h89e3, 16'h89e4, 16'h89e5, 16'h89e6, 16'h89e7 	:	val_out <= 16'h6147;
         16'h89e8, 16'h89e9, 16'h89ea, 16'h89eb, 16'h89ec, 16'h89ed, 16'h89ee, 16'h89ef 	:	val_out <= 16'h612f;
         16'h89f0, 16'h89f1, 16'h89f2, 16'h89f3, 16'h89f4, 16'h89f5, 16'h89f6, 16'h89f7 	:	val_out <= 16'h6116;
         16'h89f8, 16'h89f9, 16'h89fa, 16'h89fb, 16'h89fc, 16'h89fd, 16'h89fe, 16'h89ff 	:	val_out <= 16'h60fe;
         16'h8a00, 16'h8a01, 16'h8a02, 16'h8a03, 16'h8a04, 16'h8a05, 16'h8a06, 16'h8a07 	:	val_out <= 16'h60e6;
         16'h8a08, 16'h8a09, 16'h8a0a, 16'h8a0b, 16'h8a0c, 16'h8a0d, 16'h8a0e, 16'h8a0f 	:	val_out <= 16'h60cd;
         16'h8a10, 16'h8a11, 16'h8a12, 16'h8a13, 16'h8a14, 16'h8a15, 16'h8a16, 16'h8a17 	:	val_out <= 16'h60b5;
         16'h8a18, 16'h8a19, 16'h8a1a, 16'h8a1b, 16'h8a1c, 16'h8a1d, 16'h8a1e, 16'h8a1f 	:	val_out <= 16'h609c;
         16'h8a20, 16'h8a21, 16'h8a22, 16'h8a23, 16'h8a24, 16'h8a25, 16'h8a26, 16'h8a27 	:	val_out <= 16'h6084;
         16'h8a28, 16'h8a29, 16'h8a2a, 16'h8a2b, 16'h8a2c, 16'h8a2d, 16'h8a2e, 16'h8a2f 	:	val_out <= 16'h606c;
         16'h8a30, 16'h8a31, 16'h8a32, 16'h8a33, 16'h8a34, 16'h8a35, 16'h8a36, 16'h8a37 	:	val_out <= 16'h6053;
         16'h8a38, 16'h8a39, 16'h8a3a, 16'h8a3b, 16'h8a3c, 16'h8a3d, 16'h8a3e, 16'h8a3f 	:	val_out <= 16'h603b;
         16'h8a40, 16'h8a41, 16'h8a42, 16'h8a43, 16'h8a44, 16'h8a45, 16'h8a46, 16'h8a47 	:	val_out <= 16'h6023;
         16'h8a48, 16'h8a49, 16'h8a4a, 16'h8a4b, 16'h8a4c, 16'h8a4d, 16'h8a4e, 16'h8a4f 	:	val_out <= 16'h600a;
         16'h8a50, 16'h8a51, 16'h8a52, 16'h8a53, 16'h8a54, 16'h8a55, 16'h8a56, 16'h8a57 	:	val_out <= 16'h5ff2;
         16'h8a58, 16'h8a59, 16'h8a5a, 16'h8a5b, 16'h8a5c, 16'h8a5d, 16'h8a5e, 16'h8a5f 	:	val_out <= 16'h5fda;
         16'h8a60, 16'h8a61, 16'h8a62, 16'h8a63, 16'h8a64, 16'h8a65, 16'h8a66, 16'h8a67 	:	val_out <= 16'h5fc1;
         16'h8a68, 16'h8a69, 16'h8a6a, 16'h8a6b, 16'h8a6c, 16'h8a6d, 16'h8a6e, 16'h8a6f 	:	val_out <= 16'h5fa9;
         16'h8a70, 16'h8a71, 16'h8a72, 16'h8a73, 16'h8a74, 16'h8a75, 16'h8a76, 16'h8a77 	:	val_out <= 16'h5f91;
         16'h8a78, 16'h8a79, 16'h8a7a, 16'h8a7b, 16'h8a7c, 16'h8a7d, 16'h8a7e, 16'h8a7f 	:	val_out <= 16'h5f78;
         16'h8a80, 16'h8a81, 16'h8a82, 16'h8a83, 16'h8a84, 16'h8a85, 16'h8a86, 16'h8a87 	:	val_out <= 16'h5f60;
         16'h8a88, 16'h8a89, 16'h8a8a, 16'h8a8b, 16'h8a8c, 16'h8a8d, 16'h8a8e, 16'h8a8f 	:	val_out <= 16'h5f48;
         16'h8a90, 16'h8a91, 16'h8a92, 16'h8a93, 16'h8a94, 16'h8a95, 16'h8a96, 16'h8a97 	:	val_out <= 16'h5f2f;
         16'h8a98, 16'h8a99, 16'h8a9a, 16'h8a9b, 16'h8a9c, 16'h8a9d, 16'h8a9e, 16'h8a9f 	:	val_out <= 16'h5f17;
         16'h8aa0, 16'h8aa1, 16'h8aa2, 16'h8aa3, 16'h8aa4, 16'h8aa5, 16'h8aa6, 16'h8aa7 	:	val_out <= 16'h5eff;
         16'h8aa8, 16'h8aa9, 16'h8aaa, 16'h8aab, 16'h8aac, 16'h8aad, 16'h8aae, 16'h8aaf 	:	val_out <= 16'h5ee7;
         16'h8ab0, 16'h8ab1, 16'h8ab2, 16'h8ab3, 16'h8ab4, 16'h8ab5, 16'h8ab6, 16'h8ab7 	:	val_out <= 16'h5ece;
         16'h8ab8, 16'h8ab9, 16'h8aba, 16'h8abb, 16'h8abc, 16'h8abd, 16'h8abe, 16'h8abf 	:	val_out <= 16'h5eb6;
         16'h8ac0, 16'h8ac1, 16'h8ac2, 16'h8ac3, 16'h8ac4, 16'h8ac5, 16'h8ac6, 16'h8ac7 	:	val_out <= 16'h5e9e;
         16'h8ac8, 16'h8ac9, 16'h8aca, 16'h8acb, 16'h8acc, 16'h8acd, 16'h8ace, 16'h8acf 	:	val_out <= 16'h5e86;
         16'h8ad0, 16'h8ad1, 16'h8ad2, 16'h8ad3, 16'h8ad4, 16'h8ad5, 16'h8ad6, 16'h8ad7 	:	val_out <= 16'h5e6d;
         16'h8ad8, 16'h8ad9, 16'h8ada, 16'h8adb, 16'h8adc, 16'h8add, 16'h8ade, 16'h8adf 	:	val_out <= 16'h5e55;
         16'h8ae0, 16'h8ae1, 16'h8ae2, 16'h8ae3, 16'h8ae4, 16'h8ae5, 16'h8ae6, 16'h8ae7 	:	val_out <= 16'h5e3d;
         16'h8ae8, 16'h8ae9, 16'h8aea, 16'h8aeb, 16'h8aec, 16'h8aed, 16'h8aee, 16'h8aef 	:	val_out <= 16'h5e25;
         16'h8af0, 16'h8af1, 16'h8af2, 16'h8af3, 16'h8af4, 16'h8af5, 16'h8af6, 16'h8af7 	:	val_out <= 16'h5e0c;
         16'h8af8, 16'h8af9, 16'h8afa, 16'h8afb, 16'h8afc, 16'h8afd, 16'h8afe, 16'h8aff 	:	val_out <= 16'h5df4;
         16'h8b00, 16'h8b01, 16'h8b02, 16'h8b03, 16'h8b04, 16'h8b05, 16'h8b06, 16'h8b07 	:	val_out <= 16'h5ddc;
         16'h8b08, 16'h8b09, 16'h8b0a, 16'h8b0b, 16'h8b0c, 16'h8b0d, 16'h8b0e, 16'h8b0f 	:	val_out <= 16'h5dc4;
         16'h8b10, 16'h8b11, 16'h8b12, 16'h8b13, 16'h8b14, 16'h8b15, 16'h8b16, 16'h8b17 	:	val_out <= 16'h5dab;
         16'h8b18, 16'h8b19, 16'h8b1a, 16'h8b1b, 16'h8b1c, 16'h8b1d, 16'h8b1e, 16'h8b1f 	:	val_out <= 16'h5d93;
         16'h8b20, 16'h8b21, 16'h8b22, 16'h8b23, 16'h8b24, 16'h8b25, 16'h8b26, 16'h8b27 	:	val_out <= 16'h5d7b;
         16'h8b28, 16'h8b29, 16'h8b2a, 16'h8b2b, 16'h8b2c, 16'h8b2d, 16'h8b2e, 16'h8b2f 	:	val_out <= 16'h5d63;
         16'h8b30, 16'h8b31, 16'h8b32, 16'h8b33, 16'h8b34, 16'h8b35, 16'h8b36, 16'h8b37 	:	val_out <= 16'h5d4b;
         16'h8b38, 16'h8b39, 16'h8b3a, 16'h8b3b, 16'h8b3c, 16'h8b3d, 16'h8b3e, 16'h8b3f 	:	val_out <= 16'h5d32;
         16'h8b40, 16'h8b41, 16'h8b42, 16'h8b43, 16'h8b44, 16'h8b45, 16'h8b46, 16'h8b47 	:	val_out <= 16'h5d1a;
         16'h8b48, 16'h8b49, 16'h8b4a, 16'h8b4b, 16'h8b4c, 16'h8b4d, 16'h8b4e, 16'h8b4f 	:	val_out <= 16'h5d02;
         16'h8b50, 16'h8b51, 16'h8b52, 16'h8b53, 16'h8b54, 16'h8b55, 16'h8b56, 16'h8b57 	:	val_out <= 16'h5cea;
         16'h8b58, 16'h8b59, 16'h8b5a, 16'h8b5b, 16'h8b5c, 16'h8b5d, 16'h8b5e, 16'h8b5f 	:	val_out <= 16'h5cd2;
         16'h8b60, 16'h8b61, 16'h8b62, 16'h8b63, 16'h8b64, 16'h8b65, 16'h8b66, 16'h8b67 	:	val_out <= 16'h5cba;
         16'h8b68, 16'h8b69, 16'h8b6a, 16'h8b6b, 16'h8b6c, 16'h8b6d, 16'h8b6e, 16'h8b6f 	:	val_out <= 16'h5ca1;
         16'h8b70, 16'h8b71, 16'h8b72, 16'h8b73, 16'h8b74, 16'h8b75, 16'h8b76, 16'h8b77 	:	val_out <= 16'h5c89;
         16'h8b78, 16'h8b79, 16'h8b7a, 16'h8b7b, 16'h8b7c, 16'h8b7d, 16'h8b7e, 16'h8b7f 	:	val_out <= 16'h5c71;
         16'h8b80, 16'h8b81, 16'h8b82, 16'h8b83, 16'h8b84, 16'h8b85, 16'h8b86, 16'h8b87 	:	val_out <= 16'h5c59;
         16'h8b88, 16'h8b89, 16'h8b8a, 16'h8b8b, 16'h8b8c, 16'h8b8d, 16'h8b8e, 16'h8b8f 	:	val_out <= 16'h5c41;
         16'h8b90, 16'h8b91, 16'h8b92, 16'h8b93, 16'h8b94, 16'h8b95, 16'h8b96, 16'h8b97 	:	val_out <= 16'h5c29;
         16'h8b98, 16'h8b99, 16'h8b9a, 16'h8b9b, 16'h8b9c, 16'h8b9d, 16'h8b9e, 16'h8b9f 	:	val_out <= 16'h5c11;
         16'h8ba0, 16'h8ba1, 16'h8ba2, 16'h8ba3, 16'h8ba4, 16'h8ba5, 16'h8ba6, 16'h8ba7 	:	val_out <= 16'h5bf8;
         16'h8ba8, 16'h8ba9, 16'h8baa, 16'h8bab, 16'h8bac, 16'h8bad, 16'h8bae, 16'h8baf 	:	val_out <= 16'h5be0;
         16'h8bb0, 16'h8bb1, 16'h8bb2, 16'h8bb3, 16'h8bb4, 16'h8bb5, 16'h8bb6, 16'h8bb7 	:	val_out <= 16'h5bc8;
         16'h8bb8, 16'h8bb9, 16'h8bba, 16'h8bbb, 16'h8bbc, 16'h8bbd, 16'h8bbe, 16'h8bbf 	:	val_out <= 16'h5bb0;
         16'h8bc0, 16'h8bc1, 16'h8bc2, 16'h8bc3, 16'h8bc4, 16'h8bc5, 16'h8bc6, 16'h8bc7 	:	val_out <= 16'h5b98;
         16'h8bc8, 16'h8bc9, 16'h8bca, 16'h8bcb, 16'h8bcc, 16'h8bcd, 16'h8bce, 16'h8bcf 	:	val_out <= 16'h5b80;
         16'h8bd0, 16'h8bd1, 16'h8bd2, 16'h8bd3, 16'h8bd4, 16'h8bd5, 16'h8bd6, 16'h8bd7 	:	val_out <= 16'h5b68;
         16'h8bd8, 16'h8bd9, 16'h8bda, 16'h8bdb, 16'h8bdc, 16'h8bdd, 16'h8bde, 16'h8bdf 	:	val_out <= 16'h5b50;
         16'h8be0, 16'h8be1, 16'h8be2, 16'h8be3, 16'h8be4, 16'h8be5, 16'h8be6, 16'h8be7 	:	val_out <= 16'h5b38;
         16'h8be8, 16'h8be9, 16'h8bea, 16'h8beb, 16'h8bec, 16'h8bed, 16'h8bee, 16'h8bef 	:	val_out <= 16'h5b20;
         16'h8bf0, 16'h8bf1, 16'h8bf2, 16'h8bf3, 16'h8bf4, 16'h8bf5, 16'h8bf6, 16'h8bf7 	:	val_out <= 16'h5b08;
         16'h8bf8, 16'h8bf9, 16'h8bfa, 16'h8bfb, 16'h8bfc, 16'h8bfd, 16'h8bfe, 16'h8bff 	:	val_out <= 16'h5af0;
         16'h8c00, 16'h8c01, 16'h8c02, 16'h8c03, 16'h8c04, 16'h8c05, 16'h8c06, 16'h8c07 	:	val_out <= 16'h5ad7;
         16'h8c08, 16'h8c09, 16'h8c0a, 16'h8c0b, 16'h8c0c, 16'h8c0d, 16'h8c0e, 16'h8c0f 	:	val_out <= 16'h5abf;
         16'h8c10, 16'h8c11, 16'h8c12, 16'h8c13, 16'h8c14, 16'h8c15, 16'h8c16, 16'h8c17 	:	val_out <= 16'h5aa7;
         16'h8c18, 16'h8c19, 16'h8c1a, 16'h8c1b, 16'h8c1c, 16'h8c1d, 16'h8c1e, 16'h8c1f 	:	val_out <= 16'h5a8f;
         16'h8c20, 16'h8c21, 16'h8c22, 16'h8c23, 16'h8c24, 16'h8c25, 16'h8c26, 16'h8c27 	:	val_out <= 16'h5a77;
         16'h8c28, 16'h8c29, 16'h8c2a, 16'h8c2b, 16'h8c2c, 16'h8c2d, 16'h8c2e, 16'h8c2f 	:	val_out <= 16'h5a5f;
         16'h8c30, 16'h8c31, 16'h8c32, 16'h8c33, 16'h8c34, 16'h8c35, 16'h8c36, 16'h8c37 	:	val_out <= 16'h5a47;
         16'h8c38, 16'h8c39, 16'h8c3a, 16'h8c3b, 16'h8c3c, 16'h8c3d, 16'h8c3e, 16'h8c3f 	:	val_out <= 16'h5a2f;
         16'h8c40, 16'h8c41, 16'h8c42, 16'h8c43, 16'h8c44, 16'h8c45, 16'h8c46, 16'h8c47 	:	val_out <= 16'h5a17;
         16'h8c48, 16'h8c49, 16'h8c4a, 16'h8c4b, 16'h8c4c, 16'h8c4d, 16'h8c4e, 16'h8c4f 	:	val_out <= 16'h59ff;
         16'h8c50, 16'h8c51, 16'h8c52, 16'h8c53, 16'h8c54, 16'h8c55, 16'h8c56, 16'h8c57 	:	val_out <= 16'h59e7;
         16'h8c58, 16'h8c59, 16'h8c5a, 16'h8c5b, 16'h8c5c, 16'h8c5d, 16'h8c5e, 16'h8c5f 	:	val_out <= 16'h59cf;
         16'h8c60, 16'h8c61, 16'h8c62, 16'h8c63, 16'h8c64, 16'h8c65, 16'h8c66, 16'h8c67 	:	val_out <= 16'h59b7;
         16'h8c68, 16'h8c69, 16'h8c6a, 16'h8c6b, 16'h8c6c, 16'h8c6d, 16'h8c6e, 16'h8c6f 	:	val_out <= 16'h599f;
         16'h8c70, 16'h8c71, 16'h8c72, 16'h8c73, 16'h8c74, 16'h8c75, 16'h8c76, 16'h8c77 	:	val_out <= 16'h5987;
         16'h8c78, 16'h8c79, 16'h8c7a, 16'h8c7b, 16'h8c7c, 16'h8c7d, 16'h8c7e, 16'h8c7f 	:	val_out <= 16'h596f;
         16'h8c80, 16'h8c81, 16'h8c82, 16'h8c83, 16'h8c84, 16'h8c85, 16'h8c86, 16'h8c87 	:	val_out <= 16'h5957;
         16'h8c88, 16'h8c89, 16'h8c8a, 16'h8c8b, 16'h8c8c, 16'h8c8d, 16'h8c8e, 16'h8c8f 	:	val_out <= 16'h593f;
         16'h8c90, 16'h8c91, 16'h8c92, 16'h8c93, 16'h8c94, 16'h8c95, 16'h8c96, 16'h8c97 	:	val_out <= 16'h5927;
         16'h8c98, 16'h8c99, 16'h8c9a, 16'h8c9b, 16'h8c9c, 16'h8c9d, 16'h8c9e, 16'h8c9f 	:	val_out <= 16'h5910;
         16'h8ca0, 16'h8ca1, 16'h8ca2, 16'h8ca3, 16'h8ca4, 16'h8ca5, 16'h8ca6, 16'h8ca7 	:	val_out <= 16'h58f8;
         16'h8ca8, 16'h8ca9, 16'h8caa, 16'h8cab, 16'h8cac, 16'h8cad, 16'h8cae, 16'h8caf 	:	val_out <= 16'h58e0;
         16'h8cb0, 16'h8cb1, 16'h8cb2, 16'h8cb3, 16'h8cb4, 16'h8cb5, 16'h8cb6, 16'h8cb7 	:	val_out <= 16'h58c8;
         16'h8cb8, 16'h8cb9, 16'h8cba, 16'h8cbb, 16'h8cbc, 16'h8cbd, 16'h8cbe, 16'h8cbf 	:	val_out <= 16'h58b0;
         16'h8cc0, 16'h8cc1, 16'h8cc2, 16'h8cc3, 16'h8cc4, 16'h8cc5, 16'h8cc6, 16'h8cc7 	:	val_out <= 16'h5898;
         16'h8cc8, 16'h8cc9, 16'h8cca, 16'h8ccb, 16'h8ccc, 16'h8ccd, 16'h8cce, 16'h8ccf 	:	val_out <= 16'h5880;
         16'h8cd0, 16'h8cd1, 16'h8cd2, 16'h8cd3, 16'h8cd4, 16'h8cd5, 16'h8cd6, 16'h8cd7 	:	val_out <= 16'h5868;
         16'h8cd8, 16'h8cd9, 16'h8cda, 16'h8cdb, 16'h8cdc, 16'h8cdd, 16'h8cde, 16'h8cdf 	:	val_out <= 16'h5850;
         16'h8ce0, 16'h8ce1, 16'h8ce2, 16'h8ce3, 16'h8ce4, 16'h8ce5, 16'h8ce6, 16'h8ce7 	:	val_out <= 16'h5838;
         16'h8ce8, 16'h8ce9, 16'h8cea, 16'h8ceb, 16'h8cec, 16'h8ced, 16'h8cee, 16'h8cef 	:	val_out <= 16'h5820;
         16'h8cf0, 16'h8cf1, 16'h8cf2, 16'h8cf3, 16'h8cf4, 16'h8cf5, 16'h8cf6, 16'h8cf7 	:	val_out <= 16'h5809;
         16'h8cf8, 16'h8cf9, 16'h8cfa, 16'h8cfb, 16'h8cfc, 16'h8cfd, 16'h8cfe, 16'h8cff 	:	val_out <= 16'h57f1;
         16'h8d00, 16'h8d01, 16'h8d02, 16'h8d03, 16'h8d04, 16'h8d05, 16'h8d06, 16'h8d07 	:	val_out <= 16'h57d9;
         16'h8d08, 16'h8d09, 16'h8d0a, 16'h8d0b, 16'h8d0c, 16'h8d0d, 16'h8d0e, 16'h8d0f 	:	val_out <= 16'h57c1;
         16'h8d10, 16'h8d11, 16'h8d12, 16'h8d13, 16'h8d14, 16'h8d15, 16'h8d16, 16'h8d17 	:	val_out <= 16'h57a9;
         16'h8d18, 16'h8d19, 16'h8d1a, 16'h8d1b, 16'h8d1c, 16'h8d1d, 16'h8d1e, 16'h8d1f 	:	val_out <= 16'h5791;
         16'h8d20, 16'h8d21, 16'h8d22, 16'h8d23, 16'h8d24, 16'h8d25, 16'h8d26, 16'h8d27 	:	val_out <= 16'h5779;
         16'h8d28, 16'h8d29, 16'h8d2a, 16'h8d2b, 16'h8d2c, 16'h8d2d, 16'h8d2e, 16'h8d2f 	:	val_out <= 16'h5762;
         16'h8d30, 16'h8d31, 16'h8d32, 16'h8d33, 16'h8d34, 16'h8d35, 16'h8d36, 16'h8d37 	:	val_out <= 16'h574a;
         16'h8d38, 16'h8d39, 16'h8d3a, 16'h8d3b, 16'h8d3c, 16'h8d3d, 16'h8d3e, 16'h8d3f 	:	val_out <= 16'h5732;
         16'h8d40, 16'h8d41, 16'h8d42, 16'h8d43, 16'h8d44, 16'h8d45, 16'h8d46, 16'h8d47 	:	val_out <= 16'h571a;
         16'h8d48, 16'h8d49, 16'h8d4a, 16'h8d4b, 16'h8d4c, 16'h8d4d, 16'h8d4e, 16'h8d4f 	:	val_out <= 16'h5702;
         16'h8d50, 16'h8d51, 16'h8d52, 16'h8d53, 16'h8d54, 16'h8d55, 16'h8d56, 16'h8d57 	:	val_out <= 16'h56ea;
         16'h8d58, 16'h8d59, 16'h8d5a, 16'h8d5b, 16'h8d5c, 16'h8d5d, 16'h8d5e, 16'h8d5f 	:	val_out <= 16'h56d3;
         16'h8d60, 16'h8d61, 16'h8d62, 16'h8d63, 16'h8d64, 16'h8d65, 16'h8d66, 16'h8d67 	:	val_out <= 16'h56bb;
         16'h8d68, 16'h8d69, 16'h8d6a, 16'h8d6b, 16'h8d6c, 16'h8d6d, 16'h8d6e, 16'h8d6f 	:	val_out <= 16'h56a3;
         16'h8d70, 16'h8d71, 16'h8d72, 16'h8d73, 16'h8d74, 16'h8d75, 16'h8d76, 16'h8d77 	:	val_out <= 16'h568b;
         16'h8d78, 16'h8d79, 16'h8d7a, 16'h8d7b, 16'h8d7c, 16'h8d7d, 16'h8d7e, 16'h8d7f 	:	val_out <= 16'h5674;
         16'h8d80, 16'h8d81, 16'h8d82, 16'h8d83, 16'h8d84, 16'h8d85, 16'h8d86, 16'h8d87 	:	val_out <= 16'h565c;
         16'h8d88, 16'h8d89, 16'h8d8a, 16'h8d8b, 16'h8d8c, 16'h8d8d, 16'h8d8e, 16'h8d8f 	:	val_out <= 16'h5644;
         16'h8d90, 16'h8d91, 16'h8d92, 16'h8d93, 16'h8d94, 16'h8d95, 16'h8d96, 16'h8d97 	:	val_out <= 16'h562c;
         16'h8d98, 16'h8d99, 16'h8d9a, 16'h8d9b, 16'h8d9c, 16'h8d9d, 16'h8d9e, 16'h8d9f 	:	val_out <= 16'h5614;
         16'h8da0, 16'h8da1, 16'h8da2, 16'h8da3, 16'h8da4, 16'h8da5, 16'h8da6, 16'h8da7 	:	val_out <= 16'h55fd;
         16'h8da8, 16'h8da9, 16'h8daa, 16'h8dab, 16'h8dac, 16'h8dad, 16'h8dae, 16'h8daf 	:	val_out <= 16'h55e5;
         16'h8db0, 16'h8db1, 16'h8db2, 16'h8db3, 16'h8db4, 16'h8db5, 16'h8db6, 16'h8db7 	:	val_out <= 16'h55cd;
         16'h8db8, 16'h8db9, 16'h8dba, 16'h8dbb, 16'h8dbc, 16'h8dbd, 16'h8dbe, 16'h8dbf 	:	val_out <= 16'h55b6;
         16'h8dc0, 16'h8dc1, 16'h8dc2, 16'h8dc3, 16'h8dc4, 16'h8dc5, 16'h8dc6, 16'h8dc7 	:	val_out <= 16'h559e;
         16'h8dc8, 16'h8dc9, 16'h8dca, 16'h8dcb, 16'h8dcc, 16'h8dcd, 16'h8dce, 16'h8dcf 	:	val_out <= 16'h5586;
         16'h8dd0, 16'h8dd1, 16'h8dd2, 16'h8dd3, 16'h8dd4, 16'h8dd5, 16'h8dd6, 16'h8dd7 	:	val_out <= 16'h556e;
         16'h8dd8, 16'h8dd9, 16'h8dda, 16'h8ddb, 16'h8ddc, 16'h8ddd, 16'h8dde, 16'h8ddf 	:	val_out <= 16'h5557;
         16'h8de0, 16'h8de1, 16'h8de2, 16'h8de3, 16'h8de4, 16'h8de5, 16'h8de6, 16'h8de7 	:	val_out <= 16'h553f;
         16'h8de8, 16'h8de9, 16'h8dea, 16'h8deb, 16'h8dec, 16'h8ded, 16'h8dee, 16'h8def 	:	val_out <= 16'h5527;
         16'h8df0, 16'h8df1, 16'h8df2, 16'h8df3, 16'h8df4, 16'h8df5, 16'h8df6, 16'h8df7 	:	val_out <= 16'h5510;
         16'h8df8, 16'h8df9, 16'h8dfa, 16'h8dfb, 16'h8dfc, 16'h8dfd, 16'h8dfe, 16'h8dff 	:	val_out <= 16'h54f8;
         16'h8e00, 16'h8e01, 16'h8e02, 16'h8e03, 16'h8e04, 16'h8e05, 16'h8e06, 16'h8e07 	:	val_out <= 16'h54e0;
         16'h8e08, 16'h8e09, 16'h8e0a, 16'h8e0b, 16'h8e0c, 16'h8e0d, 16'h8e0e, 16'h8e0f 	:	val_out <= 16'h54c9;
         16'h8e10, 16'h8e11, 16'h8e12, 16'h8e13, 16'h8e14, 16'h8e15, 16'h8e16, 16'h8e17 	:	val_out <= 16'h54b1;
         16'h8e18, 16'h8e19, 16'h8e1a, 16'h8e1b, 16'h8e1c, 16'h8e1d, 16'h8e1e, 16'h8e1f 	:	val_out <= 16'h5499;
         16'h8e20, 16'h8e21, 16'h8e22, 16'h8e23, 16'h8e24, 16'h8e25, 16'h8e26, 16'h8e27 	:	val_out <= 16'h5482;
         16'h8e28, 16'h8e29, 16'h8e2a, 16'h8e2b, 16'h8e2c, 16'h8e2d, 16'h8e2e, 16'h8e2f 	:	val_out <= 16'h546a;
         16'h8e30, 16'h8e31, 16'h8e32, 16'h8e33, 16'h8e34, 16'h8e35, 16'h8e36, 16'h8e37 	:	val_out <= 16'h5452;
         16'h8e38, 16'h8e39, 16'h8e3a, 16'h8e3b, 16'h8e3c, 16'h8e3d, 16'h8e3e, 16'h8e3f 	:	val_out <= 16'h543b;
         16'h8e40, 16'h8e41, 16'h8e42, 16'h8e43, 16'h8e44, 16'h8e45, 16'h8e46, 16'h8e47 	:	val_out <= 16'h5423;
         16'h8e48, 16'h8e49, 16'h8e4a, 16'h8e4b, 16'h8e4c, 16'h8e4d, 16'h8e4e, 16'h8e4f 	:	val_out <= 16'h540c;
         16'h8e50, 16'h8e51, 16'h8e52, 16'h8e53, 16'h8e54, 16'h8e55, 16'h8e56, 16'h8e57 	:	val_out <= 16'h53f4;
         16'h8e58, 16'h8e59, 16'h8e5a, 16'h8e5b, 16'h8e5c, 16'h8e5d, 16'h8e5e, 16'h8e5f 	:	val_out <= 16'h53dc;
         16'h8e60, 16'h8e61, 16'h8e62, 16'h8e63, 16'h8e64, 16'h8e65, 16'h8e66, 16'h8e67 	:	val_out <= 16'h53c5;
         16'h8e68, 16'h8e69, 16'h8e6a, 16'h8e6b, 16'h8e6c, 16'h8e6d, 16'h8e6e, 16'h8e6f 	:	val_out <= 16'h53ad;
         16'h8e70, 16'h8e71, 16'h8e72, 16'h8e73, 16'h8e74, 16'h8e75, 16'h8e76, 16'h8e77 	:	val_out <= 16'h5396;
         16'h8e78, 16'h8e79, 16'h8e7a, 16'h8e7b, 16'h8e7c, 16'h8e7d, 16'h8e7e, 16'h8e7f 	:	val_out <= 16'h537e;
         16'h8e80, 16'h8e81, 16'h8e82, 16'h8e83, 16'h8e84, 16'h8e85, 16'h8e86, 16'h8e87 	:	val_out <= 16'h5367;
         16'h8e88, 16'h8e89, 16'h8e8a, 16'h8e8b, 16'h8e8c, 16'h8e8d, 16'h8e8e, 16'h8e8f 	:	val_out <= 16'h534f;
         16'h8e90, 16'h8e91, 16'h8e92, 16'h8e93, 16'h8e94, 16'h8e95, 16'h8e96, 16'h8e97 	:	val_out <= 16'h5337;
         16'h8e98, 16'h8e99, 16'h8e9a, 16'h8e9b, 16'h8e9c, 16'h8e9d, 16'h8e9e, 16'h8e9f 	:	val_out <= 16'h5320;
         16'h8ea0, 16'h8ea1, 16'h8ea2, 16'h8ea3, 16'h8ea4, 16'h8ea5, 16'h8ea6, 16'h8ea7 	:	val_out <= 16'h5308;
         16'h8ea8, 16'h8ea9, 16'h8eaa, 16'h8eab, 16'h8eac, 16'h8ead, 16'h8eae, 16'h8eaf 	:	val_out <= 16'h52f1;
         16'h8eb0, 16'h8eb1, 16'h8eb2, 16'h8eb3, 16'h8eb4, 16'h8eb5, 16'h8eb6, 16'h8eb7 	:	val_out <= 16'h52d9;
         16'h8eb8, 16'h8eb9, 16'h8eba, 16'h8ebb, 16'h8ebc, 16'h8ebd, 16'h8ebe, 16'h8ebf 	:	val_out <= 16'h52c2;
         16'h8ec0, 16'h8ec1, 16'h8ec2, 16'h8ec3, 16'h8ec4, 16'h8ec5, 16'h8ec6, 16'h8ec7 	:	val_out <= 16'h52aa;
         16'h8ec8, 16'h8ec9, 16'h8eca, 16'h8ecb, 16'h8ecc, 16'h8ecd, 16'h8ece, 16'h8ecf 	:	val_out <= 16'h5293;
         16'h8ed0, 16'h8ed1, 16'h8ed2, 16'h8ed3, 16'h8ed4, 16'h8ed5, 16'h8ed6, 16'h8ed7 	:	val_out <= 16'h527b;
         16'h8ed8, 16'h8ed9, 16'h8eda, 16'h8edb, 16'h8edc, 16'h8edd, 16'h8ede, 16'h8edf 	:	val_out <= 16'h5264;
         16'h8ee0, 16'h8ee1, 16'h8ee2, 16'h8ee3, 16'h8ee4, 16'h8ee5, 16'h8ee6, 16'h8ee7 	:	val_out <= 16'h524c;
         16'h8ee8, 16'h8ee9, 16'h8eea, 16'h8eeb, 16'h8eec, 16'h8eed, 16'h8eee, 16'h8eef 	:	val_out <= 16'h5235;
         16'h8ef0, 16'h8ef1, 16'h8ef2, 16'h8ef3, 16'h8ef4, 16'h8ef5, 16'h8ef6, 16'h8ef7 	:	val_out <= 16'h521d;
         16'h8ef8, 16'h8ef9, 16'h8efa, 16'h8efb, 16'h8efc, 16'h8efd, 16'h8efe, 16'h8eff 	:	val_out <= 16'h5206;
         16'h8f00, 16'h8f01, 16'h8f02, 16'h8f03, 16'h8f04, 16'h8f05, 16'h8f06, 16'h8f07 	:	val_out <= 16'h51ee;
         16'h8f08, 16'h8f09, 16'h8f0a, 16'h8f0b, 16'h8f0c, 16'h8f0d, 16'h8f0e, 16'h8f0f 	:	val_out <= 16'h51d7;
         16'h8f10, 16'h8f11, 16'h8f12, 16'h8f13, 16'h8f14, 16'h8f15, 16'h8f16, 16'h8f17 	:	val_out <= 16'h51c0;
         16'h8f18, 16'h8f19, 16'h8f1a, 16'h8f1b, 16'h8f1c, 16'h8f1d, 16'h8f1e, 16'h8f1f 	:	val_out <= 16'h51a8;
         16'h8f20, 16'h8f21, 16'h8f22, 16'h8f23, 16'h8f24, 16'h8f25, 16'h8f26, 16'h8f27 	:	val_out <= 16'h5191;
         16'h8f28, 16'h8f29, 16'h8f2a, 16'h8f2b, 16'h8f2c, 16'h8f2d, 16'h8f2e, 16'h8f2f 	:	val_out <= 16'h5179;
         16'h8f30, 16'h8f31, 16'h8f32, 16'h8f33, 16'h8f34, 16'h8f35, 16'h8f36, 16'h8f37 	:	val_out <= 16'h5162;
         16'h8f38, 16'h8f39, 16'h8f3a, 16'h8f3b, 16'h8f3c, 16'h8f3d, 16'h8f3e, 16'h8f3f 	:	val_out <= 16'h514a;
         16'h8f40, 16'h8f41, 16'h8f42, 16'h8f43, 16'h8f44, 16'h8f45, 16'h8f46, 16'h8f47 	:	val_out <= 16'h5133;
         16'h8f48, 16'h8f49, 16'h8f4a, 16'h8f4b, 16'h8f4c, 16'h8f4d, 16'h8f4e, 16'h8f4f 	:	val_out <= 16'h511c;
         16'h8f50, 16'h8f51, 16'h8f52, 16'h8f53, 16'h8f54, 16'h8f55, 16'h8f56, 16'h8f57 	:	val_out <= 16'h5104;
         16'h8f58, 16'h8f59, 16'h8f5a, 16'h8f5b, 16'h8f5c, 16'h8f5d, 16'h8f5e, 16'h8f5f 	:	val_out <= 16'h50ed;
         16'h8f60, 16'h8f61, 16'h8f62, 16'h8f63, 16'h8f64, 16'h8f65, 16'h8f66, 16'h8f67 	:	val_out <= 16'h50d6;
         16'h8f68, 16'h8f69, 16'h8f6a, 16'h8f6b, 16'h8f6c, 16'h8f6d, 16'h8f6e, 16'h8f6f 	:	val_out <= 16'h50be;
         16'h8f70, 16'h8f71, 16'h8f72, 16'h8f73, 16'h8f74, 16'h8f75, 16'h8f76, 16'h8f77 	:	val_out <= 16'h50a7;
         16'h8f78, 16'h8f79, 16'h8f7a, 16'h8f7b, 16'h8f7c, 16'h8f7d, 16'h8f7e, 16'h8f7f 	:	val_out <= 16'h5090;
         16'h8f80, 16'h8f81, 16'h8f82, 16'h8f83, 16'h8f84, 16'h8f85, 16'h8f86, 16'h8f87 	:	val_out <= 16'h5078;
         16'h8f88, 16'h8f89, 16'h8f8a, 16'h8f8b, 16'h8f8c, 16'h8f8d, 16'h8f8e, 16'h8f8f 	:	val_out <= 16'h5061;
         16'h8f90, 16'h8f91, 16'h8f92, 16'h8f93, 16'h8f94, 16'h8f95, 16'h8f96, 16'h8f97 	:	val_out <= 16'h504a;
         16'h8f98, 16'h8f99, 16'h8f9a, 16'h8f9b, 16'h8f9c, 16'h8f9d, 16'h8f9e, 16'h8f9f 	:	val_out <= 16'h5032;
         16'h8fa0, 16'h8fa1, 16'h8fa2, 16'h8fa3, 16'h8fa4, 16'h8fa5, 16'h8fa6, 16'h8fa7 	:	val_out <= 16'h501b;
         16'h8fa8, 16'h8fa9, 16'h8faa, 16'h8fab, 16'h8fac, 16'h8fad, 16'h8fae, 16'h8faf 	:	val_out <= 16'h5004;
         16'h8fb0, 16'h8fb1, 16'h8fb2, 16'h8fb3, 16'h8fb4, 16'h8fb5, 16'h8fb6, 16'h8fb7 	:	val_out <= 16'h4fec;
         16'h8fb8, 16'h8fb9, 16'h8fba, 16'h8fbb, 16'h8fbc, 16'h8fbd, 16'h8fbe, 16'h8fbf 	:	val_out <= 16'h4fd5;
         16'h8fc0, 16'h8fc1, 16'h8fc2, 16'h8fc3, 16'h8fc4, 16'h8fc5, 16'h8fc6, 16'h8fc7 	:	val_out <= 16'h4fbe;
         16'h8fc8, 16'h8fc9, 16'h8fca, 16'h8fcb, 16'h8fcc, 16'h8fcd, 16'h8fce, 16'h8fcf 	:	val_out <= 16'h4fa6;
         16'h8fd0, 16'h8fd1, 16'h8fd2, 16'h8fd3, 16'h8fd4, 16'h8fd5, 16'h8fd6, 16'h8fd7 	:	val_out <= 16'h4f8f;
         16'h8fd8, 16'h8fd9, 16'h8fda, 16'h8fdb, 16'h8fdc, 16'h8fdd, 16'h8fde, 16'h8fdf 	:	val_out <= 16'h4f78;
         16'h8fe0, 16'h8fe1, 16'h8fe2, 16'h8fe3, 16'h8fe4, 16'h8fe5, 16'h8fe6, 16'h8fe7 	:	val_out <= 16'h4f61;
         16'h8fe8, 16'h8fe9, 16'h8fea, 16'h8feb, 16'h8fec, 16'h8fed, 16'h8fee, 16'h8fef 	:	val_out <= 16'h4f49;
         16'h8ff0, 16'h8ff1, 16'h8ff2, 16'h8ff3, 16'h8ff4, 16'h8ff5, 16'h8ff6, 16'h8ff7 	:	val_out <= 16'h4f32;
         16'h8ff8, 16'h8ff9, 16'h8ffa, 16'h8ffb, 16'h8ffc, 16'h8ffd, 16'h8ffe, 16'h8fff 	:	val_out <= 16'h4f1b;
         16'h9000, 16'h9001, 16'h9002, 16'h9003, 16'h9004, 16'h9005, 16'h9006, 16'h9007 	:	val_out <= 16'h4f04;
         16'h9008, 16'h9009, 16'h900a, 16'h900b, 16'h900c, 16'h900d, 16'h900e, 16'h900f 	:	val_out <= 16'h4eed;
         16'h9010, 16'h9011, 16'h9012, 16'h9013, 16'h9014, 16'h9015, 16'h9016, 16'h9017 	:	val_out <= 16'h4ed5;
         16'h9018, 16'h9019, 16'h901a, 16'h901b, 16'h901c, 16'h901d, 16'h901e, 16'h901f 	:	val_out <= 16'h4ebe;
         16'h9020, 16'h9021, 16'h9022, 16'h9023, 16'h9024, 16'h9025, 16'h9026, 16'h9027 	:	val_out <= 16'h4ea7;
         16'h9028, 16'h9029, 16'h902a, 16'h902b, 16'h902c, 16'h902d, 16'h902e, 16'h902f 	:	val_out <= 16'h4e90;
         16'h9030, 16'h9031, 16'h9032, 16'h9033, 16'h9034, 16'h9035, 16'h9036, 16'h9037 	:	val_out <= 16'h4e79;
         16'h9038, 16'h9039, 16'h903a, 16'h903b, 16'h903c, 16'h903d, 16'h903e, 16'h903f 	:	val_out <= 16'h4e61;
         16'h9040, 16'h9041, 16'h9042, 16'h9043, 16'h9044, 16'h9045, 16'h9046, 16'h9047 	:	val_out <= 16'h4e4a;
         16'h9048, 16'h9049, 16'h904a, 16'h904b, 16'h904c, 16'h904d, 16'h904e, 16'h904f 	:	val_out <= 16'h4e33;
         16'h9050, 16'h9051, 16'h9052, 16'h9053, 16'h9054, 16'h9055, 16'h9056, 16'h9057 	:	val_out <= 16'h4e1c;
         16'h9058, 16'h9059, 16'h905a, 16'h905b, 16'h905c, 16'h905d, 16'h905e, 16'h905f 	:	val_out <= 16'h4e05;
         16'h9060, 16'h9061, 16'h9062, 16'h9063, 16'h9064, 16'h9065, 16'h9066, 16'h9067 	:	val_out <= 16'h4dee;
         16'h9068, 16'h9069, 16'h906a, 16'h906b, 16'h906c, 16'h906d, 16'h906e, 16'h906f 	:	val_out <= 16'h4dd7;
         16'h9070, 16'h9071, 16'h9072, 16'h9073, 16'h9074, 16'h9075, 16'h9076, 16'h9077 	:	val_out <= 16'h4dbf;
         16'h9078, 16'h9079, 16'h907a, 16'h907b, 16'h907c, 16'h907d, 16'h907e, 16'h907f 	:	val_out <= 16'h4da8;
         16'h9080, 16'h9081, 16'h9082, 16'h9083, 16'h9084, 16'h9085, 16'h9086, 16'h9087 	:	val_out <= 16'h4d91;
         16'h9088, 16'h9089, 16'h908a, 16'h908b, 16'h908c, 16'h908d, 16'h908e, 16'h908f 	:	val_out <= 16'h4d7a;
         16'h9090, 16'h9091, 16'h9092, 16'h9093, 16'h9094, 16'h9095, 16'h9096, 16'h9097 	:	val_out <= 16'h4d63;
         16'h9098, 16'h9099, 16'h909a, 16'h909b, 16'h909c, 16'h909d, 16'h909e, 16'h909f 	:	val_out <= 16'h4d4c;
         16'h90a0, 16'h90a1, 16'h90a2, 16'h90a3, 16'h90a4, 16'h90a5, 16'h90a6, 16'h90a7 	:	val_out <= 16'h4d35;
         16'h90a8, 16'h90a9, 16'h90aa, 16'h90ab, 16'h90ac, 16'h90ad, 16'h90ae, 16'h90af 	:	val_out <= 16'h4d1e;
         16'h90b0, 16'h90b1, 16'h90b2, 16'h90b3, 16'h90b4, 16'h90b5, 16'h90b6, 16'h90b7 	:	val_out <= 16'h4d07;
         16'h90b8, 16'h90b9, 16'h90ba, 16'h90bb, 16'h90bc, 16'h90bd, 16'h90be, 16'h90bf 	:	val_out <= 16'h4cf0;
         16'h90c0, 16'h90c1, 16'h90c2, 16'h90c3, 16'h90c4, 16'h90c5, 16'h90c6, 16'h90c7 	:	val_out <= 16'h4cd9;
         16'h90c8, 16'h90c9, 16'h90ca, 16'h90cb, 16'h90cc, 16'h90cd, 16'h90ce, 16'h90cf 	:	val_out <= 16'h4cc2;
         16'h90d0, 16'h90d1, 16'h90d2, 16'h90d3, 16'h90d4, 16'h90d5, 16'h90d6, 16'h90d7 	:	val_out <= 16'h4cab;
         16'h90d8, 16'h90d9, 16'h90da, 16'h90db, 16'h90dc, 16'h90dd, 16'h90de, 16'h90df 	:	val_out <= 16'h4c94;
         16'h90e0, 16'h90e1, 16'h90e2, 16'h90e3, 16'h90e4, 16'h90e5, 16'h90e6, 16'h90e7 	:	val_out <= 16'h4c7d;
         16'h90e8, 16'h90e9, 16'h90ea, 16'h90eb, 16'h90ec, 16'h90ed, 16'h90ee, 16'h90ef 	:	val_out <= 16'h4c66;
         16'h90f0, 16'h90f1, 16'h90f2, 16'h90f3, 16'h90f4, 16'h90f5, 16'h90f6, 16'h90f7 	:	val_out <= 16'h4c4f;
         16'h90f8, 16'h90f9, 16'h90fa, 16'h90fb, 16'h90fc, 16'h90fd, 16'h90fe, 16'h90ff 	:	val_out <= 16'h4c38;
         16'h9100, 16'h9101, 16'h9102, 16'h9103, 16'h9104, 16'h9105, 16'h9106, 16'h9107 	:	val_out <= 16'h4c21;
         16'h9108, 16'h9109, 16'h910a, 16'h910b, 16'h910c, 16'h910d, 16'h910e, 16'h910f 	:	val_out <= 16'h4c0a;
         16'h9110, 16'h9111, 16'h9112, 16'h9113, 16'h9114, 16'h9115, 16'h9116, 16'h9117 	:	val_out <= 16'h4bf3;
         16'h9118, 16'h9119, 16'h911a, 16'h911b, 16'h911c, 16'h911d, 16'h911e, 16'h911f 	:	val_out <= 16'h4bdc;
         16'h9120, 16'h9121, 16'h9122, 16'h9123, 16'h9124, 16'h9125, 16'h9126, 16'h9127 	:	val_out <= 16'h4bc5;
         16'h9128, 16'h9129, 16'h912a, 16'h912b, 16'h912c, 16'h912d, 16'h912e, 16'h912f 	:	val_out <= 16'h4bae;
         16'h9130, 16'h9131, 16'h9132, 16'h9133, 16'h9134, 16'h9135, 16'h9136, 16'h9137 	:	val_out <= 16'h4b97;
         16'h9138, 16'h9139, 16'h913a, 16'h913b, 16'h913c, 16'h913d, 16'h913e, 16'h913f 	:	val_out <= 16'h4b80;
         16'h9140, 16'h9141, 16'h9142, 16'h9143, 16'h9144, 16'h9145, 16'h9146, 16'h9147 	:	val_out <= 16'h4b69;
         16'h9148, 16'h9149, 16'h914a, 16'h914b, 16'h914c, 16'h914d, 16'h914e, 16'h914f 	:	val_out <= 16'h4b52;
         16'h9150, 16'h9151, 16'h9152, 16'h9153, 16'h9154, 16'h9155, 16'h9156, 16'h9157 	:	val_out <= 16'h4b3b;
         16'h9158, 16'h9159, 16'h915a, 16'h915b, 16'h915c, 16'h915d, 16'h915e, 16'h915f 	:	val_out <= 16'h4b24;
         16'h9160, 16'h9161, 16'h9162, 16'h9163, 16'h9164, 16'h9165, 16'h9166, 16'h9167 	:	val_out <= 16'h4b0d;
         16'h9168, 16'h9169, 16'h916a, 16'h916b, 16'h916c, 16'h916d, 16'h916e, 16'h916f 	:	val_out <= 16'h4af7;
         16'h9170, 16'h9171, 16'h9172, 16'h9173, 16'h9174, 16'h9175, 16'h9176, 16'h9177 	:	val_out <= 16'h4ae0;
         16'h9178, 16'h9179, 16'h917a, 16'h917b, 16'h917c, 16'h917d, 16'h917e, 16'h917f 	:	val_out <= 16'h4ac9;
         16'h9180, 16'h9181, 16'h9182, 16'h9183, 16'h9184, 16'h9185, 16'h9186, 16'h9187 	:	val_out <= 16'h4ab2;
         16'h9188, 16'h9189, 16'h918a, 16'h918b, 16'h918c, 16'h918d, 16'h918e, 16'h918f 	:	val_out <= 16'h4a9b;
         16'h9190, 16'h9191, 16'h9192, 16'h9193, 16'h9194, 16'h9195, 16'h9196, 16'h9197 	:	val_out <= 16'h4a84;
         16'h9198, 16'h9199, 16'h919a, 16'h919b, 16'h919c, 16'h919d, 16'h919e, 16'h919f 	:	val_out <= 16'h4a6d;
         16'h91a0, 16'h91a1, 16'h91a2, 16'h91a3, 16'h91a4, 16'h91a5, 16'h91a6, 16'h91a7 	:	val_out <= 16'h4a57;
         16'h91a8, 16'h91a9, 16'h91aa, 16'h91ab, 16'h91ac, 16'h91ad, 16'h91ae, 16'h91af 	:	val_out <= 16'h4a40;
         16'h91b0, 16'h91b1, 16'h91b2, 16'h91b3, 16'h91b4, 16'h91b5, 16'h91b6, 16'h91b7 	:	val_out <= 16'h4a29;
         16'h91b8, 16'h91b9, 16'h91ba, 16'h91bb, 16'h91bc, 16'h91bd, 16'h91be, 16'h91bf 	:	val_out <= 16'h4a12;
         16'h91c0, 16'h91c1, 16'h91c2, 16'h91c3, 16'h91c4, 16'h91c5, 16'h91c6, 16'h91c7 	:	val_out <= 16'h49fb;
         16'h91c8, 16'h91c9, 16'h91ca, 16'h91cb, 16'h91cc, 16'h91cd, 16'h91ce, 16'h91cf 	:	val_out <= 16'h49e5;
         16'h91d0, 16'h91d1, 16'h91d2, 16'h91d3, 16'h91d4, 16'h91d5, 16'h91d6, 16'h91d7 	:	val_out <= 16'h49ce;
         16'h91d8, 16'h91d9, 16'h91da, 16'h91db, 16'h91dc, 16'h91dd, 16'h91de, 16'h91df 	:	val_out <= 16'h49b7;
         16'h91e0, 16'h91e1, 16'h91e2, 16'h91e3, 16'h91e4, 16'h91e5, 16'h91e6, 16'h91e7 	:	val_out <= 16'h49a0;
         16'h91e8, 16'h91e9, 16'h91ea, 16'h91eb, 16'h91ec, 16'h91ed, 16'h91ee, 16'h91ef 	:	val_out <= 16'h498a;
         16'h91f0, 16'h91f1, 16'h91f2, 16'h91f3, 16'h91f4, 16'h91f5, 16'h91f6, 16'h91f7 	:	val_out <= 16'h4973;
         16'h91f8, 16'h91f9, 16'h91fa, 16'h91fb, 16'h91fc, 16'h91fd, 16'h91fe, 16'h91ff 	:	val_out <= 16'h495c;
         16'h9200, 16'h9201, 16'h9202, 16'h9203, 16'h9204, 16'h9205, 16'h9206, 16'h9207 	:	val_out <= 16'h4945;
         16'h9208, 16'h9209, 16'h920a, 16'h920b, 16'h920c, 16'h920d, 16'h920e, 16'h920f 	:	val_out <= 16'h492f;
         16'h9210, 16'h9211, 16'h9212, 16'h9213, 16'h9214, 16'h9215, 16'h9216, 16'h9217 	:	val_out <= 16'h4918;
         16'h9218, 16'h9219, 16'h921a, 16'h921b, 16'h921c, 16'h921d, 16'h921e, 16'h921f 	:	val_out <= 16'h4901;
         16'h9220, 16'h9221, 16'h9222, 16'h9223, 16'h9224, 16'h9225, 16'h9226, 16'h9227 	:	val_out <= 16'h48eb;
         16'h9228, 16'h9229, 16'h922a, 16'h922b, 16'h922c, 16'h922d, 16'h922e, 16'h922f 	:	val_out <= 16'h48d4;
         16'h9230, 16'h9231, 16'h9232, 16'h9233, 16'h9234, 16'h9235, 16'h9236, 16'h9237 	:	val_out <= 16'h48bd;
         16'h9238, 16'h9239, 16'h923a, 16'h923b, 16'h923c, 16'h923d, 16'h923e, 16'h923f 	:	val_out <= 16'h48a7;
         16'h9240, 16'h9241, 16'h9242, 16'h9243, 16'h9244, 16'h9245, 16'h9246, 16'h9247 	:	val_out <= 16'h4890;
         16'h9248, 16'h9249, 16'h924a, 16'h924b, 16'h924c, 16'h924d, 16'h924e, 16'h924f 	:	val_out <= 16'h4879;
         16'h9250, 16'h9251, 16'h9252, 16'h9253, 16'h9254, 16'h9255, 16'h9256, 16'h9257 	:	val_out <= 16'h4863;
         16'h9258, 16'h9259, 16'h925a, 16'h925b, 16'h925c, 16'h925d, 16'h925e, 16'h925f 	:	val_out <= 16'h484c;
         16'h9260, 16'h9261, 16'h9262, 16'h9263, 16'h9264, 16'h9265, 16'h9266, 16'h9267 	:	val_out <= 16'h4835;
         16'h9268, 16'h9269, 16'h926a, 16'h926b, 16'h926c, 16'h926d, 16'h926e, 16'h926f 	:	val_out <= 16'h481f;
         16'h9270, 16'h9271, 16'h9272, 16'h9273, 16'h9274, 16'h9275, 16'h9276, 16'h9277 	:	val_out <= 16'h4808;
         16'h9278, 16'h9279, 16'h927a, 16'h927b, 16'h927c, 16'h927d, 16'h927e, 16'h927f 	:	val_out <= 16'h47f2;
         16'h9280, 16'h9281, 16'h9282, 16'h9283, 16'h9284, 16'h9285, 16'h9286, 16'h9287 	:	val_out <= 16'h47db;
         16'h9288, 16'h9289, 16'h928a, 16'h928b, 16'h928c, 16'h928d, 16'h928e, 16'h928f 	:	val_out <= 16'h47c4;
         16'h9290, 16'h9291, 16'h9292, 16'h9293, 16'h9294, 16'h9295, 16'h9296, 16'h9297 	:	val_out <= 16'h47ae;
         16'h9298, 16'h9299, 16'h929a, 16'h929b, 16'h929c, 16'h929d, 16'h929e, 16'h929f 	:	val_out <= 16'h4797;
         16'h92a0, 16'h92a1, 16'h92a2, 16'h92a3, 16'h92a4, 16'h92a5, 16'h92a6, 16'h92a7 	:	val_out <= 16'h4781;
         16'h92a8, 16'h92a9, 16'h92aa, 16'h92ab, 16'h92ac, 16'h92ad, 16'h92ae, 16'h92af 	:	val_out <= 16'h476a;
         16'h92b0, 16'h92b1, 16'h92b2, 16'h92b3, 16'h92b4, 16'h92b5, 16'h92b6, 16'h92b7 	:	val_out <= 16'h4754;
         16'h92b8, 16'h92b9, 16'h92ba, 16'h92bb, 16'h92bc, 16'h92bd, 16'h92be, 16'h92bf 	:	val_out <= 16'h473d;
         16'h92c0, 16'h92c1, 16'h92c2, 16'h92c3, 16'h92c4, 16'h92c5, 16'h92c6, 16'h92c7 	:	val_out <= 16'h4727;
         16'h92c8, 16'h92c9, 16'h92ca, 16'h92cb, 16'h92cc, 16'h92cd, 16'h92ce, 16'h92cf 	:	val_out <= 16'h4710;
         16'h92d0, 16'h92d1, 16'h92d2, 16'h92d3, 16'h92d4, 16'h92d5, 16'h92d6, 16'h92d7 	:	val_out <= 16'h46f9;
         16'h92d8, 16'h92d9, 16'h92da, 16'h92db, 16'h92dc, 16'h92dd, 16'h92de, 16'h92df 	:	val_out <= 16'h46e3;
         16'h92e0, 16'h92e1, 16'h92e2, 16'h92e3, 16'h92e4, 16'h92e5, 16'h92e6, 16'h92e7 	:	val_out <= 16'h46cd;
         16'h92e8, 16'h92e9, 16'h92ea, 16'h92eb, 16'h92ec, 16'h92ed, 16'h92ee, 16'h92ef 	:	val_out <= 16'h46b6;
         16'h92f0, 16'h92f1, 16'h92f2, 16'h92f3, 16'h92f4, 16'h92f5, 16'h92f6, 16'h92f7 	:	val_out <= 16'h46a0;
         16'h92f8, 16'h92f9, 16'h92fa, 16'h92fb, 16'h92fc, 16'h92fd, 16'h92fe, 16'h92ff 	:	val_out <= 16'h4689;
         16'h9300, 16'h9301, 16'h9302, 16'h9303, 16'h9304, 16'h9305, 16'h9306, 16'h9307 	:	val_out <= 16'h4673;
         16'h9308, 16'h9309, 16'h930a, 16'h930b, 16'h930c, 16'h930d, 16'h930e, 16'h930f 	:	val_out <= 16'h465c;
         16'h9310, 16'h9311, 16'h9312, 16'h9313, 16'h9314, 16'h9315, 16'h9316, 16'h9317 	:	val_out <= 16'h4646;
         16'h9318, 16'h9319, 16'h931a, 16'h931b, 16'h931c, 16'h931d, 16'h931e, 16'h931f 	:	val_out <= 16'h462f;
         16'h9320, 16'h9321, 16'h9322, 16'h9323, 16'h9324, 16'h9325, 16'h9326, 16'h9327 	:	val_out <= 16'h4619;
         16'h9328, 16'h9329, 16'h932a, 16'h932b, 16'h932c, 16'h932d, 16'h932e, 16'h932f 	:	val_out <= 16'h4602;
         16'h9330, 16'h9331, 16'h9332, 16'h9333, 16'h9334, 16'h9335, 16'h9336, 16'h9337 	:	val_out <= 16'h45ec;
         16'h9338, 16'h9339, 16'h933a, 16'h933b, 16'h933c, 16'h933d, 16'h933e, 16'h933f 	:	val_out <= 16'h45d6;
         16'h9340, 16'h9341, 16'h9342, 16'h9343, 16'h9344, 16'h9345, 16'h9346, 16'h9347 	:	val_out <= 16'h45bf;
         16'h9348, 16'h9349, 16'h934a, 16'h934b, 16'h934c, 16'h934d, 16'h934e, 16'h934f 	:	val_out <= 16'h45a9;
         16'h9350, 16'h9351, 16'h9352, 16'h9353, 16'h9354, 16'h9355, 16'h9356, 16'h9357 	:	val_out <= 16'h4593;
         16'h9358, 16'h9359, 16'h935a, 16'h935b, 16'h935c, 16'h935d, 16'h935e, 16'h935f 	:	val_out <= 16'h457c;
         16'h9360, 16'h9361, 16'h9362, 16'h9363, 16'h9364, 16'h9365, 16'h9366, 16'h9367 	:	val_out <= 16'h4566;
         16'h9368, 16'h9369, 16'h936a, 16'h936b, 16'h936c, 16'h936d, 16'h936e, 16'h936f 	:	val_out <= 16'h4550;
         16'h9370, 16'h9371, 16'h9372, 16'h9373, 16'h9374, 16'h9375, 16'h9376, 16'h9377 	:	val_out <= 16'h4539;
         16'h9378, 16'h9379, 16'h937a, 16'h937b, 16'h937c, 16'h937d, 16'h937e, 16'h937f 	:	val_out <= 16'h4523;
         16'h9380, 16'h9381, 16'h9382, 16'h9383, 16'h9384, 16'h9385, 16'h9386, 16'h9387 	:	val_out <= 16'h450d;
         16'h9388, 16'h9389, 16'h938a, 16'h938b, 16'h938c, 16'h938d, 16'h938e, 16'h938f 	:	val_out <= 16'h44f6;
         16'h9390, 16'h9391, 16'h9392, 16'h9393, 16'h9394, 16'h9395, 16'h9396, 16'h9397 	:	val_out <= 16'h44e0;
         16'h9398, 16'h9399, 16'h939a, 16'h939b, 16'h939c, 16'h939d, 16'h939e, 16'h939f 	:	val_out <= 16'h44ca;
         16'h93a0, 16'h93a1, 16'h93a2, 16'h93a3, 16'h93a4, 16'h93a5, 16'h93a6, 16'h93a7 	:	val_out <= 16'h44b3;
         16'h93a8, 16'h93a9, 16'h93aa, 16'h93ab, 16'h93ac, 16'h93ad, 16'h93ae, 16'h93af 	:	val_out <= 16'h449d;
         16'h93b0, 16'h93b1, 16'h93b2, 16'h93b3, 16'h93b4, 16'h93b5, 16'h93b6, 16'h93b7 	:	val_out <= 16'h4487;
         16'h93b8, 16'h93b9, 16'h93ba, 16'h93bb, 16'h93bc, 16'h93bd, 16'h93be, 16'h93bf 	:	val_out <= 16'h4471;
         16'h93c0, 16'h93c1, 16'h93c2, 16'h93c3, 16'h93c4, 16'h93c5, 16'h93c6, 16'h93c7 	:	val_out <= 16'h445a;
         16'h93c8, 16'h93c9, 16'h93ca, 16'h93cb, 16'h93cc, 16'h93cd, 16'h93ce, 16'h93cf 	:	val_out <= 16'h4444;
         16'h93d0, 16'h93d1, 16'h93d2, 16'h93d3, 16'h93d4, 16'h93d5, 16'h93d6, 16'h93d7 	:	val_out <= 16'h442e;
         16'h93d8, 16'h93d9, 16'h93da, 16'h93db, 16'h93dc, 16'h93dd, 16'h93de, 16'h93df 	:	val_out <= 16'h4418;
         16'h93e0, 16'h93e1, 16'h93e2, 16'h93e3, 16'h93e4, 16'h93e5, 16'h93e6, 16'h93e7 	:	val_out <= 16'h4402;
         16'h93e8, 16'h93e9, 16'h93ea, 16'h93eb, 16'h93ec, 16'h93ed, 16'h93ee, 16'h93ef 	:	val_out <= 16'h43eb;
         16'h93f0, 16'h93f1, 16'h93f2, 16'h93f3, 16'h93f4, 16'h93f5, 16'h93f6, 16'h93f7 	:	val_out <= 16'h43d5;
         16'h93f8, 16'h93f9, 16'h93fa, 16'h93fb, 16'h93fc, 16'h93fd, 16'h93fe, 16'h93ff 	:	val_out <= 16'h43bf;
         16'h9400, 16'h9401, 16'h9402, 16'h9403, 16'h9404, 16'h9405, 16'h9406, 16'h9407 	:	val_out <= 16'h43a9;
         16'h9408, 16'h9409, 16'h940a, 16'h940b, 16'h940c, 16'h940d, 16'h940e, 16'h940f 	:	val_out <= 16'h4393;
         16'h9410, 16'h9411, 16'h9412, 16'h9413, 16'h9414, 16'h9415, 16'h9416, 16'h9417 	:	val_out <= 16'h437c;
         16'h9418, 16'h9419, 16'h941a, 16'h941b, 16'h941c, 16'h941d, 16'h941e, 16'h941f 	:	val_out <= 16'h4366;
         16'h9420, 16'h9421, 16'h9422, 16'h9423, 16'h9424, 16'h9425, 16'h9426, 16'h9427 	:	val_out <= 16'h4350;
         16'h9428, 16'h9429, 16'h942a, 16'h942b, 16'h942c, 16'h942d, 16'h942e, 16'h942f 	:	val_out <= 16'h433a;
         16'h9430, 16'h9431, 16'h9432, 16'h9433, 16'h9434, 16'h9435, 16'h9436, 16'h9437 	:	val_out <= 16'h4324;
         16'h9438, 16'h9439, 16'h943a, 16'h943b, 16'h943c, 16'h943d, 16'h943e, 16'h943f 	:	val_out <= 16'h430e;
         16'h9440, 16'h9441, 16'h9442, 16'h9443, 16'h9444, 16'h9445, 16'h9446, 16'h9447 	:	val_out <= 16'h42f8;
         16'h9448, 16'h9449, 16'h944a, 16'h944b, 16'h944c, 16'h944d, 16'h944e, 16'h944f 	:	val_out <= 16'h42e2;
         16'h9450, 16'h9451, 16'h9452, 16'h9453, 16'h9454, 16'h9455, 16'h9456, 16'h9457 	:	val_out <= 16'h42cc;
         16'h9458, 16'h9459, 16'h945a, 16'h945b, 16'h945c, 16'h945d, 16'h945e, 16'h945f 	:	val_out <= 16'h42b6;
         16'h9460, 16'h9461, 16'h9462, 16'h9463, 16'h9464, 16'h9465, 16'h9466, 16'h9467 	:	val_out <= 16'h429f;
         16'h9468, 16'h9469, 16'h946a, 16'h946b, 16'h946c, 16'h946d, 16'h946e, 16'h946f 	:	val_out <= 16'h4289;
         16'h9470, 16'h9471, 16'h9472, 16'h9473, 16'h9474, 16'h9475, 16'h9476, 16'h9477 	:	val_out <= 16'h4273;
         16'h9478, 16'h9479, 16'h947a, 16'h947b, 16'h947c, 16'h947d, 16'h947e, 16'h947f 	:	val_out <= 16'h425d;
         16'h9480, 16'h9481, 16'h9482, 16'h9483, 16'h9484, 16'h9485, 16'h9486, 16'h9487 	:	val_out <= 16'h4247;
         16'h9488, 16'h9489, 16'h948a, 16'h948b, 16'h948c, 16'h948d, 16'h948e, 16'h948f 	:	val_out <= 16'h4231;
         16'h9490, 16'h9491, 16'h9492, 16'h9493, 16'h9494, 16'h9495, 16'h9496, 16'h9497 	:	val_out <= 16'h421b;
         16'h9498, 16'h9499, 16'h949a, 16'h949b, 16'h949c, 16'h949d, 16'h949e, 16'h949f 	:	val_out <= 16'h4205;
         16'h94a0, 16'h94a1, 16'h94a2, 16'h94a3, 16'h94a4, 16'h94a5, 16'h94a6, 16'h94a7 	:	val_out <= 16'h41ef;
         16'h94a8, 16'h94a9, 16'h94aa, 16'h94ab, 16'h94ac, 16'h94ad, 16'h94ae, 16'h94af 	:	val_out <= 16'h41d9;
         16'h94b0, 16'h94b1, 16'h94b2, 16'h94b3, 16'h94b4, 16'h94b5, 16'h94b6, 16'h94b7 	:	val_out <= 16'h41c3;
         16'h94b8, 16'h94b9, 16'h94ba, 16'h94bb, 16'h94bc, 16'h94bd, 16'h94be, 16'h94bf 	:	val_out <= 16'h41ad;
         16'h94c0, 16'h94c1, 16'h94c2, 16'h94c3, 16'h94c4, 16'h94c5, 16'h94c6, 16'h94c7 	:	val_out <= 16'h4197;
         16'h94c8, 16'h94c9, 16'h94ca, 16'h94cb, 16'h94cc, 16'h94cd, 16'h94ce, 16'h94cf 	:	val_out <= 16'h4182;
         16'h94d0, 16'h94d1, 16'h94d2, 16'h94d3, 16'h94d4, 16'h94d5, 16'h94d6, 16'h94d7 	:	val_out <= 16'h416c;
         16'h94d8, 16'h94d9, 16'h94da, 16'h94db, 16'h94dc, 16'h94dd, 16'h94de, 16'h94df 	:	val_out <= 16'h4156;
         16'h94e0, 16'h94e1, 16'h94e2, 16'h94e3, 16'h94e4, 16'h94e5, 16'h94e6, 16'h94e7 	:	val_out <= 16'h4140;
         16'h94e8, 16'h94e9, 16'h94ea, 16'h94eb, 16'h94ec, 16'h94ed, 16'h94ee, 16'h94ef 	:	val_out <= 16'h412a;
         16'h94f0, 16'h94f1, 16'h94f2, 16'h94f3, 16'h94f4, 16'h94f5, 16'h94f6, 16'h94f7 	:	val_out <= 16'h4114;
         16'h94f8, 16'h94f9, 16'h94fa, 16'h94fb, 16'h94fc, 16'h94fd, 16'h94fe, 16'h94ff 	:	val_out <= 16'h40fe;
         16'h9500, 16'h9501, 16'h9502, 16'h9503, 16'h9504, 16'h9505, 16'h9506, 16'h9507 	:	val_out <= 16'h40e8;
         16'h9508, 16'h9509, 16'h950a, 16'h950b, 16'h950c, 16'h950d, 16'h950e, 16'h950f 	:	val_out <= 16'h40d2;
         16'h9510, 16'h9511, 16'h9512, 16'h9513, 16'h9514, 16'h9515, 16'h9516, 16'h9517 	:	val_out <= 16'h40bc;
         16'h9518, 16'h9519, 16'h951a, 16'h951b, 16'h951c, 16'h951d, 16'h951e, 16'h951f 	:	val_out <= 16'h40a7;
         16'h9520, 16'h9521, 16'h9522, 16'h9523, 16'h9524, 16'h9525, 16'h9526, 16'h9527 	:	val_out <= 16'h4091;
         16'h9528, 16'h9529, 16'h952a, 16'h952b, 16'h952c, 16'h952d, 16'h952e, 16'h952f 	:	val_out <= 16'h407b;
         16'h9530, 16'h9531, 16'h9532, 16'h9533, 16'h9534, 16'h9535, 16'h9536, 16'h9537 	:	val_out <= 16'h4065;
         16'h9538, 16'h9539, 16'h953a, 16'h953b, 16'h953c, 16'h953d, 16'h953e, 16'h953f 	:	val_out <= 16'h404f;
         16'h9540, 16'h9541, 16'h9542, 16'h9543, 16'h9544, 16'h9545, 16'h9546, 16'h9547 	:	val_out <= 16'h403a;
         16'h9548, 16'h9549, 16'h954a, 16'h954b, 16'h954c, 16'h954d, 16'h954e, 16'h954f 	:	val_out <= 16'h4024;
         16'h9550, 16'h9551, 16'h9552, 16'h9553, 16'h9554, 16'h9555, 16'h9556, 16'h9557 	:	val_out <= 16'h400e;
         16'h9558, 16'h9559, 16'h955a, 16'h955b, 16'h955c, 16'h955d, 16'h955e, 16'h955f 	:	val_out <= 16'h3ff8;
         16'h9560, 16'h9561, 16'h9562, 16'h9563, 16'h9564, 16'h9565, 16'h9566, 16'h9567 	:	val_out <= 16'h3fe2;
         16'h9568, 16'h9569, 16'h956a, 16'h956b, 16'h956c, 16'h956d, 16'h956e, 16'h956f 	:	val_out <= 16'h3fcd;
         16'h9570, 16'h9571, 16'h9572, 16'h9573, 16'h9574, 16'h9575, 16'h9576, 16'h9577 	:	val_out <= 16'h3fb7;
         16'h9578, 16'h9579, 16'h957a, 16'h957b, 16'h957c, 16'h957d, 16'h957e, 16'h957f 	:	val_out <= 16'h3fa1;
         16'h9580, 16'h9581, 16'h9582, 16'h9583, 16'h9584, 16'h9585, 16'h9586, 16'h9587 	:	val_out <= 16'h3f8c;
         16'h9588, 16'h9589, 16'h958a, 16'h958b, 16'h958c, 16'h958d, 16'h958e, 16'h958f 	:	val_out <= 16'h3f76;
         16'h9590, 16'h9591, 16'h9592, 16'h9593, 16'h9594, 16'h9595, 16'h9596, 16'h9597 	:	val_out <= 16'h3f60;
         16'h9598, 16'h9599, 16'h959a, 16'h959b, 16'h959c, 16'h959d, 16'h959e, 16'h959f 	:	val_out <= 16'h3f4a;
         16'h95a0, 16'h95a1, 16'h95a2, 16'h95a3, 16'h95a4, 16'h95a5, 16'h95a6, 16'h95a7 	:	val_out <= 16'h3f35;
         16'h95a8, 16'h95a9, 16'h95aa, 16'h95ab, 16'h95ac, 16'h95ad, 16'h95ae, 16'h95af 	:	val_out <= 16'h3f1f;
         16'h95b0, 16'h95b1, 16'h95b2, 16'h95b3, 16'h95b4, 16'h95b5, 16'h95b6, 16'h95b7 	:	val_out <= 16'h3f09;
         16'h95b8, 16'h95b9, 16'h95ba, 16'h95bb, 16'h95bc, 16'h95bd, 16'h95be, 16'h95bf 	:	val_out <= 16'h3ef4;
         16'h95c0, 16'h95c1, 16'h95c2, 16'h95c3, 16'h95c4, 16'h95c5, 16'h95c6, 16'h95c7 	:	val_out <= 16'h3ede;
         16'h95c8, 16'h95c9, 16'h95ca, 16'h95cb, 16'h95cc, 16'h95cd, 16'h95ce, 16'h95cf 	:	val_out <= 16'h3ec9;
         16'h95d0, 16'h95d1, 16'h95d2, 16'h95d3, 16'h95d4, 16'h95d5, 16'h95d6, 16'h95d7 	:	val_out <= 16'h3eb3;
         16'h95d8, 16'h95d9, 16'h95da, 16'h95db, 16'h95dc, 16'h95dd, 16'h95de, 16'h95df 	:	val_out <= 16'h3e9d;
         16'h95e0, 16'h95e1, 16'h95e2, 16'h95e3, 16'h95e4, 16'h95e5, 16'h95e6, 16'h95e7 	:	val_out <= 16'h3e88;
         16'h95e8, 16'h95e9, 16'h95ea, 16'h95eb, 16'h95ec, 16'h95ed, 16'h95ee, 16'h95ef 	:	val_out <= 16'h3e72;
         16'h95f0, 16'h95f1, 16'h95f2, 16'h95f3, 16'h95f4, 16'h95f5, 16'h95f6, 16'h95f7 	:	val_out <= 16'h3e5d;
         16'h95f8, 16'h95f9, 16'h95fa, 16'h95fb, 16'h95fc, 16'h95fd, 16'h95fe, 16'h95ff 	:	val_out <= 16'h3e47;
         16'h9600, 16'h9601, 16'h9602, 16'h9603, 16'h9604, 16'h9605, 16'h9606, 16'h9607 	:	val_out <= 16'h3e31;
         16'h9608, 16'h9609, 16'h960a, 16'h960b, 16'h960c, 16'h960d, 16'h960e, 16'h960f 	:	val_out <= 16'h3e1c;
         16'h9610, 16'h9611, 16'h9612, 16'h9613, 16'h9614, 16'h9615, 16'h9616, 16'h9617 	:	val_out <= 16'h3e06;
         16'h9618, 16'h9619, 16'h961a, 16'h961b, 16'h961c, 16'h961d, 16'h961e, 16'h961f 	:	val_out <= 16'h3df1;
         16'h9620, 16'h9621, 16'h9622, 16'h9623, 16'h9624, 16'h9625, 16'h9626, 16'h9627 	:	val_out <= 16'h3ddb;
         16'h9628, 16'h9629, 16'h962a, 16'h962b, 16'h962c, 16'h962d, 16'h962e, 16'h962f 	:	val_out <= 16'h3dc6;
         16'h9630, 16'h9631, 16'h9632, 16'h9633, 16'h9634, 16'h9635, 16'h9636, 16'h9637 	:	val_out <= 16'h3db0;
         16'h9638, 16'h9639, 16'h963a, 16'h963b, 16'h963c, 16'h963d, 16'h963e, 16'h963f 	:	val_out <= 16'h3d9b;
         16'h9640, 16'h9641, 16'h9642, 16'h9643, 16'h9644, 16'h9645, 16'h9646, 16'h9647 	:	val_out <= 16'h3d85;
         16'h9648, 16'h9649, 16'h964a, 16'h964b, 16'h964c, 16'h964d, 16'h964e, 16'h964f 	:	val_out <= 16'h3d70;
         16'h9650, 16'h9651, 16'h9652, 16'h9653, 16'h9654, 16'h9655, 16'h9656, 16'h9657 	:	val_out <= 16'h3d5a;
         16'h9658, 16'h9659, 16'h965a, 16'h965b, 16'h965c, 16'h965d, 16'h965e, 16'h965f 	:	val_out <= 16'h3d45;
         16'h9660, 16'h9661, 16'h9662, 16'h9663, 16'h9664, 16'h9665, 16'h9666, 16'h9667 	:	val_out <= 16'h3d2f;
         16'h9668, 16'h9669, 16'h966a, 16'h966b, 16'h966c, 16'h966d, 16'h966e, 16'h966f 	:	val_out <= 16'h3d1a;
         16'h9670, 16'h9671, 16'h9672, 16'h9673, 16'h9674, 16'h9675, 16'h9676, 16'h9677 	:	val_out <= 16'h3d05;
         16'h9678, 16'h9679, 16'h967a, 16'h967b, 16'h967c, 16'h967d, 16'h967e, 16'h967f 	:	val_out <= 16'h3cef;
         16'h9680, 16'h9681, 16'h9682, 16'h9683, 16'h9684, 16'h9685, 16'h9686, 16'h9687 	:	val_out <= 16'h3cda;
         16'h9688, 16'h9689, 16'h968a, 16'h968b, 16'h968c, 16'h968d, 16'h968e, 16'h968f 	:	val_out <= 16'h3cc4;
         16'h9690, 16'h9691, 16'h9692, 16'h9693, 16'h9694, 16'h9695, 16'h9696, 16'h9697 	:	val_out <= 16'h3caf;
         16'h9698, 16'h9699, 16'h969a, 16'h969b, 16'h969c, 16'h969d, 16'h969e, 16'h969f 	:	val_out <= 16'h3c9a;
         16'h96a0, 16'h96a1, 16'h96a2, 16'h96a3, 16'h96a4, 16'h96a5, 16'h96a6, 16'h96a7 	:	val_out <= 16'h3c84;
         16'h96a8, 16'h96a9, 16'h96aa, 16'h96ab, 16'h96ac, 16'h96ad, 16'h96ae, 16'h96af 	:	val_out <= 16'h3c6f;
         16'h96b0, 16'h96b1, 16'h96b2, 16'h96b3, 16'h96b4, 16'h96b5, 16'h96b6, 16'h96b7 	:	val_out <= 16'h3c5a;
         16'h96b8, 16'h96b9, 16'h96ba, 16'h96bb, 16'h96bc, 16'h96bd, 16'h96be, 16'h96bf 	:	val_out <= 16'h3c44;
         16'h96c0, 16'h96c1, 16'h96c2, 16'h96c3, 16'h96c4, 16'h96c5, 16'h96c6, 16'h96c7 	:	val_out <= 16'h3c2f;
         16'h96c8, 16'h96c9, 16'h96ca, 16'h96cb, 16'h96cc, 16'h96cd, 16'h96ce, 16'h96cf 	:	val_out <= 16'h3c1a;
         16'h96d0, 16'h96d1, 16'h96d2, 16'h96d3, 16'h96d4, 16'h96d5, 16'h96d6, 16'h96d7 	:	val_out <= 16'h3c04;
         16'h96d8, 16'h96d9, 16'h96da, 16'h96db, 16'h96dc, 16'h96dd, 16'h96de, 16'h96df 	:	val_out <= 16'h3bef;
         16'h96e0, 16'h96e1, 16'h96e2, 16'h96e3, 16'h96e4, 16'h96e5, 16'h96e6, 16'h96e7 	:	val_out <= 16'h3bda;
         16'h96e8, 16'h96e9, 16'h96ea, 16'h96eb, 16'h96ec, 16'h96ed, 16'h96ee, 16'h96ef 	:	val_out <= 16'h3bc4;
         16'h96f0, 16'h96f1, 16'h96f2, 16'h96f3, 16'h96f4, 16'h96f5, 16'h96f6, 16'h96f7 	:	val_out <= 16'h3baf;
         16'h96f8, 16'h96f9, 16'h96fa, 16'h96fb, 16'h96fc, 16'h96fd, 16'h96fe, 16'h96ff 	:	val_out <= 16'h3b9a;
         16'h9700, 16'h9701, 16'h9702, 16'h9703, 16'h9704, 16'h9705, 16'h9706, 16'h9707 	:	val_out <= 16'h3b85;
         16'h9708, 16'h9709, 16'h970a, 16'h970b, 16'h970c, 16'h970d, 16'h970e, 16'h970f 	:	val_out <= 16'h3b6f;
         16'h9710, 16'h9711, 16'h9712, 16'h9713, 16'h9714, 16'h9715, 16'h9716, 16'h9717 	:	val_out <= 16'h3b5a;
         16'h9718, 16'h9719, 16'h971a, 16'h971b, 16'h971c, 16'h971d, 16'h971e, 16'h971f 	:	val_out <= 16'h3b45;
         16'h9720, 16'h9721, 16'h9722, 16'h9723, 16'h9724, 16'h9725, 16'h9726, 16'h9727 	:	val_out <= 16'h3b30;
         16'h9728, 16'h9729, 16'h972a, 16'h972b, 16'h972c, 16'h972d, 16'h972e, 16'h972f 	:	val_out <= 16'h3b1b;
         16'h9730, 16'h9731, 16'h9732, 16'h9733, 16'h9734, 16'h9735, 16'h9736, 16'h9737 	:	val_out <= 16'h3b05;
         16'h9738, 16'h9739, 16'h973a, 16'h973b, 16'h973c, 16'h973d, 16'h973e, 16'h973f 	:	val_out <= 16'h3af0;
         16'h9740, 16'h9741, 16'h9742, 16'h9743, 16'h9744, 16'h9745, 16'h9746, 16'h9747 	:	val_out <= 16'h3adb;
         16'h9748, 16'h9749, 16'h974a, 16'h974b, 16'h974c, 16'h974d, 16'h974e, 16'h974f 	:	val_out <= 16'h3ac6;
         16'h9750, 16'h9751, 16'h9752, 16'h9753, 16'h9754, 16'h9755, 16'h9756, 16'h9757 	:	val_out <= 16'h3ab1;
         16'h9758, 16'h9759, 16'h975a, 16'h975b, 16'h975c, 16'h975d, 16'h975e, 16'h975f 	:	val_out <= 16'h3a9c;
         16'h9760, 16'h9761, 16'h9762, 16'h9763, 16'h9764, 16'h9765, 16'h9766, 16'h9767 	:	val_out <= 16'h3a87;
         16'h9768, 16'h9769, 16'h976a, 16'h976b, 16'h976c, 16'h976d, 16'h976e, 16'h976f 	:	val_out <= 16'h3a72;
         16'h9770, 16'h9771, 16'h9772, 16'h9773, 16'h9774, 16'h9775, 16'h9776, 16'h9777 	:	val_out <= 16'h3a5c;
         16'h9778, 16'h9779, 16'h977a, 16'h977b, 16'h977c, 16'h977d, 16'h977e, 16'h977f 	:	val_out <= 16'h3a47;
         16'h9780, 16'h9781, 16'h9782, 16'h9783, 16'h9784, 16'h9785, 16'h9786, 16'h9787 	:	val_out <= 16'h3a32;
         16'h9788, 16'h9789, 16'h978a, 16'h978b, 16'h978c, 16'h978d, 16'h978e, 16'h978f 	:	val_out <= 16'h3a1d;
         16'h9790, 16'h9791, 16'h9792, 16'h9793, 16'h9794, 16'h9795, 16'h9796, 16'h9797 	:	val_out <= 16'h3a08;
         16'h9798, 16'h9799, 16'h979a, 16'h979b, 16'h979c, 16'h979d, 16'h979e, 16'h979f 	:	val_out <= 16'h39f3;
         16'h97a0, 16'h97a1, 16'h97a2, 16'h97a3, 16'h97a4, 16'h97a5, 16'h97a6, 16'h97a7 	:	val_out <= 16'h39de;
         16'h97a8, 16'h97a9, 16'h97aa, 16'h97ab, 16'h97ac, 16'h97ad, 16'h97ae, 16'h97af 	:	val_out <= 16'h39c9;
         16'h97b0, 16'h97b1, 16'h97b2, 16'h97b3, 16'h97b4, 16'h97b5, 16'h97b6, 16'h97b7 	:	val_out <= 16'h39b4;
         16'h97b8, 16'h97b9, 16'h97ba, 16'h97bb, 16'h97bc, 16'h97bd, 16'h97be, 16'h97bf 	:	val_out <= 16'h399f;
         16'h97c0, 16'h97c1, 16'h97c2, 16'h97c3, 16'h97c4, 16'h97c5, 16'h97c6, 16'h97c7 	:	val_out <= 16'h398a;
         16'h97c8, 16'h97c9, 16'h97ca, 16'h97cb, 16'h97cc, 16'h97cd, 16'h97ce, 16'h97cf 	:	val_out <= 16'h3975;
         16'h97d0, 16'h97d1, 16'h97d2, 16'h97d3, 16'h97d4, 16'h97d5, 16'h97d6, 16'h97d7 	:	val_out <= 16'h3960;
         16'h97d8, 16'h97d9, 16'h97da, 16'h97db, 16'h97dc, 16'h97dd, 16'h97de, 16'h97df 	:	val_out <= 16'h394b;
         16'h97e0, 16'h97e1, 16'h97e2, 16'h97e3, 16'h97e4, 16'h97e5, 16'h97e6, 16'h97e7 	:	val_out <= 16'h3936;
         16'h97e8, 16'h97e9, 16'h97ea, 16'h97eb, 16'h97ec, 16'h97ed, 16'h97ee, 16'h97ef 	:	val_out <= 16'h3921;
         16'h97f0, 16'h97f1, 16'h97f2, 16'h97f3, 16'h97f4, 16'h97f5, 16'h97f6, 16'h97f7 	:	val_out <= 16'h390c;
         16'h97f8, 16'h97f9, 16'h97fa, 16'h97fb, 16'h97fc, 16'h97fd, 16'h97fe, 16'h97ff 	:	val_out <= 16'h38f7;
         16'h9800, 16'h9801, 16'h9802, 16'h9803, 16'h9804, 16'h9805, 16'h9806, 16'h9807 	:	val_out <= 16'h38e3;
         16'h9808, 16'h9809, 16'h980a, 16'h980b, 16'h980c, 16'h980d, 16'h980e, 16'h980f 	:	val_out <= 16'h38ce;
         16'h9810, 16'h9811, 16'h9812, 16'h9813, 16'h9814, 16'h9815, 16'h9816, 16'h9817 	:	val_out <= 16'h38b9;
         16'h9818, 16'h9819, 16'h981a, 16'h981b, 16'h981c, 16'h981d, 16'h981e, 16'h981f 	:	val_out <= 16'h38a4;
         16'h9820, 16'h9821, 16'h9822, 16'h9823, 16'h9824, 16'h9825, 16'h9826, 16'h9827 	:	val_out <= 16'h388f;
         16'h9828, 16'h9829, 16'h982a, 16'h982b, 16'h982c, 16'h982d, 16'h982e, 16'h982f 	:	val_out <= 16'h387a;
         16'h9830, 16'h9831, 16'h9832, 16'h9833, 16'h9834, 16'h9835, 16'h9836, 16'h9837 	:	val_out <= 16'h3865;
         16'h9838, 16'h9839, 16'h983a, 16'h983b, 16'h983c, 16'h983d, 16'h983e, 16'h983f 	:	val_out <= 16'h3851;
         16'h9840, 16'h9841, 16'h9842, 16'h9843, 16'h9844, 16'h9845, 16'h9846, 16'h9847 	:	val_out <= 16'h383c;
         16'h9848, 16'h9849, 16'h984a, 16'h984b, 16'h984c, 16'h984d, 16'h984e, 16'h984f 	:	val_out <= 16'h3827;
         16'h9850, 16'h9851, 16'h9852, 16'h9853, 16'h9854, 16'h9855, 16'h9856, 16'h9857 	:	val_out <= 16'h3812;
         16'h9858, 16'h9859, 16'h985a, 16'h985b, 16'h985c, 16'h985d, 16'h985e, 16'h985f 	:	val_out <= 16'h37fd;
         16'h9860, 16'h9861, 16'h9862, 16'h9863, 16'h9864, 16'h9865, 16'h9866, 16'h9867 	:	val_out <= 16'h37e9;
         16'h9868, 16'h9869, 16'h986a, 16'h986b, 16'h986c, 16'h986d, 16'h986e, 16'h986f 	:	val_out <= 16'h37d4;
         16'h9870, 16'h9871, 16'h9872, 16'h9873, 16'h9874, 16'h9875, 16'h9876, 16'h9877 	:	val_out <= 16'h37bf;
         16'h9878, 16'h9879, 16'h987a, 16'h987b, 16'h987c, 16'h987d, 16'h987e, 16'h987f 	:	val_out <= 16'h37aa;
         16'h9880, 16'h9881, 16'h9882, 16'h9883, 16'h9884, 16'h9885, 16'h9886, 16'h9887 	:	val_out <= 16'h3796;
         16'h9888, 16'h9889, 16'h988a, 16'h988b, 16'h988c, 16'h988d, 16'h988e, 16'h988f 	:	val_out <= 16'h3781;
         16'h9890, 16'h9891, 16'h9892, 16'h9893, 16'h9894, 16'h9895, 16'h9896, 16'h9897 	:	val_out <= 16'h376c;
         16'h9898, 16'h9899, 16'h989a, 16'h989b, 16'h989c, 16'h989d, 16'h989e, 16'h989f 	:	val_out <= 16'h3757;
         16'h98a0, 16'h98a1, 16'h98a2, 16'h98a3, 16'h98a4, 16'h98a5, 16'h98a6, 16'h98a7 	:	val_out <= 16'h3743;
         16'h98a8, 16'h98a9, 16'h98aa, 16'h98ab, 16'h98ac, 16'h98ad, 16'h98ae, 16'h98af 	:	val_out <= 16'h372e;
         16'h98b0, 16'h98b1, 16'h98b2, 16'h98b3, 16'h98b4, 16'h98b5, 16'h98b6, 16'h98b7 	:	val_out <= 16'h3719;
         16'h98b8, 16'h98b9, 16'h98ba, 16'h98bb, 16'h98bc, 16'h98bd, 16'h98be, 16'h98bf 	:	val_out <= 16'h3705;
         16'h98c0, 16'h98c1, 16'h98c2, 16'h98c3, 16'h98c4, 16'h98c5, 16'h98c6, 16'h98c7 	:	val_out <= 16'h36f0;
         16'h98c8, 16'h98c9, 16'h98ca, 16'h98cb, 16'h98cc, 16'h98cd, 16'h98ce, 16'h98cf 	:	val_out <= 16'h36dc;
         16'h98d0, 16'h98d1, 16'h98d2, 16'h98d3, 16'h98d4, 16'h98d5, 16'h98d6, 16'h98d7 	:	val_out <= 16'h36c7;
         16'h98d8, 16'h98d9, 16'h98da, 16'h98db, 16'h98dc, 16'h98dd, 16'h98de, 16'h98df 	:	val_out <= 16'h36b2;
         16'h98e0, 16'h98e1, 16'h98e2, 16'h98e3, 16'h98e4, 16'h98e5, 16'h98e6, 16'h98e7 	:	val_out <= 16'h369e;
         16'h98e8, 16'h98e9, 16'h98ea, 16'h98eb, 16'h98ec, 16'h98ed, 16'h98ee, 16'h98ef 	:	val_out <= 16'h3689;
         16'h98f0, 16'h98f1, 16'h98f2, 16'h98f3, 16'h98f4, 16'h98f5, 16'h98f6, 16'h98f7 	:	val_out <= 16'h3675;
         16'h98f8, 16'h98f9, 16'h98fa, 16'h98fb, 16'h98fc, 16'h98fd, 16'h98fe, 16'h98ff 	:	val_out <= 16'h3660;
         16'h9900, 16'h9901, 16'h9902, 16'h9903, 16'h9904, 16'h9905, 16'h9906, 16'h9907 	:	val_out <= 16'h364b;
         16'h9908, 16'h9909, 16'h990a, 16'h990b, 16'h990c, 16'h990d, 16'h990e, 16'h990f 	:	val_out <= 16'h3637;
         16'h9910, 16'h9911, 16'h9912, 16'h9913, 16'h9914, 16'h9915, 16'h9916, 16'h9917 	:	val_out <= 16'h3622;
         16'h9918, 16'h9919, 16'h991a, 16'h991b, 16'h991c, 16'h991d, 16'h991e, 16'h991f 	:	val_out <= 16'h360e;
         16'h9920, 16'h9921, 16'h9922, 16'h9923, 16'h9924, 16'h9925, 16'h9926, 16'h9927 	:	val_out <= 16'h35f9;
         16'h9928, 16'h9929, 16'h992a, 16'h992b, 16'h992c, 16'h992d, 16'h992e, 16'h992f 	:	val_out <= 16'h35e5;
         16'h9930, 16'h9931, 16'h9932, 16'h9933, 16'h9934, 16'h9935, 16'h9936, 16'h9937 	:	val_out <= 16'h35d0;
         16'h9938, 16'h9939, 16'h993a, 16'h993b, 16'h993c, 16'h993d, 16'h993e, 16'h993f 	:	val_out <= 16'h35bc;
         16'h9940, 16'h9941, 16'h9942, 16'h9943, 16'h9944, 16'h9945, 16'h9946, 16'h9947 	:	val_out <= 16'h35a7;
         16'h9948, 16'h9949, 16'h994a, 16'h994b, 16'h994c, 16'h994d, 16'h994e, 16'h994f 	:	val_out <= 16'h3593;
         16'h9950, 16'h9951, 16'h9952, 16'h9953, 16'h9954, 16'h9955, 16'h9956, 16'h9957 	:	val_out <= 16'h357e;
         16'h9958, 16'h9959, 16'h995a, 16'h995b, 16'h995c, 16'h995d, 16'h995e, 16'h995f 	:	val_out <= 16'h356a;
         16'h9960, 16'h9961, 16'h9962, 16'h9963, 16'h9964, 16'h9965, 16'h9966, 16'h9967 	:	val_out <= 16'h3556;
         16'h9968, 16'h9969, 16'h996a, 16'h996b, 16'h996c, 16'h996d, 16'h996e, 16'h996f 	:	val_out <= 16'h3541;
         16'h9970, 16'h9971, 16'h9972, 16'h9973, 16'h9974, 16'h9975, 16'h9976, 16'h9977 	:	val_out <= 16'h352d;
         16'h9978, 16'h9979, 16'h997a, 16'h997b, 16'h997c, 16'h997d, 16'h997e, 16'h997f 	:	val_out <= 16'h3518;
         16'h9980, 16'h9981, 16'h9982, 16'h9983, 16'h9984, 16'h9985, 16'h9986, 16'h9987 	:	val_out <= 16'h3504;
         16'h9988, 16'h9989, 16'h998a, 16'h998b, 16'h998c, 16'h998d, 16'h998e, 16'h998f 	:	val_out <= 16'h34f0;
         16'h9990, 16'h9991, 16'h9992, 16'h9993, 16'h9994, 16'h9995, 16'h9996, 16'h9997 	:	val_out <= 16'h34db;
         16'h9998, 16'h9999, 16'h999a, 16'h999b, 16'h999c, 16'h999d, 16'h999e, 16'h999f 	:	val_out <= 16'h34c7;
         16'h99a0, 16'h99a1, 16'h99a2, 16'h99a3, 16'h99a4, 16'h99a5, 16'h99a6, 16'h99a7 	:	val_out <= 16'h34b3;
         16'h99a8, 16'h99a9, 16'h99aa, 16'h99ab, 16'h99ac, 16'h99ad, 16'h99ae, 16'h99af 	:	val_out <= 16'h349e;
         16'h99b0, 16'h99b1, 16'h99b2, 16'h99b3, 16'h99b4, 16'h99b5, 16'h99b6, 16'h99b7 	:	val_out <= 16'h348a;
         16'h99b8, 16'h99b9, 16'h99ba, 16'h99bb, 16'h99bc, 16'h99bd, 16'h99be, 16'h99bf 	:	val_out <= 16'h3476;
         16'h99c0, 16'h99c1, 16'h99c2, 16'h99c3, 16'h99c4, 16'h99c5, 16'h99c6, 16'h99c7 	:	val_out <= 16'h3461;
         16'h99c8, 16'h99c9, 16'h99ca, 16'h99cb, 16'h99cc, 16'h99cd, 16'h99ce, 16'h99cf 	:	val_out <= 16'h344d;
         16'h99d0, 16'h99d1, 16'h99d2, 16'h99d3, 16'h99d4, 16'h99d5, 16'h99d6, 16'h99d7 	:	val_out <= 16'h3439;
         16'h99d8, 16'h99d9, 16'h99da, 16'h99db, 16'h99dc, 16'h99dd, 16'h99de, 16'h99df 	:	val_out <= 16'h3425;
         16'h99e0, 16'h99e1, 16'h99e2, 16'h99e3, 16'h99e4, 16'h99e5, 16'h99e6, 16'h99e7 	:	val_out <= 16'h3410;
         16'h99e8, 16'h99e9, 16'h99ea, 16'h99eb, 16'h99ec, 16'h99ed, 16'h99ee, 16'h99ef 	:	val_out <= 16'h33fc;
         16'h99f0, 16'h99f1, 16'h99f2, 16'h99f3, 16'h99f4, 16'h99f5, 16'h99f6, 16'h99f7 	:	val_out <= 16'h33e8;
         16'h99f8, 16'h99f9, 16'h99fa, 16'h99fb, 16'h99fc, 16'h99fd, 16'h99fe, 16'h99ff 	:	val_out <= 16'h33d4;
         16'h9a00, 16'h9a01, 16'h9a02, 16'h9a03, 16'h9a04, 16'h9a05, 16'h9a06, 16'h9a07 	:	val_out <= 16'h33c0;
         16'h9a08, 16'h9a09, 16'h9a0a, 16'h9a0b, 16'h9a0c, 16'h9a0d, 16'h9a0e, 16'h9a0f 	:	val_out <= 16'h33ab;
         16'h9a10, 16'h9a11, 16'h9a12, 16'h9a13, 16'h9a14, 16'h9a15, 16'h9a16, 16'h9a17 	:	val_out <= 16'h3397;
         16'h9a18, 16'h9a19, 16'h9a1a, 16'h9a1b, 16'h9a1c, 16'h9a1d, 16'h9a1e, 16'h9a1f 	:	val_out <= 16'h3383;
         16'h9a20, 16'h9a21, 16'h9a22, 16'h9a23, 16'h9a24, 16'h9a25, 16'h9a26, 16'h9a27 	:	val_out <= 16'h336f;
         16'h9a28, 16'h9a29, 16'h9a2a, 16'h9a2b, 16'h9a2c, 16'h9a2d, 16'h9a2e, 16'h9a2f 	:	val_out <= 16'h335b;
         16'h9a30, 16'h9a31, 16'h9a32, 16'h9a33, 16'h9a34, 16'h9a35, 16'h9a36, 16'h9a37 	:	val_out <= 16'h3347;
         16'h9a38, 16'h9a39, 16'h9a3a, 16'h9a3b, 16'h9a3c, 16'h9a3d, 16'h9a3e, 16'h9a3f 	:	val_out <= 16'h3333;
         16'h9a40, 16'h9a41, 16'h9a42, 16'h9a43, 16'h9a44, 16'h9a45, 16'h9a46, 16'h9a47 	:	val_out <= 16'h331e;
         16'h9a48, 16'h9a49, 16'h9a4a, 16'h9a4b, 16'h9a4c, 16'h9a4d, 16'h9a4e, 16'h9a4f 	:	val_out <= 16'h330a;
         16'h9a50, 16'h9a51, 16'h9a52, 16'h9a53, 16'h9a54, 16'h9a55, 16'h9a56, 16'h9a57 	:	val_out <= 16'h32f6;
         16'h9a58, 16'h9a59, 16'h9a5a, 16'h9a5b, 16'h9a5c, 16'h9a5d, 16'h9a5e, 16'h9a5f 	:	val_out <= 16'h32e2;
         16'h9a60, 16'h9a61, 16'h9a62, 16'h9a63, 16'h9a64, 16'h9a65, 16'h9a66, 16'h9a67 	:	val_out <= 16'h32ce;
         16'h9a68, 16'h9a69, 16'h9a6a, 16'h9a6b, 16'h9a6c, 16'h9a6d, 16'h9a6e, 16'h9a6f 	:	val_out <= 16'h32ba;
         16'h9a70, 16'h9a71, 16'h9a72, 16'h9a73, 16'h9a74, 16'h9a75, 16'h9a76, 16'h9a77 	:	val_out <= 16'h32a6;
         16'h9a78, 16'h9a79, 16'h9a7a, 16'h9a7b, 16'h9a7c, 16'h9a7d, 16'h9a7e, 16'h9a7f 	:	val_out <= 16'h3292;
         16'h9a80, 16'h9a81, 16'h9a82, 16'h9a83, 16'h9a84, 16'h9a85, 16'h9a86, 16'h9a87 	:	val_out <= 16'h327e;
         16'h9a88, 16'h9a89, 16'h9a8a, 16'h9a8b, 16'h9a8c, 16'h9a8d, 16'h9a8e, 16'h9a8f 	:	val_out <= 16'h326a;
         16'h9a90, 16'h9a91, 16'h9a92, 16'h9a93, 16'h9a94, 16'h9a95, 16'h9a96, 16'h9a97 	:	val_out <= 16'h3256;
         16'h9a98, 16'h9a99, 16'h9a9a, 16'h9a9b, 16'h9a9c, 16'h9a9d, 16'h9a9e, 16'h9a9f 	:	val_out <= 16'h3242;
         16'h9aa0, 16'h9aa1, 16'h9aa2, 16'h9aa3, 16'h9aa4, 16'h9aa5, 16'h9aa6, 16'h9aa7 	:	val_out <= 16'h322e;
         16'h9aa8, 16'h9aa9, 16'h9aaa, 16'h9aab, 16'h9aac, 16'h9aad, 16'h9aae, 16'h9aaf 	:	val_out <= 16'h321a;
         16'h9ab0, 16'h9ab1, 16'h9ab2, 16'h9ab3, 16'h9ab4, 16'h9ab5, 16'h9ab6, 16'h9ab7 	:	val_out <= 16'h3206;
         16'h9ab8, 16'h9ab9, 16'h9aba, 16'h9abb, 16'h9abc, 16'h9abd, 16'h9abe, 16'h9abf 	:	val_out <= 16'h31f2;
         16'h9ac0, 16'h9ac1, 16'h9ac2, 16'h9ac3, 16'h9ac4, 16'h9ac5, 16'h9ac6, 16'h9ac7 	:	val_out <= 16'h31de;
         16'h9ac8, 16'h9ac9, 16'h9aca, 16'h9acb, 16'h9acc, 16'h9acd, 16'h9ace, 16'h9acf 	:	val_out <= 16'h31cb;
         16'h9ad0, 16'h9ad1, 16'h9ad2, 16'h9ad3, 16'h9ad4, 16'h9ad5, 16'h9ad6, 16'h9ad7 	:	val_out <= 16'h31b7;
         16'h9ad8, 16'h9ad9, 16'h9ada, 16'h9adb, 16'h9adc, 16'h9add, 16'h9ade, 16'h9adf 	:	val_out <= 16'h31a3;
         16'h9ae0, 16'h9ae1, 16'h9ae2, 16'h9ae3, 16'h9ae4, 16'h9ae5, 16'h9ae6, 16'h9ae7 	:	val_out <= 16'h318f;
         16'h9ae8, 16'h9ae9, 16'h9aea, 16'h9aeb, 16'h9aec, 16'h9aed, 16'h9aee, 16'h9aef 	:	val_out <= 16'h317b;
         16'h9af0, 16'h9af1, 16'h9af2, 16'h9af3, 16'h9af4, 16'h9af5, 16'h9af6, 16'h9af7 	:	val_out <= 16'h3167;
         16'h9af8, 16'h9af9, 16'h9afa, 16'h9afb, 16'h9afc, 16'h9afd, 16'h9afe, 16'h9aff 	:	val_out <= 16'h3153;
         16'h9b00, 16'h9b01, 16'h9b02, 16'h9b03, 16'h9b04, 16'h9b05, 16'h9b06, 16'h9b07 	:	val_out <= 16'h3140;
         16'h9b08, 16'h9b09, 16'h9b0a, 16'h9b0b, 16'h9b0c, 16'h9b0d, 16'h9b0e, 16'h9b0f 	:	val_out <= 16'h312c;
         16'h9b10, 16'h9b11, 16'h9b12, 16'h9b13, 16'h9b14, 16'h9b15, 16'h9b16, 16'h9b17 	:	val_out <= 16'h3118;
         16'h9b18, 16'h9b19, 16'h9b1a, 16'h9b1b, 16'h9b1c, 16'h9b1d, 16'h9b1e, 16'h9b1f 	:	val_out <= 16'h3104;
         16'h9b20, 16'h9b21, 16'h9b22, 16'h9b23, 16'h9b24, 16'h9b25, 16'h9b26, 16'h9b27 	:	val_out <= 16'h30f0;
         16'h9b28, 16'h9b29, 16'h9b2a, 16'h9b2b, 16'h9b2c, 16'h9b2d, 16'h9b2e, 16'h9b2f 	:	val_out <= 16'h30dd;
         16'h9b30, 16'h9b31, 16'h9b32, 16'h9b33, 16'h9b34, 16'h9b35, 16'h9b36, 16'h9b37 	:	val_out <= 16'h30c9;
         16'h9b38, 16'h9b39, 16'h9b3a, 16'h9b3b, 16'h9b3c, 16'h9b3d, 16'h9b3e, 16'h9b3f 	:	val_out <= 16'h30b5;
         16'h9b40, 16'h9b41, 16'h9b42, 16'h9b43, 16'h9b44, 16'h9b45, 16'h9b46, 16'h9b47 	:	val_out <= 16'h30a1;
         16'h9b48, 16'h9b49, 16'h9b4a, 16'h9b4b, 16'h9b4c, 16'h9b4d, 16'h9b4e, 16'h9b4f 	:	val_out <= 16'h308e;
         16'h9b50, 16'h9b51, 16'h9b52, 16'h9b53, 16'h9b54, 16'h9b55, 16'h9b56, 16'h9b57 	:	val_out <= 16'h307a;
         16'h9b58, 16'h9b59, 16'h9b5a, 16'h9b5b, 16'h9b5c, 16'h9b5d, 16'h9b5e, 16'h9b5f 	:	val_out <= 16'h3066;
         16'h9b60, 16'h9b61, 16'h9b62, 16'h9b63, 16'h9b64, 16'h9b65, 16'h9b66, 16'h9b67 	:	val_out <= 16'h3053;
         16'h9b68, 16'h9b69, 16'h9b6a, 16'h9b6b, 16'h9b6c, 16'h9b6d, 16'h9b6e, 16'h9b6f 	:	val_out <= 16'h303f;
         16'h9b70, 16'h9b71, 16'h9b72, 16'h9b73, 16'h9b74, 16'h9b75, 16'h9b76, 16'h9b77 	:	val_out <= 16'h302b;
         16'h9b78, 16'h9b79, 16'h9b7a, 16'h9b7b, 16'h9b7c, 16'h9b7d, 16'h9b7e, 16'h9b7f 	:	val_out <= 16'h3018;
         16'h9b80, 16'h9b81, 16'h9b82, 16'h9b83, 16'h9b84, 16'h9b85, 16'h9b86, 16'h9b87 	:	val_out <= 16'h3004;
         16'h9b88, 16'h9b89, 16'h9b8a, 16'h9b8b, 16'h9b8c, 16'h9b8d, 16'h9b8e, 16'h9b8f 	:	val_out <= 16'h2ff0;
         16'h9b90, 16'h9b91, 16'h9b92, 16'h9b93, 16'h9b94, 16'h9b95, 16'h9b96, 16'h9b97 	:	val_out <= 16'h2fdd;
         16'h9b98, 16'h9b99, 16'h9b9a, 16'h9b9b, 16'h9b9c, 16'h9b9d, 16'h9b9e, 16'h9b9f 	:	val_out <= 16'h2fc9;
         16'h9ba0, 16'h9ba1, 16'h9ba2, 16'h9ba3, 16'h9ba4, 16'h9ba5, 16'h9ba6, 16'h9ba7 	:	val_out <= 16'h2fb6;
         16'h9ba8, 16'h9ba9, 16'h9baa, 16'h9bab, 16'h9bac, 16'h9bad, 16'h9bae, 16'h9baf 	:	val_out <= 16'h2fa2;
         16'h9bb0, 16'h9bb1, 16'h9bb2, 16'h9bb3, 16'h9bb4, 16'h9bb5, 16'h9bb6, 16'h9bb7 	:	val_out <= 16'h2f8f;
         16'h9bb8, 16'h9bb9, 16'h9bba, 16'h9bbb, 16'h9bbc, 16'h9bbd, 16'h9bbe, 16'h9bbf 	:	val_out <= 16'h2f7b;
         16'h9bc0, 16'h9bc1, 16'h9bc2, 16'h9bc3, 16'h9bc4, 16'h9bc5, 16'h9bc6, 16'h9bc7 	:	val_out <= 16'h2f68;
         16'h9bc8, 16'h9bc9, 16'h9bca, 16'h9bcb, 16'h9bcc, 16'h9bcd, 16'h9bce, 16'h9bcf 	:	val_out <= 16'h2f54;
         16'h9bd0, 16'h9bd1, 16'h9bd2, 16'h9bd3, 16'h9bd4, 16'h9bd5, 16'h9bd6, 16'h9bd7 	:	val_out <= 16'h2f40;
         16'h9bd8, 16'h9bd9, 16'h9bda, 16'h9bdb, 16'h9bdc, 16'h9bdd, 16'h9bde, 16'h9bdf 	:	val_out <= 16'h2f2d;
         16'h9be0, 16'h9be1, 16'h9be2, 16'h9be3, 16'h9be4, 16'h9be5, 16'h9be6, 16'h9be7 	:	val_out <= 16'h2f1a;
         16'h9be8, 16'h9be9, 16'h9bea, 16'h9beb, 16'h9bec, 16'h9bed, 16'h9bee, 16'h9bef 	:	val_out <= 16'h2f06;
         16'h9bf0, 16'h9bf1, 16'h9bf2, 16'h9bf3, 16'h9bf4, 16'h9bf5, 16'h9bf6, 16'h9bf7 	:	val_out <= 16'h2ef3;
         16'h9bf8, 16'h9bf9, 16'h9bfa, 16'h9bfb, 16'h9bfc, 16'h9bfd, 16'h9bfe, 16'h9bff 	:	val_out <= 16'h2edf;
         16'h9c00, 16'h9c01, 16'h9c02, 16'h9c03, 16'h9c04, 16'h9c05, 16'h9c06, 16'h9c07 	:	val_out <= 16'h2ecc;
         16'h9c08, 16'h9c09, 16'h9c0a, 16'h9c0b, 16'h9c0c, 16'h9c0d, 16'h9c0e, 16'h9c0f 	:	val_out <= 16'h2eb8;
         16'h9c10, 16'h9c11, 16'h9c12, 16'h9c13, 16'h9c14, 16'h9c15, 16'h9c16, 16'h9c17 	:	val_out <= 16'h2ea5;
         16'h9c18, 16'h9c19, 16'h9c1a, 16'h9c1b, 16'h9c1c, 16'h9c1d, 16'h9c1e, 16'h9c1f 	:	val_out <= 16'h2e91;
         16'h9c20, 16'h9c21, 16'h9c22, 16'h9c23, 16'h9c24, 16'h9c25, 16'h9c26, 16'h9c27 	:	val_out <= 16'h2e7e;
         16'h9c28, 16'h9c29, 16'h9c2a, 16'h9c2b, 16'h9c2c, 16'h9c2d, 16'h9c2e, 16'h9c2f 	:	val_out <= 16'h2e6b;
         16'h9c30, 16'h9c31, 16'h9c32, 16'h9c33, 16'h9c34, 16'h9c35, 16'h9c36, 16'h9c37 	:	val_out <= 16'h2e57;
         16'h9c38, 16'h9c39, 16'h9c3a, 16'h9c3b, 16'h9c3c, 16'h9c3d, 16'h9c3e, 16'h9c3f 	:	val_out <= 16'h2e44;
         16'h9c40, 16'h9c41, 16'h9c42, 16'h9c43, 16'h9c44, 16'h9c45, 16'h9c46, 16'h9c47 	:	val_out <= 16'h2e31;
         16'h9c48, 16'h9c49, 16'h9c4a, 16'h9c4b, 16'h9c4c, 16'h9c4d, 16'h9c4e, 16'h9c4f 	:	val_out <= 16'h2e1d;
         16'h9c50, 16'h9c51, 16'h9c52, 16'h9c53, 16'h9c54, 16'h9c55, 16'h9c56, 16'h9c57 	:	val_out <= 16'h2e0a;
         16'h9c58, 16'h9c59, 16'h9c5a, 16'h9c5b, 16'h9c5c, 16'h9c5d, 16'h9c5e, 16'h9c5f 	:	val_out <= 16'h2df7;
         16'h9c60, 16'h9c61, 16'h9c62, 16'h9c63, 16'h9c64, 16'h9c65, 16'h9c66, 16'h9c67 	:	val_out <= 16'h2de3;
         16'h9c68, 16'h9c69, 16'h9c6a, 16'h9c6b, 16'h9c6c, 16'h9c6d, 16'h9c6e, 16'h9c6f 	:	val_out <= 16'h2dd0;
         16'h9c70, 16'h9c71, 16'h9c72, 16'h9c73, 16'h9c74, 16'h9c75, 16'h9c76, 16'h9c77 	:	val_out <= 16'h2dbd;
         16'h9c78, 16'h9c79, 16'h9c7a, 16'h9c7b, 16'h9c7c, 16'h9c7d, 16'h9c7e, 16'h9c7f 	:	val_out <= 16'h2daa;
         16'h9c80, 16'h9c81, 16'h9c82, 16'h9c83, 16'h9c84, 16'h9c85, 16'h9c86, 16'h9c87 	:	val_out <= 16'h2d96;
         16'h9c88, 16'h9c89, 16'h9c8a, 16'h9c8b, 16'h9c8c, 16'h9c8d, 16'h9c8e, 16'h9c8f 	:	val_out <= 16'h2d83;
         16'h9c90, 16'h9c91, 16'h9c92, 16'h9c93, 16'h9c94, 16'h9c95, 16'h9c96, 16'h9c97 	:	val_out <= 16'h2d70;
         16'h9c98, 16'h9c99, 16'h9c9a, 16'h9c9b, 16'h9c9c, 16'h9c9d, 16'h9c9e, 16'h9c9f 	:	val_out <= 16'h2d5d;
         16'h9ca0, 16'h9ca1, 16'h9ca2, 16'h9ca3, 16'h9ca4, 16'h9ca5, 16'h9ca6, 16'h9ca7 	:	val_out <= 16'h2d4a;
         16'h9ca8, 16'h9ca9, 16'h9caa, 16'h9cab, 16'h9cac, 16'h9cad, 16'h9cae, 16'h9caf 	:	val_out <= 16'h2d36;
         16'h9cb0, 16'h9cb1, 16'h9cb2, 16'h9cb3, 16'h9cb4, 16'h9cb5, 16'h9cb6, 16'h9cb7 	:	val_out <= 16'h2d23;
         16'h9cb8, 16'h9cb9, 16'h9cba, 16'h9cbb, 16'h9cbc, 16'h9cbd, 16'h9cbe, 16'h9cbf 	:	val_out <= 16'h2d10;
         16'h9cc0, 16'h9cc1, 16'h9cc2, 16'h9cc3, 16'h9cc4, 16'h9cc5, 16'h9cc6, 16'h9cc7 	:	val_out <= 16'h2cfd;
         16'h9cc8, 16'h9cc9, 16'h9cca, 16'h9ccb, 16'h9ccc, 16'h9ccd, 16'h9cce, 16'h9ccf 	:	val_out <= 16'h2cea;
         16'h9cd0, 16'h9cd1, 16'h9cd2, 16'h9cd3, 16'h9cd4, 16'h9cd5, 16'h9cd6, 16'h9cd7 	:	val_out <= 16'h2cd7;
         16'h9cd8, 16'h9cd9, 16'h9cda, 16'h9cdb, 16'h9cdc, 16'h9cdd, 16'h9cde, 16'h9cdf 	:	val_out <= 16'h2cc4;
         16'h9ce0, 16'h9ce1, 16'h9ce2, 16'h9ce3, 16'h9ce4, 16'h9ce5, 16'h9ce6, 16'h9ce7 	:	val_out <= 16'h2cb1;
         16'h9ce8, 16'h9ce9, 16'h9cea, 16'h9ceb, 16'h9cec, 16'h9ced, 16'h9cee, 16'h9cef 	:	val_out <= 16'h2c9d;
         16'h9cf0, 16'h9cf1, 16'h9cf2, 16'h9cf3, 16'h9cf4, 16'h9cf5, 16'h9cf6, 16'h9cf7 	:	val_out <= 16'h2c8a;
         16'h9cf8, 16'h9cf9, 16'h9cfa, 16'h9cfb, 16'h9cfc, 16'h9cfd, 16'h9cfe, 16'h9cff 	:	val_out <= 16'h2c77;
         16'h9d00, 16'h9d01, 16'h9d02, 16'h9d03, 16'h9d04, 16'h9d05, 16'h9d06, 16'h9d07 	:	val_out <= 16'h2c64;
         16'h9d08, 16'h9d09, 16'h9d0a, 16'h9d0b, 16'h9d0c, 16'h9d0d, 16'h9d0e, 16'h9d0f 	:	val_out <= 16'h2c51;
         16'h9d10, 16'h9d11, 16'h9d12, 16'h9d13, 16'h9d14, 16'h9d15, 16'h9d16, 16'h9d17 	:	val_out <= 16'h2c3e;
         16'h9d18, 16'h9d19, 16'h9d1a, 16'h9d1b, 16'h9d1c, 16'h9d1d, 16'h9d1e, 16'h9d1f 	:	val_out <= 16'h2c2b;
         16'h9d20, 16'h9d21, 16'h9d22, 16'h9d23, 16'h9d24, 16'h9d25, 16'h9d26, 16'h9d27 	:	val_out <= 16'h2c18;
         16'h9d28, 16'h9d29, 16'h9d2a, 16'h9d2b, 16'h9d2c, 16'h9d2d, 16'h9d2e, 16'h9d2f 	:	val_out <= 16'h2c05;
         16'h9d30, 16'h9d31, 16'h9d32, 16'h9d33, 16'h9d34, 16'h9d35, 16'h9d36, 16'h9d37 	:	val_out <= 16'h2bf2;
         16'h9d38, 16'h9d39, 16'h9d3a, 16'h9d3b, 16'h9d3c, 16'h9d3d, 16'h9d3e, 16'h9d3f 	:	val_out <= 16'h2bdf;
         16'h9d40, 16'h9d41, 16'h9d42, 16'h9d43, 16'h9d44, 16'h9d45, 16'h9d46, 16'h9d47 	:	val_out <= 16'h2bcc;
         16'h9d48, 16'h9d49, 16'h9d4a, 16'h9d4b, 16'h9d4c, 16'h9d4d, 16'h9d4e, 16'h9d4f 	:	val_out <= 16'h2bba;
         16'h9d50, 16'h9d51, 16'h9d52, 16'h9d53, 16'h9d54, 16'h9d55, 16'h9d56, 16'h9d57 	:	val_out <= 16'h2ba7;
         16'h9d58, 16'h9d59, 16'h9d5a, 16'h9d5b, 16'h9d5c, 16'h9d5d, 16'h9d5e, 16'h9d5f 	:	val_out <= 16'h2b94;
         16'h9d60, 16'h9d61, 16'h9d62, 16'h9d63, 16'h9d64, 16'h9d65, 16'h9d66, 16'h9d67 	:	val_out <= 16'h2b81;
         16'h9d68, 16'h9d69, 16'h9d6a, 16'h9d6b, 16'h9d6c, 16'h9d6d, 16'h9d6e, 16'h9d6f 	:	val_out <= 16'h2b6e;
         16'h9d70, 16'h9d71, 16'h9d72, 16'h9d73, 16'h9d74, 16'h9d75, 16'h9d76, 16'h9d77 	:	val_out <= 16'h2b5b;
         16'h9d78, 16'h9d79, 16'h9d7a, 16'h9d7b, 16'h9d7c, 16'h9d7d, 16'h9d7e, 16'h9d7f 	:	val_out <= 16'h2b48;
         16'h9d80, 16'h9d81, 16'h9d82, 16'h9d83, 16'h9d84, 16'h9d85, 16'h9d86, 16'h9d87 	:	val_out <= 16'h2b35;
         16'h9d88, 16'h9d89, 16'h9d8a, 16'h9d8b, 16'h9d8c, 16'h9d8d, 16'h9d8e, 16'h9d8f 	:	val_out <= 16'h2b23;
         16'h9d90, 16'h9d91, 16'h9d92, 16'h9d93, 16'h9d94, 16'h9d95, 16'h9d96, 16'h9d97 	:	val_out <= 16'h2b10;
         16'h9d98, 16'h9d99, 16'h9d9a, 16'h9d9b, 16'h9d9c, 16'h9d9d, 16'h9d9e, 16'h9d9f 	:	val_out <= 16'h2afd;
         16'h9da0, 16'h9da1, 16'h9da2, 16'h9da3, 16'h9da4, 16'h9da5, 16'h9da6, 16'h9da7 	:	val_out <= 16'h2aea;
         16'h9da8, 16'h9da9, 16'h9daa, 16'h9dab, 16'h9dac, 16'h9dad, 16'h9dae, 16'h9daf 	:	val_out <= 16'h2ad7;
         16'h9db0, 16'h9db1, 16'h9db2, 16'h9db3, 16'h9db4, 16'h9db5, 16'h9db6, 16'h9db7 	:	val_out <= 16'h2ac5;
         16'h9db8, 16'h9db9, 16'h9dba, 16'h9dbb, 16'h9dbc, 16'h9dbd, 16'h9dbe, 16'h9dbf 	:	val_out <= 16'h2ab2;
         16'h9dc0, 16'h9dc1, 16'h9dc2, 16'h9dc3, 16'h9dc4, 16'h9dc5, 16'h9dc6, 16'h9dc7 	:	val_out <= 16'h2a9f;
         16'h9dc8, 16'h9dc9, 16'h9dca, 16'h9dcb, 16'h9dcc, 16'h9dcd, 16'h9dce, 16'h9dcf 	:	val_out <= 16'h2a8d;
         16'h9dd0, 16'h9dd1, 16'h9dd2, 16'h9dd3, 16'h9dd4, 16'h9dd5, 16'h9dd6, 16'h9dd7 	:	val_out <= 16'h2a7a;
         16'h9dd8, 16'h9dd9, 16'h9dda, 16'h9ddb, 16'h9ddc, 16'h9ddd, 16'h9dde, 16'h9ddf 	:	val_out <= 16'h2a67;
         16'h9de0, 16'h9de1, 16'h9de2, 16'h9de3, 16'h9de4, 16'h9de5, 16'h9de6, 16'h9de7 	:	val_out <= 16'h2a54;
         16'h9de8, 16'h9de9, 16'h9dea, 16'h9deb, 16'h9dec, 16'h9ded, 16'h9dee, 16'h9def 	:	val_out <= 16'h2a42;
         16'h9df0, 16'h9df1, 16'h9df2, 16'h9df3, 16'h9df4, 16'h9df5, 16'h9df6, 16'h9df7 	:	val_out <= 16'h2a2f;
         16'h9df8, 16'h9df9, 16'h9dfa, 16'h9dfb, 16'h9dfc, 16'h9dfd, 16'h9dfe, 16'h9dff 	:	val_out <= 16'h2a1c;
         16'h9e00, 16'h9e01, 16'h9e02, 16'h9e03, 16'h9e04, 16'h9e05, 16'h9e06, 16'h9e07 	:	val_out <= 16'h2a0a;
         16'h9e08, 16'h9e09, 16'h9e0a, 16'h9e0b, 16'h9e0c, 16'h9e0d, 16'h9e0e, 16'h9e0f 	:	val_out <= 16'h29f7;
         16'h9e10, 16'h9e11, 16'h9e12, 16'h9e13, 16'h9e14, 16'h9e15, 16'h9e16, 16'h9e17 	:	val_out <= 16'h29e5;
         16'h9e18, 16'h9e19, 16'h9e1a, 16'h9e1b, 16'h9e1c, 16'h9e1d, 16'h9e1e, 16'h9e1f 	:	val_out <= 16'h29d2;
         16'h9e20, 16'h9e21, 16'h9e22, 16'h9e23, 16'h9e24, 16'h9e25, 16'h9e26, 16'h9e27 	:	val_out <= 16'h29bf;
         16'h9e28, 16'h9e29, 16'h9e2a, 16'h9e2b, 16'h9e2c, 16'h9e2d, 16'h9e2e, 16'h9e2f 	:	val_out <= 16'h29ad;
         16'h9e30, 16'h9e31, 16'h9e32, 16'h9e33, 16'h9e34, 16'h9e35, 16'h9e36, 16'h9e37 	:	val_out <= 16'h299a;
         16'h9e38, 16'h9e39, 16'h9e3a, 16'h9e3b, 16'h9e3c, 16'h9e3d, 16'h9e3e, 16'h9e3f 	:	val_out <= 16'h2988;
         16'h9e40, 16'h9e41, 16'h9e42, 16'h9e43, 16'h9e44, 16'h9e45, 16'h9e46, 16'h9e47 	:	val_out <= 16'h2975;
         16'h9e48, 16'h9e49, 16'h9e4a, 16'h9e4b, 16'h9e4c, 16'h9e4d, 16'h9e4e, 16'h9e4f 	:	val_out <= 16'h2963;
         16'h9e50, 16'h9e51, 16'h9e52, 16'h9e53, 16'h9e54, 16'h9e55, 16'h9e56, 16'h9e57 	:	val_out <= 16'h2950;
         16'h9e58, 16'h9e59, 16'h9e5a, 16'h9e5b, 16'h9e5c, 16'h9e5d, 16'h9e5e, 16'h9e5f 	:	val_out <= 16'h293e;
         16'h9e60, 16'h9e61, 16'h9e62, 16'h9e63, 16'h9e64, 16'h9e65, 16'h9e66, 16'h9e67 	:	val_out <= 16'h292b;
         16'h9e68, 16'h9e69, 16'h9e6a, 16'h9e6b, 16'h9e6c, 16'h9e6d, 16'h9e6e, 16'h9e6f 	:	val_out <= 16'h2919;
         16'h9e70, 16'h9e71, 16'h9e72, 16'h9e73, 16'h9e74, 16'h9e75, 16'h9e76, 16'h9e77 	:	val_out <= 16'h2906;
         16'h9e78, 16'h9e79, 16'h9e7a, 16'h9e7b, 16'h9e7c, 16'h9e7d, 16'h9e7e, 16'h9e7f 	:	val_out <= 16'h28f4;
         16'h9e80, 16'h9e81, 16'h9e82, 16'h9e83, 16'h9e84, 16'h9e85, 16'h9e86, 16'h9e87 	:	val_out <= 16'h28e2;
         16'h9e88, 16'h9e89, 16'h9e8a, 16'h9e8b, 16'h9e8c, 16'h9e8d, 16'h9e8e, 16'h9e8f 	:	val_out <= 16'h28cf;
         16'h9e90, 16'h9e91, 16'h9e92, 16'h9e93, 16'h9e94, 16'h9e95, 16'h9e96, 16'h9e97 	:	val_out <= 16'h28bd;
         16'h9e98, 16'h9e99, 16'h9e9a, 16'h9e9b, 16'h9e9c, 16'h9e9d, 16'h9e9e, 16'h9e9f 	:	val_out <= 16'h28aa;
         16'h9ea0, 16'h9ea1, 16'h9ea2, 16'h9ea3, 16'h9ea4, 16'h9ea5, 16'h9ea6, 16'h9ea7 	:	val_out <= 16'h2898;
         16'h9ea8, 16'h9ea9, 16'h9eaa, 16'h9eab, 16'h9eac, 16'h9ead, 16'h9eae, 16'h9eaf 	:	val_out <= 16'h2886;
         16'h9eb0, 16'h9eb1, 16'h9eb2, 16'h9eb3, 16'h9eb4, 16'h9eb5, 16'h9eb6, 16'h9eb7 	:	val_out <= 16'h2873;
         16'h9eb8, 16'h9eb9, 16'h9eba, 16'h9ebb, 16'h9ebc, 16'h9ebd, 16'h9ebe, 16'h9ebf 	:	val_out <= 16'h2861;
         16'h9ec0, 16'h9ec1, 16'h9ec2, 16'h9ec3, 16'h9ec4, 16'h9ec5, 16'h9ec6, 16'h9ec7 	:	val_out <= 16'h284f;
         16'h9ec8, 16'h9ec9, 16'h9eca, 16'h9ecb, 16'h9ecc, 16'h9ecd, 16'h9ece, 16'h9ecf 	:	val_out <= 16'h283c;
         16'h9ed0, 16'h9ed1, 16'h9ed2, 16'h9ed3, 16'h9ed4, 16'h9ed5, 16'h9ed6, 16'h9ed7 	:	val_out <= 16'h282a;
         16'h9ed8, 16'h9ed9, 16'h9eda, 16'h9edb, 16'h9edc, 16'h9edd, 16'h9ede, 16'h9edf 	:	val_out <= 16'h2818;
         16'h9ee0, 16'h9ee1, 16'h9ee2, 16'h9ee3, 16'h9ee4, 16'h9ee5, 16'h9ee6, 16'h9ee7 	:	val_out <= 16'h2806;
         16'h9ee8, 16'h9ee9, 16'h9eea, 16'h9eeb, 16'h9eec, 16'h9eed, 16'h9eee, 16'h9eef 	:	val_out <= 16'h27f3;
         16'h9ef0, 16'h9ef1, 16'h9ef2, 16'h9ef3, 16'h9ef4, 16'h9ef5, 16'h9ef6, 16'h9ef7 	:	val_out <= 16'h27e1;
         16'h9ef8, 16'h9ef9, 16'h9efa, 16'h9efb, 16'h9efc, 16'h9efd, 16'h9efe, 16'h9eff 	:	val_out <= 16'h27cf;
         16'h9f00, 16'h9f01, 16'h9f02, 16'h9f03, 16'h9f04, 16'h9f05, 16'h9f06, 16'h9f07 	:	val_out <= 16'h27bd;
         16'h9f08, 16'h9f09, 16'h9f0a, 16'h9f0b, 16'h9f0c, 16'h9f0d, 16'h9f0e, 16'h9f0f 	:	val_out <= 16'h27aa;
         16'h9f10, 16'h9f11, 16'h9f12, 16'h9f13, 16'h9f14, 16'h9f15, 16'h9f16, 16'h9f17 	:	val_out <= 16'h2798;
         16'h9f18, 16'h9f19, 16'h9f1a, 16'h9f1b, 16'h9f1c, 16'h9f1d, 16'h9f1e, 16'h9f1f 	:	val_out <= 16'h2786;
         16'h9f20, 16'h9f21, 16'h9f22, 16'h9f23, 16'h9f24, 16'h9f25, 16'h9f26, 16'h9f27 	:	val_out <= 16'h2774;
         16'h9f28, 16'h9f29, 16'h9f2a, 16'h9f2b, 16'h9f2c, 16'h9f2d, 16'h9f2e, 16'h9f2f 	:	val_out <= 16'h2762;
         16'h9f30, 16'h9f31, 16'h9f32, 16'h9f33, 16'h9f34, 16'h9f35, 16'h9f36, 16'h9f37 	:	val_out <= 16'h2750;
         16'h9f38, 16'h9f39, 16'h9f3a, 16'h9f3b, 16'h9f3c, 16'h9f3d, 16'h9f3e, 16'h9f3f 	:	val_out <= 16'h273e;
         16'h9f40, 16'h9f41, 16'h9f42, 16'h9f43, 16'h9f44, 16'h9f45, 16'h9f46, 16'h9f47 	:	val_out <= 16'h272b;
         16'h9f48, 16'h9f49, 16'h9f4a, 16'h9f4b, 16'h9f4c, 16'h9f4d, 16'h9f4e, 16'h9f4f 	:	val_out <= 16'h2719;
         16'h9f50, 16'h9f51, 16'h9f52, 16'h9f53, 16'h9f54, 16'h9f55, 16'h9f56, 16'h9f57 	:	val_out <= 16'h2707;
         16'h9f58, 16'h9f59, 16'h9f5a, 16'h9f5b, 16'h9f5c, 16'h9f5d, 16'h9f5e, 16'h9f5f 	:	val_out <= 16'h26f5;
         16'h9f60, 16'h9f61, 16'h9f62, 16'h9f63, 16'h9f64, 16'h9f65, 16'h9f66, 16'h9f67 	:	val_out <= 16'h26e3;
         16'h9f68, 16'h9f69, 16'h9f6a, 16'h9f6b, 16'h9f6c, 16'h9f6d, 16'h9f6e, 16'h9f6f 	:	val_out <= 16'h26d1;
         16'h9f70, 16'h9f71, 16'h9f72, 16'h9f73, 16'h9f74, 16'h9f75, 16'h9f76, 16'h9f77 	:	val_out <= 16'h26bf;
         16'h9f78, 16'h9f79, 16'h9f7a, 16'h9f7b, 16'h9f7c, 16'h9f7d, 16'h9f7e, 16'h9f7f 	:	val_out <= 16'h26ad;
         16'h9f80, 16'h9f81, 16'h9f82, 16'h9f83, 16'h9f84, 16'h9f85, 16'h9f86, 16'h9f87 	:	val_out <= 16'h269b;
         16'h9f88, 16'h9f89, 16'h9f8a, 16'h9f8b, 16'h9f8c, 16'h9f8d, 16'h9f8e, 16'h9f8f 	:	val_out <= 16'h2689;
         16'h9f90, 16'h9f91, 16'h9f92, 16'h9f93, 16'h9f94, 16'h9f95, 16'h9f96, 16'h9f97 	:	val_out <= 16'h2677;
         16'h9f98, 16'h9f99, 16'h9f9a, 16'h9f9b, 16'h9f9c, 16'h9f9d, 16'h9f9e, 16'h9f9f 	:	val_out <= 16'h2665;
         16'h9fa0, 16'h9fa1, 16'h9fa2, 16'h9fa3, 16'h9fa4, 16'h9fa5, 16'h9fa6, 16'h9fa7 	:	val_out <= 16'h2653;
         16'h9fa8, 16'h9fa9, 16'h9faa, 16'h9fab, 16'h9fac, 16'h9fad, 16'h9fae, 16'h9faf 	:	val_out <= 16'h2641;
         16'h9fb0, 16'h9fb1, 16'h9fb2, 16'h9fb3, 16'h9fb4, 16'h9fb5, 16'h9fb6, 16'h9fb7 	:	val_out <= 16'h262f;
         16'h9fb8, 16'h9fb9, 16'h9fba, 16'h9fbb, 16'h9fbc, 16'h9fbd, 16'h9fbe, 16'h9fbf 	:	val_out <= 16'h261e;
         16'h9fc0, 16'h9fc1, 16'h9fc2, 16'h9fc3, 16'h9fc4, 16'h9fc5, 16'h9fc6, 16'h9fc7 	:	val_out <= 16'h260c;
         16'h9fc8, 16'h9fc9, 16'h9fca, 16'h9fcb, 16'h9fcc, 16'h9fcd, 16'h9fce, 16'h9fcf 	:	val_out <= 16'h25fa;
         16'h9fd0, 16'h9fd1, 16'h9fd2, 16'h9fd3, 16'h9fd4, 16'h9fd5, 16'h9fd6, 16'h9fd7 	:	val_out <= 16'h25e8;
         16'h9fd8, 16'h9fd9, 16'h9fda, 16'h9fdb, 16'h9fdc, 16'h9fdd, 16'h9fde, 16'h9fdf 	:	val_out <= 16'h25d6;
         16'h9fe0, 16'h9fe1, 16'h9fe2, 16'h9fe3, 16'h9fe4, 16'h9fe5, 16'h9fe6, 16'h9fe7 	:	val_out <= 16'h25c4;
         16'h9fe8, 16'h9fe9, 16'h9fea, 16'h9feb, 16'h9fec, 16'h9fed, 16'h9fee, 16'h9fef 	:	val_out <= 16'h25b2;
         16'h9ff0, 16'h9ff1, 16'h9ff2, 16'h9ff3, 16'h9ff4, 16'h9ff5, 16'h9ff6, 16'h9ff7 	:	val_out <= 16'h25a1;
         16'h9ff8, 16'h9ff9, 16'h9ffa, 16'h9ffb, 16'h9ffc, 16'h9ffd, 16'h9ffe, 16'h9fff 	:	val_out <= 16'h258f;
         16'ha000, 16'ha001, 16'ha002, 16'ha003, 16'ha004, 16'ha005, 16'ha006, 16'ha007 	:	val_out <= 16'h257d;
         16'ha008, 16'ha009, 16'ha00a, 16'ha00b, 16'ha00c, 16'ha00d, 16'ha00e, 16'ha00f 	:	val_out <= 16'h256b;
         16'ha010, 16'ha011, 16'ha012, 16'ha013, 16'ha014, 16'ha015, 16'ha016, 16'ha017 	:	val_out <= 16'h255a;
         16'ha018, 16'ha019, 16'ha01a, 16'ha01b, 16'ha01c, 16'ha01d, 16'ha01e, 16'ha01f 	:	val_out <= 16'h2548;
         16'ha020, 16'ha021, 16'ha022, 16'ha023, 16'ha024, 16'ha025, 16'ha026, 16'ha027 	:	val_out <= 16'h2536;
         16'ha028, 16'ha029, 16'ha02a, 16'ha02b, 16'ha02c, 16'ha02d, 16'ha02e, 16'ha02f 	:	val_out <= 16'h2524;
         16'ha030, 16'ha031, 16'ha032, 16'ha033, 16'ha034, 16'ha035, 16'ha036, 16'ha037 	:	val_out <= 16'h2513;
         16'ha038, 16'ha039, 16'ha03a, 16'ha03b, 16'ha03c, 16'ha03d, 16'ha03e, 16'ha03f 	:	val_out <= 16'h2501;
         16'ha040, 16'ha041, 16'ha042, 16'ha043, 16'ha044, 16'ha045, 16'ha046, 16'ha047 	:	val_out <= 16'h24ef;
         16'ha048, 16'ha049, 16'ha04a, 16'ha04b, 16'ha04c, 16'ha04d, 16'ha04e, 16'ha04f 	:	val_out <= 16'h24de;
         16'ha050, 16'ha051, 16'ha052, 16'ha053, 16'ha054, 16'ha055, 16'ha056, 16'ha057 	:	val_out <= 16'h24cc;
         16'ha058, 16'ha059, 16'ha05a, 16'ha05b, 16'ha05c, 16'ha05d, 16'ha05e, 16'ha05f 	:	val_out <= 16'h24ba;
         16'ha060, 16'ha061, 16'ha062, 16'ha063, 16'ha064, 16'ha065, 16'ha066, 16'ha067 	:	val_out <= 16'h24a9;
         16'ha068, 16'ha069, 16'ha06a, 16'ha06b, 16'ha06c, 16'ha06d, 16'ha06e, 16'ha06f 	:	val_out <= 16'h2497;
         16'ha070, 16'ha071, 16'ha072, 16'ha073, 16'ha074, 16'ha075, 16'ha076, 16'ha077 	:	val_out <= 16'h2486;
         16'ha078, 16'ha079, 16'ha07a, 16'ha07b, 16'ha07c, 16'ha07d, 16'ha07e, 16'ha07f 	:	val_out <= 16'h2474;
         16'ha080, 16'ha081, 16'ha082, 16'ha083, 16'ha084, 16'ha085, 16'ha086, 16'ha087 	:	val_out <= 16'h2462;
         16'ha088, 16'ha089, 16'ha08a, 16'ha08b, 16'ha08c, 16'ha08d, 16'ha08e, 16'ha08f 	:	val_out <= 16'h2451;
         16'ha090, 16'ha091, 16'ha092, 16'ha093, 16'ha094, 16'ha095, 16'ha096, 16'ha097 	:	val_out <= 16'h243f;
         16'ha098, 16'ha099, 16'ha09a, 16'ha09b, 16'ha09c, 16'ha09d, 16'ha09e, 16'ha09f 	:	val_out <= 16'h242e;
         16'ha0a0, 16'ha0a1, 16'ha0a2, 16'ha0a3, 16'ha0a4, 16'ha0a5, 16'ha0a6, 16'ha0a7 	:	val_out <= 16'h241c;
         16'ha0a8, 16'ha0a9, 16'ha0aa, 16'ha0ab, 16'ha0ac, 16'ha0ad, 16'ha0ae, 16'ha0af 	:	val_out <= 16'h240b;
         16'ha0b0, 16'ha0b1, 16'ha0b2, 16'ha0b3, 16'ha0b4, 16'ha0b5, 16'ha0b6, 16'ha0b7 	:	val_out <= 16'h23f9;
         16'ha0b8, 16'ha0b9, 16'ha0ba, 16'ha0bb, 16'ha0bc, 16'ha0bd, 16'ha0be, 16'ha0bf 	:	val_out <= 16'h23e8;
         16'ha0c0, 16'ha0c1, 16'ha0c2, 16'ha0c3, 16'ha0c4, 16'ha0c5, 16'ha0c6, 16'ha0c7 	:	val_out <= 16'h23d6;
         16'ha0c8, 16'ha0c9, 16'ha0ca, 16'ha0cb, 16'ha0cc, 16'ha0cd, 16'ha0ce, 16'ha0cf 	:	val_out <= 16'h23c5;
         16'ha0d0, 16'ha0d1, 16'ha0d2, 16'ha0d3, 16'ha0d4, 16'ha0d5, 16'ha0d6, 16'ha0d7 	:	val_out <= 16'h23b4;
         16'ha0d8, 16'ha0d9, 16'ha0da, 16'ha0db, 16'ha0dc, 16'ha0dd, 16'ha0de, 16'ha0df 	:	val_out <= 16'h23a2;
         16'ha0e0, 16'ha0e1, 16'ha0e2, 16'ha0e3, 16'ha0e4, 16'ha0e5, 16'ha0e6, 16'ha0e7 	:	val_out <= 16'h2391;
         16'ha0e8, 16'ha0e9, 16'ha0ea, 16'ha0eb, 16'ha0ec, 16'ha0ed, 16'ha0ee, 16'ha0ef 	:	val_out <= 16'h237f;
         16'ha0f0, 16'ha0f1, 16'ha0f2, 16'ha0f3, 16'ha0f4, 16'ha0f5, 16'ha0f6, 16'ha0f7 	:	val_out <= 16'h236e;
         16'ha0f8, 16'ha0f9, 16'ha0fa, 16'ha0fb, 16'ha0fc, 16'ha0fd, 16'ha0fe, 16'ha0ff 	:	val_out <= 16'h235d;
         16'ha100, 16'ha101, 16'ha102, 16'ha103, 16'ha104, 16'ha105, 16'ha106, 16'ha107 	:	val_out <= 16'h234b;
         16'ha108, 16'ha109, 16'ha10a, 16'ha10b, 16'ha10c, 16'ha10d, 16'ha10e, 16'ha10f 	:	val_out <= 16'h233a;
         16'ha110, 16'ha111, 16'ha112, 16'ha113, 16'ha114, 16'ha115, 16'ha116, 16'ha117 	:	val_out <= 16'h2329;
         16'ha118, 16'ha119, 16'ha11a, 16'ha11b, 16'ha11c, 16'ha11d, 16'ha11e, 16'ha11f 	:	val_out <= 16'h2317;
         16'ha120, 16'ha121, 16'ha122, 16'ha123, 16'ha124, 16'ha125, 16'ha126, 16'ha127 	:	val_out <= 16'h2306;
         16'ha128, 16'ha129, 16'ha12a, 16'ha12b, 16'ha12c, 16'ha12d, 16'ha12e, 16'ha12f 	:	val_out <= 16'h22f5;
         16'ha130, 16'ha131, 16'ha132, 16'ha133, 16'ha134, 16'ha135, 16'ha136, 16'ha137 	:	val_out <= 16'h22e4;
         16'ha138, 16'ha139, 16'ha13a, 16'ha13b, 16'ha13c, 16'ha13d, 16'ha13e, 16'ha13f 	:	val_out <= 16'h22d2;
         16'ha140, 16'ha141, 16'ha142, 16'ha143, 16'ha144, 16'ha145, 16'ha146, 16'ha147 	:	val_out <= 16'h22c1;
         16'ha148, 16'ha149, 16'ha14a, 16'ha14b, 16'ha14c, 16'ha14d, 16'ha14e, 16'ha14f 	:	val_out <= 16'h22b0;
         16'ha150, 16'ha151, 16'ha152, 16'ha153, 16'ha154, 16'ha155, 16'ha156, 16'ha157 	:	val_out <= 16'h229f;
         16'ha158, 16'ha159, 16'ha15a, 16'ha15b, 16'ha15c, 16'ha15d, 16'ha15e, 16'ha15f 	:	val_out <= 16'h228e;
         16'ha160, 16'ha161, 16'ha162, 16'ha163, 16'ha164, 16'ha165, 16'ha166, 16'ha167 	:	val_out <= 16'h227c;
         16'ha168, 16'ha169, 16'ha16a, 16'ha16b, 16'ha16c, 16'ha16d, 16'ha16e, 16'ha16f 	:	val_out <= 16'h226b;
         16'ha170, 16'ha171, 16'ha172, 16'ha173, 16'ha174, 16'ha175, 16'ha176, 16'ha177 	:	val_out <= 16'h225a;
         16'ha178, 16'ha179, 16'ha17a, 16'ha17b, 16'ha17c, 16'ha17d, 16'ha17e, 16'ha17f 	:	val_out <= 16'h2249;
         16'ha180, 16'ha181, 16'ha182, 16'ha183, 16'ha184, 16'ha185, 16'ha186, 16'ha187 	:	val_out <= 16'h2238;
         16'ha188, 16'ha189, 16'ha18a, 16'ha18b, 16'ha18c, 16'ha18d, 16'ha18e, 16'ha18f 	:	val_out <= 16'h2227;
         16'ha190, 16'ha191, 16'ha192, 16'ha193, 16'ha194, 16'ha195, 16'ha196, 16'ha197 	:	val_out <= 16'h2216;
         16'ha198, 16'ha199, 16'ha19a, 16'ha19b, 16'ha19c, 16'ha19d, 16'ha19e, 16'ha19f 	:	val_out <= 16'h2205;
         16'ha1a0, 16'ha1a1, 16'ha1a2, 16'ha1a3, 16'ha1a4, 16'ha1a5, 16'ha1a6, 16'ha1a7 	:	val_out <= 16'h21f4;
         16'ha1a8, 16'ha1a9, 16'ha1aa, 16'ha1ab, 16'ha1ac, 16'ha1ad, 16'ha1ae, 16'ha1af 	:	val_out <= 16'h21e3;
         16'ha1b0, 16'ha1b1, 16'ha1b2, 16'ha1b3, 16'ha1b4, 16'ha1b5, 16'ha1b6, 16'ha1b7 	:	val_out <= 16'h21d2;
         16'ha1b8, 16'ha1b9, 16'ha1ba, 16'ha1bb, 16'ha1bc, 16'ha1bd, 16'ha1be, 16'ha1bf 	:	val_out <= 16'h21c0;
         16'ha1c0, 16'ha1c1, 16'ha1c2, 16'ha1c3, 16'ha1c4, 16'ha1c5, 16'ha1c6, 16'ha1c7 	:	val_out <= 16'h21af;
         16'ha1c8, 16'ha1c9, 16'ha1ca, 16'ha1cb, 16'ha1cc, 16'ha1cd, 16'ha1ce, 16'ha1cf 	:	val_out <= 16'h219f;
         16'ha1d0, 16'ha1d1, 16'ha1d2, 16'ha1d3, 16'ha1d4, 16'ha1d5, 16'ha1d6, 16'ha1d7 	:	val_out <= 16'h218e;
         16'ha1d8, 16'ha1d9, 16'ha1da, 16'ha1db, 16'ha1dc, 16'ha1dd, 16'ha1de, 16'ha1df 	:	val_out <= 16'h217d;
         16'ha1e0, 16'ha1e1, 16'ha1e2, 16'ha1e3, 16'ha1e4, 16'ha1e5, 16'ha1e6, 16'ha1e7 	:	val_out <= 16'h216c;
         16'ha1e8, 16'ha1e9, 16'ha1ea, 16'ha1eb, 16'ha1ec, 16'ha1ed, 16'ha1ee, 16'ha1ef 	:	val_out <= 16'h215b;
         16'ha1f0, 16'ha1f1, 16'ha1f2, 16'ha1f3, 16'ha1f4, 16'ha1f5, 16'ha1f6, 16'ha1f7 	:	val_out <= 16'h214a;
         16'ha1f8, 16'ha1f9, 16'ha1fa, 16'ha1fb, 16'ha1fc, 16'ha1fd, 16'ha1fe, 16'ha1ff 	:	val_out <= 16'h2139;
         16'ha200, 16'ha201, 16'ha202, 16'ha203, 16'ha204, 16'ha205, 16'ha206, 16'ha207 	:	val_out <= 16'h2128;
         16'ha208, 16'ha209, 16'ha20a, 16'ha20b, 16'ha20c, 16'ha20d, 16'ha20e, 16'ha20f 	:	val_out <= 16'h2117;
         16'ha210, 16'ha211, 16'ha212, 16'ha213, 16'ha214, 16'ha215, 16'ha216, 16'ha217 	:	val_out <= 16'h2106;
         16'ha218, 16'ha219, 16'ha21a, 16'ha21b, 16'ha21c, 16'ha21d, 16'ha21e, 16'ha21f 	:	val_out <= 16'h20f5;
         16'ha220, 16'ha221, 16'ha222, 16'ha223, 16'ha224, 16'ha225, 16'ha226, 16'ha227 	:	val_out <= 16'h20e5;
         16'ha228, 16'ha229, 16'ha22a, 16'ha22b, 16'ha22c, 16'ha22d, 16'ha22e, 16'ha22f 	:	val_out <= 16'h20d4;
         16'ha230, 16'ha231, 16'ha232, 16'ha233, 16'ha234, 16'ha235, 16'ha236, 16'ha237 	:	val_out <= 16'h20c3;
         16'ha238, 16'ha239, 16'ha23a, 16'ha23b, 16'ha23c, 16'ha23d, 16'ha23e, 16'ha23f 	:	val_out <= 16'h20b2;
         16'ha240, 16'ha241, 16'ha242, 16'ha243, 16'ha244, 16'ha245, 16'ha246, 16'ha247 	:	val_out <= 16'h20a1;
         16'ha248, 16'ha249, 16'ha24a, 16'ha24b, 16'ha24c, 16'ha24d, 16'ha24e, 16'ha24f 	:	val_out <= 16'h2091;
         16'ha250, 16'ha251, 16'ha252, 16'ha253, 16'ha254, 16'ha255, 16'ha256, 16'ha257 	:	val_out <= 16'h2080;
         16'ha258, 16'ha259, 16'ha25a, 16'ha25b, 16'ha25c, 16'ha25d, 16'ha25e, 16'ha25f 	:	val_out <= 16'h206f;
         16'ha260, 16'ha261, 16'ha262, 16'ha263, 16'ha264, 16'ha265, 16'ha266, 16'ha267 	:	val_out <= 16'h205f;
         16'ha268, 16'ha269, 16'ha26a, 16'ha26b, 16'ha26c, 16'ha26d, 16'ha26e, 16'ha26f 	:	val_out <= 16'h204e;
         16'ha270, 16'ha271, 16'ha272, 16'ha273, 16'ha274, 16'ha275, 16'ha276, 16'ha277 	:	val_out <= 16'h203d;
         16'ha278, 16'ha279, 16'ha27a, 16'ha27b, 16'ha27c, 16'ha27d, 16'ha27e, 16'ha27f 	:	val_out <= 16'h202c;
         16'ha280, 16'ha281, 16'ha282, 16'ha283, 16'ha284, 16'ha285, 16'ha286, 16'ha287 	:	val_out <= 16'h201c;
         16'ha288, 16'ha289, 16'ha28a, 16'ha28b, 16'ha28c, 16'ha28d, 16'ha28e, 16'ha28f 	:	val_out <= 16'h200b;
         16'ha290, 16'ha291, 16'ha292, 16'ha293, 16'ha294, 16'ha295, 16'ha296, 16'ha297 	:	val_out <= 16'h1ffb;
         16'ha298, 16'ha299, 16'ha29a, 16'ha29b, 16'ha29c, 16'ha29d, 16'ha29e, 16'ha29f 	:	val_out <= 16'h1fea;
         16'ha2a0, 16'ha2a1, 16'ha2a2, 16'ha2a3, 16'ha2a4, 16'ha2a5, 16'ha2a6, 16'ha2a7 	:	val_out <= 16'h1fd9;
         16'ha2a8, 16'ha2a9, 16'ha2aa, 16'ha2ab, 16'ha2ac, 16'ha2ad, 16'ha2ae, 16'ha2af 	:	val_out <= 16'h1fc9;
         16'ha2b0, 16'ha2b1, 16'ha2b2, 16'ha2b3, 16'ha2b4, 16'ha2b5, 16'ha2b6, 16'ha2b7 	:	val_out <= 16'h1fb8;
         16'ha2b8, 16'ha2b9, 16'ha2ba, 16'ha2bb, 16'ha2bc, 16'ha2bd, 16'ha2be, 16'ha2bf 	:	val_out <= 16'h1fa8;
         16'ha2c0, 16'ha2c1, 16'ha2c2, 16'ha2c3, 16'ha2c4, 16'ha2c5, 16'ha2c6, 16'ha2c7 	:	val_out <= 16'h1f97;
         16'ha2c8, 16'ha2c9, 16'ha2ca, 16'ha2cb, 16'ha2cc, 16'ha2cd, 16'ha2ce, 16'ha2cf 	:	val_out <= 16'h1f87;
         16'ha2d0, 16'ha2d1, 16'ha2d2, 16'ha2d3, 16'ha2d4, 16'ha2d5, 16'ha2d6, 16'ha2d7 	:	val_out <= 16'h1f76;
         16'ha2d8, 16'ha2d9, 16'ha2da, 16'ha2db, 16'ha2dc, 16'ha2dd, 16'ha2de, 16'ha2df 	:	val_out <= 16'h1f66;
         16'ha2e0, 16'ha2e1, 16'ha2e2, 16'ha2e3, 16'ha2e4, 16'ha2e5, 16'ha2e6, 16'ha2e7 	:	val_out <= 16'h1f55;
         16'ha2e8, 16'ha2e9, 16'ha2ea, 16'ha2eb, 16'ha2ec, 16'ha2ed, 16'ha2ee, 16'ha2ef 	:	val_out <= 16'h1f45;
         16'ha2f0, 16'ha2f1, 16'ha2f2, 16'ha2f3, 16'ha2f4, 16'ha2f5, 16'ha2f6, 16'ha2f7 	:	val_out <= 16'h1f34;
         16'ha2f8, 16'ha2f9, 16'ha2fa, 16'ha2fb, 16'ha2fc, 16'ha2fd, 16'ha2fe, 16'ha2ff 	:	val_out <= 16'h1f24;
         16'ha300, 16'ha301, 16'ha302, 16'ha303, 16'ha304, 16'ha305, 16'ha306, 16'ha307 	:	val_out <= 16'h1f13;
         16'ha308, 16'ha309, 16'ha30a, 16'ha30b, 16'ha30c, 16'ha30d, 16'ha30e, 16'ha30f 	:	val_out <= 16'h1f03;
         16'ha310, 16'ha311, 16'ha312, 16'ha313, 16'ha314, 16'ha315, 16'ha316, 16'ha317 	:	val_out <= 16'h1ef2;
         16'ha318, 16'ha319, 16'ha31a, 16'ha31b, 16'ha31c, 16'ha31d, 16'ha31e, 16'ha31f 	:	val_out <= 16'h1ee2;
         16'ha320, 16'ha321, 16'ha322, 16'ha323, 16'ha324, 16'ha325, 16'ha326, 16'ha327 	:	val_out <= 16'h1ed2;
         16'ha328, 16'ha329, 16'ha32a, 16'ha32b, 16'ha32c, 16'ha32d, 16'ha32e, 16'ha32f 	:	val_out <= 16'h1ec1;
         16'ha330, 16'ha331, 16'ha332, 16'ha333, 16'ha334, 16'ha335, 16'ha336, 16'ha337 	:	val_out <= 16'h1eb1;
         16'ha338, 16'ha339, 16'ha33a, 16'ha33b, 16'ha33c, 16'ha33d, 16'ha33e, 16'ha33f 	:	val_out <= 16'h1ea1;
         16'ha340, 16'ha341, 16'ha342, 16'ha343, 16'ha344, 16'ha345, 16'ha346, 16'ha347 	:	val_out <= 16'h1e90;
         16'ha348, 16'ha349, 16'ha34a, 16'ha34b, 16'ha34c, 16'ha34d, 16'ha34e, 16'ha34f 	:	val_out <= 16'h1e80;
         16'ha350, 16'ha351, 16'ha352, 16'ha353, 16'ha354, 16'ha355, 16'ha356, 16'ha357 	:	val_out <= 16'h1e70;
         16'ha358, 16'ha359, 16'ha35a, 16'ha35b, 16'ha35c, 16'ha35d, 16'ha35e, 16'ha35f 	:	val_out <= 16'h1e60;
         16'ha360, 16'ha361, 16'ha362, 16'ha363, 16'ha364, 16'ha365, 16'ha366, 16'ha367 	:	val_out <= 16'h1e4f;
         16'ha368, 16'ha369, 16'ha36a, 16'ha36b, 16'ha36c, 16'ha36d, 16'ha36e, 16'ha36f 	:	val_out <= 16'h1e3f;
         16'ha370, 16'ha371, 16'ha372, 16'ha373, 16'ha374, 16'ha375, 16'ha376, 16'ha377 	:	val_out <= 16'h1e2f;
         16'ha378, 16'ha379, 16'ha37a, 16'ha37b, 16'ha37c, 16'ha37d, 16'ha37e, 16'ha37f 	:	val_out <= 16'h1e1f;
         16'ha380, 16'ha381, 16'ha382, 16'ha383, 16'ha384, 16'ha385, 16'ha386, 16'ha387 	:	val_out <= 16'h1e0e;
         16'ha388, 16'ha389, 16'ha38a, 16'ha38b, 16'ha38c, 16'ha38d, 16'ha38e, 16'ha38f 	:	val_out <= 16'h1dfe;
         16'ha390, 16'ha391, 16'ha392, 16'ha393, 16'ha394, 16'ha395, 16'ha396, 16'ha397 	:	val_out <= 16'h1dee;
         16'ha398, 16'ha399, 16'ha39a, 16'ha39b, 16'ha39c, 16'ha39d, 16'ha39e, 16'ha39f 	:	val_out <= 16'h1dde;
         16'ha3a0, 16'ha3a1, 16'ha3a2, 16'ha3a3, 16'ha3a4, 16'ha3a5, 16'ha3a6, 16'ha3a7 	:	val_out <= 16'h1dce;
         16'ha3a8, 16'ha3a9, 16'ha3aa, 16'ha3ab, 16'ha3ac, 16'ha3ad, 16'ha3ae, 16'ha3af 	:	val_out <= 16'h1dbe;
         16'ha3b0, 16'ha3b1, 16'ha3b2, 16'ha3b3, 16'ha3b4, 16'ha3b5, 16'ha3b6, 16'ha3b7 	:	val_out <= 16'h1dae;
         16'ha3b8, 16'ha3b9, 16'ha3ba, 16'ha3bb, 16'ha3bc, 16'ha3bd, 16'ha3be, 16'ha3bf 	:	val_out <= 16'h1d9e;
         16'ha3c0, 16'ha3c1, 16'ha3c2, 16'ha3c3, 16'ha3c4, 16'ha3c5, 16'ha3c6, 16'ha3c7 	:	val_out <= 16'h1d8e;
         16'ha3c8, 16'ha3c9, 16'ha3ca, 16'ha3cb, 16'ha3cc, 16'ha3cd, 16'ha3ce, 16'ha3cf 	:	val_out <= 16'h1d7d;
         16'ha3d0, 16'ha3d1, 16'ha3d2, 16'ha3d3, 16'ha3d4, 16'ha3d5, 16'ha3d6, 16'ha3d7 	:	val_out <= 16'h1d6d;
         16'ha3d8, 16'ha3d9, 16'ha3da, 16'ha3db, 16'ha3dc, 16'ha3dd, 16'ha3de, 16'ha3df 	:	val_out <= 16'h1d5d;
         16'ha3e0, 16'ha3e1, 16'ha3e2, 16'ha3e3, 16'ha3e4, 16'ha3e5, 16'ha3e6, 16'ha3e7 	:	val_out <= 16'h1d4d;
         16'ha3e8, 16'ha3e9, 16'ha3ea, 16'ha3eb, 16'ha3ec, 16'ha3ed, 16'ha3ee, 16'ha3ef 	:	val_out <= 16'h1d3d;
         16'ha3f0, 16'ha3f1, 16'ha3f2, 16'ha3f3, 16'ha3f4, 16'ha3f5, 16'ha3f6, 16'ha3f7 	:	val_out <= 16'h1d2d;
         16'ha3f8, 16'ha3f9, 16'ha3fa, 16'ha3fb, 16'ha3fc, 16'ha3fd, 16'ha3fe, 16'ha3ff 	:	val_out <= 16'h1d1d;
         16'ha400, 16'ha401, 16'ha402, 16'ha403, 16'ha404, 16'ha405, 16'ha406, 16'ha407 	:	val_out <= 16'h1d0d;
         16'ha408, 16'ha409, 16'ha40a, 16'ha40b, 16'ha40c, 16'ha40d, 16'ha40e, 16'ha40f 	:	val_out <= 16'h1cfe;
         16'ha410, 16'ha411, 16'ha412, 16'ha413, 16'ha414, 16'ha415, 16'ha416, 16'ha417 	:	val_out <= 16'h1cee;
         16'ha418, 16'ha419, 16'ha41a, 16'ha41b, 16'ha41c, 16'ha41d, 16'ha41e, 16'ha41f 	:	val_out <= 16'h1cde;
         16'ha420, 16'ha421, 16'ha422, 16'ha423, 16'ha424, 16'ha425, 16'ha426, 16'ha427 	:	val_out <= 16'h1cce;
         16'ha428, 16'ha429, 16'ha42a, 16'ha42b, 16'ha42c, 16'ha42d, 16'ha42e, 16'ha42f 	:	val_out <= 16'h1cbe;
         16'ha430, 16'ha431, 16'ha432, 16'ha433, 16'ha434, 16'ha435, 16'ha436, 16'ha437 	:	val_out <= 16'h1cae;
         16'ha438, 16'ha439, 16'ha43a, 16'ha43b, 16'ha43c, 16'ha43d, 16'ha43e, 16'ha43f 	:	val_out <= 16'h1c9e;
         16'ha440, 16'ha441, 16'ha442, 16'ha443, 16'ha444, 16'ha445, 16'ha446, 16'ha447 	:	val_out <= 16'h1c8e;
         16'ha448, 16'ha449, 16'ha44a, 16'ha44b, 16'ha44c, 16'ha44d, 16'ha44e, 16'ha44f 	:	val_out <= 16'h1c7f;
         16'ha450, 16'ha451, 16'ha452, 16'ha453, 16'ha454, 16'ha455, 16'ha456, 16'ha457 	:	val_out <= 16'h1c6f;
         16'ha458, 16'ha459, 16'ha45a, 16'ha45b, 16'ha45c, 16'ha45d, 16'ha45e, 16'ha45f 	:	val_out <= 16'h1c5f;
         16'ha460, 16'ha461, 16'ha462, 16'ha463, 16'ha464, 16'ha465, 16'ha466, 16'ha467 	:	val_out <= 16'h1c4f;
         16'ha468, 16'ha469, 16'ha46a, 16'ha46b, 16'ha46c, 16'ha46d, 16'ha46e, 16'ha46f 	:	val_out <= 16'h1c3f;
         16'ha470, 16'ha471, 16'ha472, 16'ha473, 16'ha474, 16'ha475, 16'ha476, 16'ha477 	:	val_out <= 16'h1c30;
         16'ha478, 16'ha479, 16'ha47a, 16'ha47b, 16'ha47c, 16'ha47d, 16'ha47e, 16'ha47f 	:	val_out <= 16'h1c20;
         16'ha480, 16'ha481, 16'ha482, 16'ha483, 16'ha484, 16'ha485, 16'ha486, 16'ha487 	:	val_out <= 16'h1c10;
         16'ha488, 16'ha489, 16'ha48a, 16'ha48b, 16'ha48c, 16'ha48d, 16'ha48e, 16'ha48f 	:	val_out <= 16'h1c01;
         16'ha490, 16'ha491, 16'ha492, 16'ha493, 16'ha494, 16'ha495, 16'ha496, 16'ha497 	:	val_out <= 16'h1bf1;
         16'ha498, 16'ha499, 16'ha49a, 16'ha49b, 16'ha49c, 16'ha49d, 16'ha49e, 16'ha49f 	:	val_out <= 16'h1be1;
         16'ha4a0, 16'ha4a1, 16'ha4a2, 16'ha4a3, 16'ha4a4, 16'ha4a5, 16'ha4a6, 16'ha4a7 	:	val_out <= 16'h1bd2;
         16'ha4a8, 16'ha4a9, 16'ha4aa, 16'ha4ab, 16'ha4ac, 16'ha4ad, 16'ha4ae, 16'ha4af 	:	val_out <= 16'h1bc2;
         16'ha4b0, 16'ha4b1, 16'ha4b2, 16'ha4b3, 16'ha4b4, 16'ha4b5, 16'ha4b6, 16'ha4b7 	:	val_out <= 16'h1bb2;
         16'ha4b8, 16'ha4b9, 16'ha4ba, 16'ha4bb, 16'ha4bc, 16'ha4bd, 16'ha4be, 16'ha4bf 	:	val_out <= 16'h1ba3;
         16'ha4c0, 16'ha4c1, 16'ha4c2, 16'ha4c3, 16'ha4c4, 16'ha4c5, 16'ha4c6, 16'ha4c7 	:	val_out <= 16'h1b93;
         16'ha4c8, 16'ha4c9, 16'ha4ca, 16'ha4cb, 16'ha4cc, 16'ha4cd, 16'ha4ce, 16'ha4cf 	:	val_out <= 16'h1b84;
         16'ha4d0, 16'ha4d1, 16'ha4d2, 16'ha4d3, 16'ha4d4, 16'ha4d5, 16'ha4d6, 16'ha4d7 	:	val_out <= 16'h1b74;
         16'ha4d8, 16'ha4d9, 16'ha4da, 16'ha4db, 16'ha4dc, 16'ha4dd, 16'ha4de, 16'ha4df 	:	val_out <= 16'h1b64;
         16'ha4e0, 16'ha4e1, 16'ha4e2, 16'ha4e3, 16'ha4e4, 16'ha4e5, 16'ha4e6, 16'ha4e7 	:	val_out <= 16'h1b55;
         16'ha4e8, 16'ha4e9, 16'ha4ea, 16'ha4eb, 16'ha4ec, 16'ha4ed, 16'ha4ee, 16'ha4ef 	:	val_out <= 16'h1b45;
         16'ha4f0, 16'ha4f1, 16'ha4f2, 16'ha4f3, 16'ha4f4, 16'ha4f5, 16'ha4f6, 16'ha4f7 	:	val_out <= 16'h1b36;
         16'ha4f8, 16'ha4f9, 16'ha4fa, 16'ha4fb, 16'ha4fc, 16'ha4fd, 16'ha4fe, 16'ha4ff 	:	val_out <= 16'h1b26;
         16'ha500, 16'ha501, 16'ha502, 16'ha503, 16'ha504, 16'ha505, 16'ha506, 16'ha507 	:	val_out <= 16'h1b17;
         16'ha508, 16'ha509, 16'ha50a, 16'ha50b, 16'ha50c, 16'ha50d, 16'ha50e, 16'ha50f 	:	val_out <= 16'h1b08;
         16'ha510, 16'ha511, 16'ha512, 16'ha513, 16'ha514, 16'ha515, 16'ha516, 16'ha517 	:	val_out <= 16'h1af8;
         16'ha518, 16'ha519, 16'ha51a, 16'ha51b, 16'ha51c, 16'ha51d, 16'ha51e, 16'ha51f 	:	val_out <= 16'h1ae9;
         16'ha520, 16'ha521, 16'ha522, 16'ha523, 16'ha524, 16'ha525, 16'ha526, 16'ha527 	:	val_out <= 16'h1ad9;
         16'ha528, 16'ha529, 16'ha52a, 16'ha52b, 16'ha52c, 16'ha52d, 16'ha52e, 16'ha52f 	:	val_out <= 16'h1aca;
         16'ha530, 16'ha531, 16'ha532, 16'ha533, 16'ha534, 16'ha535, 16'ha536, 16'ha537 	:	val_out <= 16'h1aba;
         16'ha538, 16'ha539, 16'ha53a, 16'ha53b, 16'ha53c, 16'ha53d, 16'ha53e, 16'ha53f 	:	val_out <= 16'h1aab;
         16'ha540, 16'ha541, 16'ha542, 16'ha543, 16'ha544, 16'ha545, 16'ha546, 16'ha547 	:	val_out <= 16'h1a9c;
         16'ha548, 16'ha549, 16'ha54a, 16'ha54b, 16'ha54c, 16'ha54d, 16'ha54e, 16'ha54f 	:	val_out <= 16'h1a8c;
         16'ha550, 16'ha551, 16'ha552, 16'ha553, 16'ha554, 16'ha555, 16'ha556, 16'ha557 	:	val_out <= 16'h1a7d;
         16'ha558, 16'ha559, 16'ha55a, 16'ha55b, 16'ha55c, 16'ha55d, 16'ha55e, 16'ha55f 	:	val_out <= 16'h1a6e;
         16'ha560, 16'ha561, 16'ha562, 16'ha563, 16'ha564, 16'ha565, 16'ha566, 16'ha567 	:	val_out <= 16'h1a5f;
         16'ha568, 16'ha569, 16'ha56a, 16'ha56b, 16'ha56c, 16'ha56d, 16'ha56e, 16'ha56f 	:	val_out <= 16'h1a4f;
         16'ha570, 16'ha571, 16'ha572, 16'ha573, 16'ha574, 16'ha575, 16'ha576, 16'ha577 	:	val_out <= 16'h1a40;
         16'ha578, 16'ha579, 16'ha57a, 16'ha57b, 16'ha57c, 16'ha57d, 16'ha57e, 16'ha57f 	:	val_out <= 16'h1a31;
         16'ha580, 16'ha581, 16'ha582, 16'ha583, 16'ha584, 16'ha585, 16'ha586, 16'ha587 	:	val_out <= 16'h1a22;
         16'ha588, 16'ha589, 16'ha58a, 16'ha58b, 16'ha58c, 16'ha58d, 16'ha58e, 16'ha58f 	:	val_out <= 16'h1a12;
         16'ha590, 16'ha591, 16'ha592, 16'ha593, 16'ha594, 16'ha595, 16'ha596, 16'ha597 	:	val_out <= 16'h1a03;
         16'ha598, 16'ha599, 16'ha59a, 16'ha59b, 16'ha59c, 16'ha59d, 16'ha59e, 16'ha59f 	:	val_out <= 16'h19f4;
         16'ha5a0, 16'ha5a1, 16'ha5a2, 16'ha5a3, 16'ha5a4, 16'ha5a5, 16'ha5a6, 16'ha5a7 	:	val_out <= 16'h19e5;
         16'ha5a8, 16'ha5a9, 16'ha5aa, 16'ha5ab, 16'ha5ac, 16'ha5ad, 16'ha5ae, 16'ha5af 	:	val_out <= 16'h19d6;
         16'ha5b0, 16'ha5b1, 16'ha5b2, 16'ha5b3, 16'ha5b4, 16'ha5b5, 16'ha5b6, 16'ha5b7 	:	val_out <= 16'h19c6;
         16'ha5b8, 16'ha5b9, 16'ha5ba, 16'ha5bb, 16'ha5bc, 16'ha5bd, 16'ha5be, 16'ha5bf 	:	val_out <= 16'h19b7;
         16'ha5c0, 16'ha5c1, 16'ha5c2, 16'ha5c3, 16'ha5c4, 16'ha5c5, 16'ha5c6, 16'ha5c7 	:	val_out <= 16'h19a8;
         16'ha5c8, 16'ha5c9, 16'ha5ca, 16'ha5cb, 16'ha5cc, 16'ha5cd, 16'ha5ce, 16'ha5cf 	:	val_out <= 16'h1999;
         16'ha5d0, 16'ha5d1, 16'ha5d2, 16'ha5d3, 16'ha5d4, 16'ha5d5, 16'ha5d6, 16'ha5d7 	:	val_out <= 16'h198a;
         16'ha5d8, 16'ha5d9, 16'ha5da, 16'ha5db, 16'ha5dc, 16'ha5dd, 16'ha5de, 16'ha5df 	:	val_out <= 16'h197b;
         16'ha5e0, 16'ha5e1, 16'ha5e2, 16'ha5e3, 16'ha5e4, 16'ha5e5, 16'ha5e6, 16'ha5e7 	:	val_out <= 16'h196c;
         16'ha5e8, 16'ha5e9, 16'ha5ea, 16'ha5eb, 16'ha5ec, 16'ha5ed, 16'ha5ee, 16'ha5ef 	:	val_out <= 16'h195d;
         16'ha5f0, 16'ha5f1, 16'ha5f2, 16'ha5f3, 16'ha5f4, 16'ha5f5, 16'ha5f6, 16'ha5f7 	:	val_out <= 16'h194e;
         16'ha5f8, 16'ha5f9, 16'ha5fa, 16'ha5fb, 16'ha5fc, 16'ha5fd, 16'ha5fe, 16'ha5ff 	:	val_out <= 16'h193f;
         16'ha600, 16'ha601, 16'ha602, 16'ha603, 16'ha604, 16'ha605, 16'ha606, 16'ha607 	:	val_out <= 16'h1930;
         16'ha608, 16'ha609, 16'ha60a, 16'ha60b, 16'ha60c, 16'ha60d, 16'ha60e, 16'ha60f 	:	val_out <= 16'h1921;
         16'ha610, 16'ha611, 16'ha612, 16'ha613, 16'ha614, 16'ha615, 16'ha616, 16'ha617 	:	val_out <= 16'h1912;
         16'ha618, 16'ha619, 16'ha61a, 16'ha61b, 16'ha61c, 16'ha61d, 16'ha61e, 16'ha61f 	:	val_out <= 16'h1903;
         16'ha620, 16'ha621, 16'ha622, 16'ha623, 16'ha624, 16'ha625, 16'ha626, 16'ha627 	:	val_out <= 16'h18f4;
         16'ha628, 16'ha629, 16'ha62a, 16'ha62b, 16'ha62c, 16'ha62d, 16'ha62e, 16'ha62f 	:	val_out <= 16'h18e5;
         16'ha630, 16'ha631, 16'ha632, 16'ha633, 16'ha634, 16'ha635, 16'ha636, 16'ha637 	:	val_out <= 16'h18d6;
         16'ha638, 16'ha639, 16'ha63a, 16'ha63b, 16'ha63c, 16'ha63d, 16'ha63e, 16'ha63f 	:	val_out <= 16'h18c8;
         16'ha640, 16'ha641, 16'ha642, 16'ha643, 16'ha644, 16'ha645, 16'ha646, 16'ha647 	:	val_out <= 16'h18b9;
         16'ha648, 16'ha649, 16'ha64a, 16'ha64b, 16'ha64c, 16'ha64d, 16'ha64e, 16'ha64f 	:	val_out <= 16'h18aa;
         16'ha650, 16'ha651, 16'ha652, 16'ha653, 16'ha654, 16'ha655, 16'ha656, 16'ha657 	:	val_out <= 16'h189b;
         16'ha658, 16'ha659, 16'ha65a, 16'ha65b, 16'ha65c, 16'ha65d, 16'ha65e, 16'ha65f 	:	val_out <= 16'h188c;
         16'ha660, 16'ha661, 16'ha662, 16'ha663, 16'ha664, 16'ha665, 16'ha666, 16'ha667 	:	val_out <= 16'h187d;
         16'ha668, 16'ha669, 16'ha66a, 16'ha66b, 16'ha66c, 16'ha66d, 16'ha66e, 16'ha66f 	:	val_out <= 16'h186f;
         16'ha670, 16'ha671, 16'ha672, 16'ha673, 16'ha674, 16'ha675, 16'ha676, 16'ha677 	:	val_out <= 16'h1860;
         16'ha678, 16'ha679, 16'ha67a, 16'ha67b, 16'ha67c, 16'ha67d, 16'ha67e, 16'ha67f 	:	val_out <= 16'h1851;
         16'ha680, 16'ha681, 16'ha682, 16'ha683, 16'ha684, 16'ha685, 16'ha686, 16'ha687 	:	val_out <= 16'h1842;
         16'ha688, 16'ha689, 16'ha68a, 16'ha68b, 16'ha68c, 16'ha68d, 16'ha68e, 16'ha68f 	:	val_out <= 16'h1834;
         16'ha690, 16'ha691, 16'ha692, 16'ha693, 16'ha694, 16'ha695, 16'ha696, 16'ha697 	:	val_out <= 16'h1825;
         16'ha698, 16'ha699, 16'ha69a, 16'ha69b, 16'ha69c, 16'ha69d, 16'ha69e, 16'ha69f 	:	val_out <= 16'h1816;
         16'ha6a0, 16'ha6a1, 16'ha6a2, 16'ha6a3, 16'ha6a4, 16'ha6a5, 16'ha6a6, 16'ha6a7 	:	val_out <= 16'h1808;
         16'ha6a8, 16'ha6a9, 16'ha6aa, 16'ha6ab, 16'ha6ac, 16'ha6ad, 16'ha6ae, 16'ha6af 	:	val_out <= 16'h17f9;
         16'ha6b0, 16'ha6b1, 16'ha6b2, 16'ha6b3, 16'ha6b4, 16'ha6b5, 16'ha6b6, 16'ha6b7 	:	val_out <= 16'h17ea;
         16'ha6b8, 16'ha6b9, 16'ha6ba, 16'ha6bb, 16'ha6bc, 16'ha6bd, 16'ha6be, 16'ha6bf 	:	val_out <= 16'h17dc;
         16'ha6c0, 16'ha6c1, 16'ha6c2, 16'ha6c3, 16'ha6c4, 16'ha6c5, 16'ha6c6, 16'ha6c7 	:	val_out <= 16'h17cd;
         16'ha6c8, 16'ha6c9, 16'ha6ca, 16'ha6cb, 16'ha6cc, 16'ha6cd, 16'ha6ce, 16'ha6cf 	:	val_out <= 16'h17bf;
         16'ha6d0, 16'ha6d1, 16'ha6d2, 16'ha6d3, 16'ha6d4, 16'ha6d5, 16'ha6d6, 16'ha6d7 	:	val_out <= 16'h17b0;
         16'ha6d8, 16'ha6d9, 16'ha6da, 16'ha6db, 16'ha6dc, 16'ha6dd, 16'ha6de, 16'ha6df 	:	val_out <= 16'h17a1;
         16'ha6e0, 16'ha6e1, 16'ha6e2, 16'ha6e3, 16'ha6e4, 16'ha6e5, 16'ha6e6, 16'ha6e7 	:	val_out <= 16'h1793;
         16'ha6e8, 16'ha6e9, 16'ha6ea, 16'ha6eb, 16'ha6ec, 16'ha6ed, 16'ha6ee, 16'ha6ef 	:	val_out <= 16'h1784;
         16'ha6f0, 16'ha6f1, 16'ha6f2, 16'ha6f3, 16'ha6f4, 16'ha6f5, 16'ha6f6, 16'ha6f7 	:	val_out <= 16'h1776;
         16'ha6f8, 16'ha6f9, 16'ha6fa, 16'ha6fb, 16'ha6fc, 16'ha6fd, 16'ha6fe, 16'ha6ff 	:	val_out <= 16'h1767;
         16'ha700, 16'ha701, 16'ha702, 16'ha703, 16'ha704, 16'ha705, 16'ha706, 16'ha707 	:	val_out <= 16'h1759;
         16'ha708, 16'ha709, 16'ha70a, 16'ha70b, 16'ha70c, 16'ha70d, 16'ha70e, 16'ha70f 	:	val_out <= 16'h174a;
         16'ha710, 16'ha711, 16'ha712, 16'ha713, 16'ha714, 16'ha715, 16'ha716, 16'ha717 	:	val_out <= 16'h173c;
         16'ha718, 16'ha719, 16'ha71a, 16'ha71b, 16'ha71c, 16'ha71d, 16'ha71e, 16'ha71f 	:	val_out <= 16'h172e;
         16'ha720, 16'ha721, 16'ha722, 16'ha723, 16'ha724, 16'ha725, 16'ha726, 16'ha727 	:	val_out <= 16'h171f;
         16'ha728, 16'ha729, 16'ha72a, 16'ha72b, 16'ha72c, 16'ha72d, 16'ha72e, 16'ha72f 	:	val_out <= 16'h1711;
         16'ha730, 16'ha731, 16'ha732, 16'ha733, 16'ha734, 16'ha735, 16'ha736, 16'ha737 	:	val_out <= 16'h1702;
         16'ha738, 16'ha739, 16'ha73a, 16'ha73b, 16'ha73c, 16'ha73d, 16'ha73e, 16'ha73f 	:	val_out <= 16'h16f4;
         16'ha740, 16'ha741, 16'ha742, 16'ha743, 16'ha744, 16'ha745, 16'ha746, 16'ha747 	:	val_out <= 16'h16e6;
         16'ha748, 16'ha749, 16'ha74a, 16'ha74b, 16'ha74c, 16'ha74d, 16'ha74e, 16'ha74f 	:	val_out <= 16'h16d7;
         16'ha750, 16'ha751, 16'ha752, 16'ha753, 16'ha754, 16'ha755, 16'ha756, 16'ha757 	:	val_out <= 16'h16c9;
         16'ha758, 16'ha759, 16'ha75a, 16'ha75b, 16'ha75c, 16'ha75d, 16'ha75e, 16'ha75f 	:	val_out <= 16'h16bb;
         16'ha760, 16'ha761, 16'ha762, 16'ha763, 16'ha764, 16'ha765, 16'ha766, 16'ha767 	:	val_out <= 16'h16ac;
         16'ha768, 16'ha769, 16'ha76a, 16'ha76b, 16'ha76c, 16'ha76d, 16'ha76e, 16'ha76f 	:	val_out <= 16'h169e;
         16'ha770, 16'ha771, 16'ha772, 16'ha773, 16'ha774, 16'ha775, 16'ha776, 16'ha777 	:	val_out <= 16'h1690;
         16'ha778, 16'ha779, 16'ha77a, 16'ha77b, 16'ha77c, 16'ha77d, 16'ha77e, 16'ha77f 	:	val_out <= 16'h1682;
         16'ha780, 16'ha781, 16'ha782, 16'ha783, 16'ha784, 16'ha785, 16'ha786, 16'ha787 	:	val_out <= 16'h1673;
         16'ha788, 16'ha789, 16'ha78a, 16'ha78b, 16'ha78c, 16'ha78d, 16'ha78e, 16'ha78f 	:	val_out <= 16'h1665;
         16'ha790, 16'ha791, 16'ha792, 16'ha793, 16'ha794, 16'ha795, 16'ha796, 16'ha797 	:	val_out <= 16'h1657;
         16'ha798, 16'ha799, 16'ha79a, 16'ha79b, 16'ha79c, 16'ha79d, 16'ha79e, 16'ha79f 	:	val_out <= 16'h1649;
         16'ha7a0, 16'ha7a1, 16'ha7a2, 16'ha7a3, 16'ha7a4, 16'ha7a5, 16'ha7a6, 16'ha7a7 	:	val_out <= 16'h163b;
         16'ha7a8, 16'ha7a9, 16'ha7aa, 16'ha7ab, 16'ha7ac, 16'ha7ad, 16'ha7ae, 16'ha7af 	:	val_out <= 16'h162c;
         16'ha7b0, 16'ha7b1, 16'ha7b2, 16'ha7b3, 16'ha7b4, 16'ha7b5, 16'ha7b6, 16'ha7b7 	:	val_out <= 16'h161e;
         16'ha7b8, 16'ha7b9, 16'ha7ba, 16'ha7bb, 16'ha7bc, 16'ha7bd, 16'ha7be, 16'ha7bf 	:	val_out <= 16'h1610;
         16'ha7c0, 16'ha7c1, 16'ha7c2, 16'ha7c3, 16'ha7c4, 16'ha7c5, 16'ha7c6, 16'ha7c7 	:	val_out <= 16'h1602;
         16'ha7c8, 16'ha7c9, 16'ha7ca, 16'ha7cb, 16'ha7cc, 16'ha7cd, 16'ha7ce, 16'ha7cf 	:	val_out <= 16'h15f4;
         16'ha7d0, 16'ha7d1, 16'ha7d2, 16'ha7d3, 16'ha7d4, 16'ha7d5, 16'ha7d6, 16'ha7d7 	:	val_out <= 16'h15e6;
         16'ha7d8, 16'ha7d9, 16'ha7da, 16'ha7db, 16'ha7dc, 16'ha7dd, 16'ha7de, 16'ha7df 	:	val_out <= 16'h15d8;
         16'ha7e0, 16'ha7e1, 16'ha7e2, 16'ha7e3, 16'ha7e4, 16'ha7e5, 16'ha7e6, 16'ha7e7 	:	val_out <= 16'h15ca;
         16'ha7e8, 16'ha7e9, 16'ha7ea, 16'ha7eb, 16'ha7ec, 16'ha7ed, 16'ha7ee, 16'ha7ef 	:	val_out <= 16'h15bc;
         16'ha7f0, 16'ha7f1, 16'ha7f2, 16'ha7f3, 16'ha7f4, 16'ha7f5, 16'ha7f6, 16'ha7f7 	:	val_out <= 16'h15ae;
         16'ha7f8, 16'ha7f9, 16'ha7fa, 16'ha7fb, 16'ha7fc, 16'ha7fd, 16'ha7fe, 16'ha7ff 	:	val_out <= 16'h15a0;
         16'ha800, 16'ha801, 16'ha802, 16'ha803, 16'ha804, 16'ha805, 16'ha806, 16'ha807 	:	val_out <= 16'h1592;
         16'ha808, 16'ha809, 16'ha80a, 16'ha80b, 16'ha80c, 16'ha80d, 16'ha80e, 16'ha80f 	:	val_out <= 16'h1584;
         16'ha810, 16'ha811, 16'ha812, 16'ha813, 16'ha814, 16'ha815, 16'ha816, 16'ha817 	:	val_out <= 16'h1576;
         16'ha818, 16'ha819, 16'ha81a, 16'ha81b, 16'ha81c, 16'ha81d, 16'ha81e, 16'ha81f 	:	val_out <= 16'h1568;
         16'ha820, 16'ha821, 16'ha822, 16'ha823, 16'ha824, 16'ha825, 16'ha826, 16'ha827 	:	val_out <= 16'h155a;
         16'ha828, 16'ha829, 16'ha82a, 16'ha82b, 16'ha82c, 16'ha82d, 16'ha82e, 16'ha82f 	:	val_out <= 16'h154c;
         16'ha830, 16'ha831, 16'ha832, 16'ha833, 16'ha834, 16'ha835, 16'ha836, 16'ha837 	:	val_out <= 16'h153e;
         16'ha838, 16'ha839, 16'ha83a, 16'ha83b, 16'ha83c, 16'ha83d, 16'ha83e, 16'ha83f 	:	val_out <= 16'h1531;
         16'ha840, 16'ha841, 16'ha842, 16'ha843, 16'ha844, 16'ha845, 16'ha846, 16'ha847 	:	val_out <= 16'h1523;
         16'ha848, 16'ha849, 16'ha84a, 16'ha84b, 16'ha84c, 16'ha84d, 16'ha84e, 16'ha84f 	:	val_out <= 16'h1515;
         16'ha850, 16'ha851, 16'ha852, 16'ha853, 16'ha854, 16'ha855, 16'ha856, 16'ha857 	:	val_out <= 16'h1507;
         16'ha858, 16'ha859, 16'ha85a, 16'ha85b, 16'ha85c, 16'ha85d, 16'ha85e, 16'ha85f 	:	val_out <= 16'h14f9;
         16'ha860, 16'ha861, 16'ha862, 16'ha863, 16'ha864, 16'ha865, 16'ha866, 16'ha867 	:	val_out <= 16'h14ec;
         16'ha868, 16'ha869, 16'ha86a, 16'ha86b, 16'ha86c, 16'ha86d, 16'ha86e, 16'ha86f 	:	val_out <= 16'h14de;
         16'ha870, 16'ha871, 16'ha872, 16'ha873, 16'ha874, 16'ha875, 16'ha876, 16'ha877 	:	val_out <= 16'h14d0;
         16'ha878, 16'ha879, 16'ha87a, 16'ha87b, 16'ha87c, 16'ha87d, 16'ha87e, 16'ha87f 	:	val_out <= 16'h14c2;
         16'ha880, 16'ha881, 16'ha882, 16'ha883, 16'ha884, 16'ha885, 16'ha886, 16'ha887 	:	val_out <= 16'h14b5;
         16'ha888, 16'ha889, 16'ha88a, 16'ha88b, 16'ha88c, 16'ha88d, 16'ha88e, 16'ha88f 	:	val_out <= 16'h14a7;
         16'ha890, 16'ha891, 16'ha892, 16'ha893, 16'ha894, 16'ha895, 16'ha896, 16'ha897 	:	val_out <= 16'h1499;
         16'ha898, 16'ha899, 16'ha89a, 16'ha89b, 16'ha89c, 16'ha89d, 16'ha89e, 16'ha89f 	:	val_out <= 16'h148c;
         16'ha8a0, 16'ha8a1, 16'ha8a2, 16'ha8a3, 16'ha8a4, 16'ha8a5, 16'ha8a6, 16'ha8a7 	:	val_out <= 16'h147e;
         16'ha8a8, 16'ha8a9, 16'ha8aa, 16'ha8ab, 16'ha8ac, 16'ha8ad, 16'ha8ae, 16'ha8af 	:	val_out <= 16'h1470;
         16'ha8b0, 16'ha8b1, 16'ha8b2, 16'ha8b3, 16'ha8b4, 16'ha8b5, 16'ha8b6, 16'ha8b7 	:	val_out <= 16'h1463;
         16'ha8b8, 16'ha8b9, 16'ha8ba, 16'ha8bb, 16'ha8bc, 16'ha8bd, 16'ha8be, 16'ha8bf 	:	val_out <= 16'h1455;
         16'ha8c0, 16'ha8c1, 16'ha8c2, 16'ha8c3, 16'ha8c4, 16'ha8c5, 16'ha8c6, 16'ha8c7 	:	val_out <= 16'h1447;
         16'ha8c8, 16'ha8c9, 16'ha8ca, 16'ha8cb, 16'ha8cc, 16'ha8cd, 16'ha8ce, 16'ha8cf 	:	val_out <= 16'h143a;
         16'ha8d0, 16'ha8d1, 16'ha8d2, 16'ha8d3, 16'ha8d4, 16'ha8d5, 16'ha8d6, 16'ha8d7 	:	val_out <= 16'h142c;
         16'ha8d8, 16'ha8d9, 16'ha8da, 16'ha8db, 16'ha8dc, 16'ha8dd, 16'ha8de, 16'ha8df 	:	val_out <= 16'h141f;
         16'ha8e0, 16'ha8e1, 16'ha8e2, 16'ha8e3, 16'ha8e4, 16'ha8e5, 16'ha8e6, 16'ha8e7 	:	val_out <= 16'h1411;
         16'ha8e8, 16'ha8e9, 16'ha8ea, 16'ha8eb, 16'ha8ec, 16'ha8ed, 16'ha8ee, 16'ha8ef 	:	val_out <= 16'h1404;
         16'ha8f0, 16'ha8f1, 16'ha8f2, 16'ha8f3, 16'ha8f4, 16'ha8f5, 16'ha8f6, 16'ha8f7 	:	val_out <= 16'h13f6;
         16'ha8f8, 16'ha8f9, 16'ha8fa, 16'ha8fb, 16'ha8fc, 16'ha8fd, 16'ha8fe, 16'ha8ff 	:	val_out <= 16'h13e9;
         16'ha900, 16'ha901, 16'ha902, 16'ha903, 16'ha904, 16'ha905, 16'ha906, 16'ha907 	:	val_out <= 16'h13db;
         16'ha908, 16'ha909, 16'ha90a, 16'ha90b, 16'ha90c, 16'ha90d, 16'ha90e, 16'ha90f 	:	val_out <= 16'h13ce;
         16'ha910, 16'ha911, 16'ha912, 16'ha913, 16'ha914, 16'ha915, 16'ha916, 16'ha917 	:	val_out <= 16'h13c0;
         16'ha918, 16'ha919, 16'ha91a, 16'ha91b, 16'ha91c, 16'ha91d, 16'ha91e, 16'ha91f 	:	val_out <= 16'h13b3;
         16'ha920, 16'ha921, 16'ha922, 16'ha923, 16'ha924, 16'ha925, 16'ha926, 16'ha927 	:	val_out <= 16'h13a6;
         16'ha928, 16'ha929, 16'ha92a, 16'ha92b, 16'ha92c, 16'ha92d, 16'ha92e, 16'ha92f 	:	val_out <= 16'h1398;
         16'ha930, 16'ha931, 16'ha932, 16'ha933, 16'ha934, 16'ha935, 16'ha936, 16'ha937 	:	val_out <= 16'h138b;
         16'ha938, 16'ha939, 16'ha93a, 16'ha93b, 16'ha93c, 16'ha93d, 16'ha93e, 16'ha93f 	:	val_out <= 16'h137e;
         16'ha940, 16'ha941, 16'ha942, 16'ha943, 16'ha944, 16'ha945, 16'ha946, 16'ha947 	:	val_out <= 16'h1370;
         16'ha948, 16'ha949, 16'ha94a, 16'ha94b, 16'ha94c, 16'ha94d, 16'ha94e, 16'ha94f 	:	val_out <= 16'h1363;
         16'ha950, 16'ha951, 16'ha952, 16'ha953, 16'ha954, 16'ha955, 16'ha956, 16'ha957 	:	val_out <= 16'h1356;
         16'ha958, 16'ha959, 16'ha95a, 16'ha95b, 16'ha95c, 16'ha95d, 16'ha95e, 16'ha95f 	:	val_out <= 16'h1348;
         16'ha960, 16'ha961, 16'ha962, 16'ha963, 16'ha964, 16'ha965, 16'ha966, 16'ha967 	:	val_out <= 16'h133b;
         16'ha968, 16'ha969, 16'ha96a, 16'ha96b, 16'ha96c, 16'ha96d, 16'ha96e, 16'ha96f 	:	val_out <= 16'h132e;
         16'ha970, 16'ha971, 16'ha972, 16'ha973, 16'ha974, 16'ha975, 16'ha976, 16'ha977 	:	val_out <= 16'h1321;
         16'ha978, 16'ha979, 16'ha97a, 16'ha97b, 16'ha97c, 16'ha97d, 16'ha97e, 16'ha97f 	:	val_out <= 16'h1313;
         16'ha980, 16'ha981, 16'ha982, 16'ha983, 16'ha984, 16'ha985, 16'ha986, 16'ha987 	:	val_out <= 16'h1306;
         16'ha988, 16'ha989, 16'ha98a, 16'ha98b, 16'ha98c, 16'ha98d, 16'ha98e, 16'ha98f 	:	val_out <= 16'h12f9;
         16'ha990, 16'ha991, 16'ha992, 16'ha993, 16'ha994, 16'ha995, 16'ha996, 16'ha997 	:	val_out <= 16'h12ec;
         16'ha998, 16'ha999, 16'ha99a, 16'ha99b, 16'ha99c, 16'ha99d, 16'ha99e, 16'ha99f 	:	val_out <= 16'h12df;
         16'ha9a0, 16'ha9a1, 16'ha9a2, 16'ha9a3, 16'ha9a4, 16'ha9a5, 16'ha9a6, 16'ha9a7 	:	val_out <= 16'h12d2;
         16'ha9a8, 16'ha9a9, 16'ha9aa, 16'ha9ab, 16'ha9ac, 16'ha9ad, 16'ha9ae, 16'ha9af 	:	val_out <= 16'h12c5;
         16'ha9b0, 16'ha9b1, 16'ha9b2, 16'ha9b3, 16'ha9b4, 16'ha9b5, 16'ha9b6, 16'ha9b7 	:	val_out <= 16'h12b7;
         16'ha9b8, 16'ha9b9, 16'ha9ba, 16'ha9bb, 16'ha9bc, 16'ha9bd, 16'ha9be, 16'ha9bf 	:	val_out <= 16'h12aa;
         16'ha9c0, 16'ha9c1, 16'ha9c2, 16'ha9c3, 16'ha9c4, 16'ha9c5, 16'ha9c6, 16'ha9c7 	:	val_out <= 16'h129d;
         16'ha9c8, 16'ha9c9, 16'ha9ca, 16'ha9cb, 16'ha9cc, 16'ha9cd, 16'ha9ce, 16'ha9cf 	:	val_out <= 16'h1290;
         16'ha9d0, 16'ha9d1, 16'ha9d2, 16'ha9d3, 16'ha9d4, 16'ha9d5, 16'ha9d6, 16'ha9d7 	:	val_out <= 16'h1283;
         16'ha9d8, 16'ha9d9, 16'ha9da, 16'ha9db, 16'ha9dc, 16'ha9dd, 16'ha9de, 16'ha9df 	:	val_out <= 16'h1276;
         16'ha9e0, 16'ha9e1, 16'ha9e2, 16'ha9e3, 16'ha9e4, 16'ha9e5, 16'ha9e6, 16'ha9e7 	:	val_out <= 16'h1269;
         16'ha9e8, 16'ha9e9, 16'ha9ea, 16'ha9eb, 16'ha9ec, 16'ha9ed, 16'ha9ee, 16'ha9ef 	:	val_out <= 16'h125c;
         16'ha9f0, 16'ha9f1, 16'ha9f2, 16'ha9f3, 16'ha9f4, 16'ha9f5, 16'ha9f6, 16'ha9f7 	:	val_out <= 16'h124f;
         16'ha9f8, 16'ha9f9, 16'ha9fa, 16'ha9fb, 16'ha9fc, 16'ha9fd, 16'ha9fe, 16'ha9ff 	:	val_out <= 16'h1242;
         16'haa00, 16'haa01, 16'haa02, 16'haa03, 16'haa04, 16'haa05, 16'haa06, 16'haa07 	:	val_out <= 16'h1235;
         16'haa08, 16'haa09, 16'haa0a, 16'haa0b, 16'haa0c, 16'haa0d, 16'haa0e, 16'haa0f 	:	val_out <= 16'h1229;
         16'haa10, 16'haa11, 16'haa12, 16'haa13, 16'haa14, 16'haa15, 16'haa16, 16'haa17 	:	val_out <= 16'h121c;
         16'haa18, 16'haa19, 16'haa1a, 16'haa1b, 16'haa1c, 16'haa1d, 16'haa1e, 16'haa1f 	:	val_out <= 16'h120f;
         16'haa20, 16'haa21, 16'haa22, 16'haa23, 16'haa24, 16'haa25, 16'haa26, 16'haa27 	:	val_out <= 16'h1202;
         16'haa28, 16'haa29, 16'haa2a, 16'haa2b, 16'haa2c, 16'haa2d, 16'haa2e, 16'haa2f 	:	val_out <= 16'h11f5;
         16'haa30, 16'haa31, 16'haa32, 16'haa33, 16'haa34, 16'haa35, 16'haa36, 16'haa37 	:	val_out <= 16'h11e8;
         16'haa38, 16'haa39, 16'haa3a, 16'haa3b, 16'haa3c, 16'haa3d, 16'haa3e, 16'haa3f 	:	val_out <= 16'h11db;
         16'haa40, 16'haa41, 16'haa42, 16'haa43, 16'haa44, 16'haa45, 16'haa46, 16'haa47 	:	val_out <= 16'h11cf;
         16'haa48, 16'haa49, 16'haa4a, 16'haa4b, 16'haa4c, 16'haa4d, 16'haa4e, 16'haa4f 	:	val_out <= 16'h11c2;
         16'haa50, 16'haa51, 16'haa52, 16'haa53, 16'haa54, 16'haa55, 16'haa56, 16'haa57 	:	val_out <= 16'h11b5;
         16'haa58, 16'haa59, 16'haa5a, 16'haa5b, 16'haa5c, 16'haa5d, 16'haa5e, 16'haa5f 	:	val_out <= 16'h11a8;
         16'haa60, 16'haa61, 16'haa62, 16'haa63, 16'haa64, 16'haa65, 16'haa66, 16'haa67 	:	val_out <= 16'h119c;
         16'haa68, 16'haa69, 16'haa6a, 16'haa6b, 16'haa6c, 16'haa6d, 16'haa6e, 16'haa6f 	:	val_out <= 16'h118f;
         16'haa70, 16'haa71, 16'haa72, 16'haa73, 16'haa74, 16'haa75, 16'haa76, 16'haa77 	:	val_out <= 16'h1182;
         16'haa78, 16'haa79, 16'haa7a, 16'haa7b, 16'haa7c, 16'haa7d, 16'haa7e, 16'haa7f 	:	val_out <= 16'h1176;
         16'haa80, 16'haa81, 16'haa82, 16'haa83, 16'haa84, 16'haa85, 16'haa86, 16'haa87 	:	val_out <= 16'h1169;
         16'haa88, 16'haa89, 16'haa8a, 16'haa8b, 16'haa8c, 16'haa8d, 16'haa8e, 16'haa8f 	:	val_out <= 16'h115c;
         16'haa90, 16'haa91, 16'haa92, 16'haa93, 16'haa94, 16'haa95, 16'haa96, 16'haa97 	:	val_out <= 16'h1150;
         16'haa98, 16'haa99, 16'haa9a, 16'haa9b, 16'haa9c, 16'haa9d, 16'haa9e, 16'haa9f 	:	val_out <= 16'h1143;
         16'haaa0, 16'haaa1, 16'haaa2, 16'haaa3, 16'haaa4, 16'haaa5, 16'haaa6, 16'haaa7 	:	val_out <= 16'h1136;
         16'haaa8, 16'haaa9, 16'haaaa, 16'haaab, 16'haaac, 16'haaad, 16'haaae, 16'haaaf 	:	val_out <= 16'h112a;
         16'haab0, 16'haab1, 16'haab2, 16'haab3, 16'haab4, 16'haab5, 16'haab6, 16'haab7 	:	val_out <= 16'h111d;
         16'haab8, 16'haab9, 16'haaba, 16'haabb, 16'haabc, 16'haabd, 16'haabe, 16'haabf 	:	val_out <= 16'h1111;
         16'haac0, 16'haac1, 16'haac2, 16'haac3, 16'haac4, 16'haac5, 16'haac6, 16'haac7 	:	val_out <= 16'h1104;
         16'haac8, 16'haac9, 16'haaca, 16'haacb, 16'haacc, 16'haacd, 16'haace, 16'haacf 	:	val_out <= 16'h10f8;
         16'haad0, 16'haad1, 16'haad2, 16'haad3, 16'haad4, 16'haad5, 16'haad6, 16'haad7 	:	val_out <= 16'h10eb;
         16'haad8, 16'haad9, 16'haada, 16'haadb, 16'haadc, 16'haadd, 16'haade, 16'haadf 	:	val_out <= 16'h10df;
         16'haae0, 16'haae1, 16'haae2, 16'haae3, 16'haae4, 16'haae5, 16'haae6, 16'haae7 	:	val_out <= 16'h10d2;
         16'haae8, 16'haae9, 16'haaea, 16'haaeb, 16'haaec, 16'haaed, 16'haaee, 16'haaef 	:	val_out <= 16'h10c6;
         16'haaf0, 16'haaf1, 16'haaf2, 16'haaf3, 16'haaf4, 16'haaf5, 16'haaf6, 16'haaf7 	:	val_out <= 16'h10b9;
         16'haaf8, 16'haaf9, 16'haafa, 16'haafb, 16'haafc, 16'haafd, 16'haafe, 16'haaff 	:	val_out <= 16'h10ad;
         16'hab00, 16'hab01, 16'hab02, 16'hab03, 16'hab04, 16'hab05, 16'hab06, 16'hab07 	:	val_out <= 16'h10a0;
         16'hab08, 16'hab09, 16'hab0a, 16'hab0b, 16'hab0c, 16'hab0d, 16'hab0e, 16'hab0f 	:	val_out <= 16'h1094;
         16'hab10, 16'hab11, 16'hab12, 16'hab13, 16'hab14, 16'hab15, 16'hab16, 16'hab17 	:	val_out <= 16'h1088;
         16'hab18, 16'hab19, 16'hab1a, 16'hab1b, 16'hab1c, 16'hab1d, 16'hab1e, 16'hab1f 	:	val_out <= 16'h107b;
         16'hab20, 16'hab21, 16'hab22, 16'hab23, 16'hab24, 16'hab25, 16'hab26, 16'hab27 	:	val_out <= 16'h106f;
         16'hab28, 16'hab29, 16'hab2a, 16'hab2b, 16'hab2c, 16'hab2d, 16'hab2e, 16'hab2f 	:	val_out <= 16'h1063;
         16'hab30, 16'hab31, 16'hab32, 16'hab33, 16'hab34, 16'hab35, 16'hab36, 16'hab37 	:	val_out <= 16'h1056;
         16'hab38, 16'hab39, 16'hab3a, 16'hab3b, 16'hab3c, 16'hab3d, 16'hab3e, 16'hab3f 	:	val_out <= 16'h104a;
         16'hab40, 16'hab41, 16'hab42, 16'hab43, 16'hab44, 16'hab45, 16'hab46, 16'hab47 	:	val_out <= 16'h103e;
         16'hab48, 16'hab49, 16'hab4a, 16'hab4b, 16'hab4c, 16'hab4d, 16'hab4e, 16'hab4f 	:	val_out <= 16'h1032;
         16'hab50, 16'hab51, 16'hab52, 16'hab53, 16'hab54, 16'hab55, 16'hab56, 16'hab57 	:	val_out <= 16'h1025;
         16'hab58, 16'hab59, 16'hab5a, 16'hab5b, 16'hab5c, 16'hab5d, 16'hab5e, 16'hab5f 	:	val_out <= 16'h1019;
         16'hab60, 16'hab61, 16'hab62, 16'hab63, 16'hab64, 16'hab65, 16'hab66, 16'hab67 	:	val_out <= 16'h100d;
         16'hab68, 16'hab69, 16'hab6a, 16'hab6b, 16'hab6c, 16'hab6d, 16'hab6e, 16'hab6f 	:	val_out <= 16'h1001;
         16'hab70, 16'hab71, 16'hab72, 16'hab73, 16'hab74, 16'hab75, 16'hab76, 16'hab77 	:	val_out <= 16'h0ff5;
         16'hab78, 16'hab79, 16'hab7a, 16'hab7b, 16'hab7c, 16'hab7d, 16'hab7e, 16'hab7f 	:	val_out <= 16'h0fe9;
         16'hab80, 16'hab81, 16'hab82, 16'hab83, 16'hab84, 16'hab85, 16'hab86, 16'hab87 	:	val_out <= 16'h0fdc;
         16'hab88, 16'hab89, 16'hab8a, 16'hab8b, 16'hab8c, 16'hab8d, 16'hab8e, 16'hab8f 	:	val_out <= 16'h0fd0;
         16'hab90, 16'hab91, 16'hab92, 16'hab93, 16'hab94, 16'hab95, 16'hab96, 16'hab97 	:	val_out <= 16'h0fc4;
         16'hab98, 16'hab99, 16'hab9a, 16'hab9b, 16'hab9c, 16'hab9d, 16'hab9e, 16'hab9f 	:	val_out <= 16'h0fb8;
         16'haba0, 16'haba1, 16'haba2, 16'haba3, 16'haba4, 16'haba5, 16'haba6, 16'haba7 	:	val_out <= 16'h0fac;
         16'haba8, 16'haba9, 16'habaa, 16'habab, 16'habac, 16'habad, 16'habae, 16'habaf 	:	val_out <= 16'h0fa0;
         16'habb0, 16'habb1, 16'habb2, 16'habb3, 16'habb4, 16'habb5, 16'habb6, 16'habb7 	:	val_out <= 16'h0f94;
         16'habb8, 16'habb9, 16'habba, 16'habbb, 16'habbc, 16'habbd, 16'habbe, 16'habbf 	:	val_out <= 16'h0f88;
         16'habc0, 16'habc1, 16'habc2, 16'habc3, 16'habc4, 16'habc5, 16'habc6, 16'habc7 	:	val_out <= 16'h0f7c;
         16'habc8, 16'habc9, 16'habca, 16'habcb, 16'habcc, 16'habcd, 16'habce, 16'habcf 	:	val_out <= 16'h0f70;
         16'habd0, 16'habd1, 16'habd2, 16'habd3, 16'habd4, 16'habd5, 16'habd6, 16'habd7 	:	val_out <= 16'h0f64;
         16'habd8, 16'habd9, 16'habda, 16'habdb, 16'habdc, 16'habdd, 16'habde, 16'habdf 	:	val_out <= 16'h0f58;
         16'habe0, 16'habe1, 16'habe2, 16'habe3, 16'habe4, 16'habe5, 16'habe6, 16'habe7 	:	val_out <= 16'h0f4c;
         16'habe8, 16'habe9, 16'habea, 16'habeb, 16'habec, 16'habed, 16'habee, 16'habef 	:	val_out <= 16'h0f40;
         16'habf0, 16'habf1, 16'habf2, 16'habf3, 16'habf4, 16'habf5, 16'habf6, 16'habf7 	:	val_out <= 16'h0f34;
         16'habf8, 16'habf9, 16'habfa, 16'habfb, 16'habfc, 16'habfd, 16'habfe, 16'habff 	:	val_out <= 16'h0f29;
         16'hac00, 16'hac01, 16'hac02, 16'hac03, 16'hac04, 16'hac05, 16'hac06, 16'hac07 	:	val_out <= 16'h0f1d;
         16'hac08, 16'hac09, 16'hac0a, 16'hac0b, 16'hac0c, 16'hac0d, 16'hac0e, 16'hac0f 	:	val_out <= 16'h0f11;
         16'hac10, 16'hac11, 16'hac12, 16'hac13, 16'hac14, 16'hac15, 16'hac16, 16'hac17 	:	val_out <= 16'h0f05;
         16'hac18, 16'hac19, 16'hac1a, 16'hac1b, 16'hac1c, 16'hac1d, 16'hac1e, 16'hac1f 	:	val_out <= 16'h0ef9;
         16'hac20, 16'hac21, 16'hac22, 16'hac23, 16'hac24, 16'hac25, 16'hac26, 16'hac27 	:	val_out <= 16'h0eed;
         16'hac28, 16'hac29, 16'hac2a, 16'hac2b, 16'hac2c, 16'hac2d, 16'hac2e, 16'hac2f 	:	val_out <= 16'h0ee2;
         16'hac30, 16'hac31, 16'hac32, 16'hac33, 16'hac34, 16'hac35, 16'hac36, 16'hac37 	:	val_out <= 16'h0ed6;
         16'hac38, 16'hac39, 16'hac3a, 16'hac3b, 16'hac3c, 16'hac3d, 16'hac3e, 16'hac3f 	:	val_out <= 16'h0eca;
         16'hac40, 16'hac41, 16'hac42, 16'hac43, 16'hac44, 16'hac45, 16'hac46, 16'hac47 	:	val_out <= 16'h0ebe;
         16'hac48, 16'hac49, 16'hac4a, 16'hac4b, 16'hac4c, 16'hac4d, 16'hac4e, 16'hac4f 	:	val_out <= 16'h0eb3;
         16'hac50, 16'hac51, 16'hac52, 16'hac53, 16'hac54, 16'hac55, 16'hac56, 16'hac57 	:	val_out <= 16'h0ea7;
         16'hac58, 16'hac59, 16'hac5a, 16'hac5b, 16'hac5c, 16'hac5d, 16'hac5e, 16'hac5f 	:	val_out <= 16'h0e9b;
         16'hac60, 16'hac61, 16'hac62, 16'hac63, 16'hac64, 16'hac65, 16'hac66, 16'hac67 	:	val_out <= 16'h0e90;
         16'hac68, 16'hac69, 16'hac6a, 16'hac6b, 16'hac6c, 16'hac6d, 16'hac6e, 16'hac6f 	:	val_out <= 16'h0e84;
         16'hac70, 16'hac71, 16'hac72, 16'hac73, 16'hac74, 16'hac75, 16'hac76, 16'hac77 	:	val_out <= 16'h0e79;
         16'hac78, 16'hac79, 16'hac7a, 16'hac7b, 16'hac7c, 16'hac7d, 16'hac7e, 16'hac7f 	:	val_out <= 16'h0e6d;
         16'hac80, 16'hac81, 16'hac82, 16'hac83, 16'hac84, 16'hac85, 16'hac86, 16'hac87 	:	val_out <= 16'h0e61;
         16'hac88, 16'hac89, 16'hac8a, 16'hac8b, 16'hac8c, 16'hac8d, 16'hac8e, 16'hac8f 	:	val_out <= 16'h0e56;
         16'hac90, 16'hac91, 16'hac92, 16'hac93, 16'hac94, 16'hac95, 16'hac96, 16'hac97 	:	val_out <= 16'h0e4a;
         16'hac98, 16'hac99, 16'hac9a, 16'hac9b, 16'hac9c, 16'hac9d, 16'hac9e, 16'hac9f 	:	val_out <= 16'h0e3f;
         16'haca0, 16'haca1, 16'haca2, 16'haca3, 16'haca4, 16'haca5, 16'haca6, 16'haca7 	:	val_out <= 16'h0e33;
         16'haca8, 16'haca9, 16'hacaa, 16'hacab, 16'hacac, 16'hacad, 16'hacae, 16'hacaf 	:	val_out <= 16'h0e28;
         16'hacb0, 16'hacb1, 16'hacb2, 16'hacb3, 16'hacb4, 16'hacb5, 16'hacb6, 16'hacb7 	:	val_out <= 16'h0e1c;
         16'hacb8, 16'hacb9, 16'hacba, 16'hacbb, 16'hacbc, 16'hacbd, 16'hacbe, 16'hacbf 	:	val_out <= 16'h0e11;
         16'hacc0, 16'hacc1, 16'hacc2, 16'hacc3, 16'hacc4, 16'hacc5, 16'hacc6, 16'hacc7 	:	val_out <= 16'h0e05;
         16'hacc8, 16'hacc9, 16'hacca, 16'haccb, 16'haccc, 16'haccd, 16'hacce, 16'haccf 	:	val_out <= 16'h0dfa;
         16'hacd0, 16'hacd1, 16'hacd2, 16'hacd3, 16'hacd4, 16'hacd5, 16'hacd6, 16'hacd7 	:	val_out <= 16'h0dee;
         16'hacd8, 16'hacd9, 16'hacda, 16'hacdb, 16'hacdc, 16'hacdd, 16'hacde, 16'hacdf 	:	val_out <= 16'h0de3;
         16'hace0, 16'hace1, 16'hace2, 16'hace3, 16'hace4, 16'hace5, 16'hace6, 16'hace7 	:	val_out <= 16'h0dd8;
         16'hace8, 16'hace9, 16'hacea, 16'haceb, 16'hacec, 16'haced, 16'hacee, 16'hacef 	:	val_out <= 16'h0dcc;
         16'hacf0, 16'hacf1, 16'hacf2, 16'hacf3, 16'hacf4, 16'hacf5, 16'hacf6, 16'hacf7 	:	val_out <= 16'h0dc1;
         16'hacf8, 16'hacf9, 16'hacfa, 16'hacfb, 16'hacfc, 16'hacfd, 16'hacfe, 16'hacff 	:	val_out <= 16'h0db6;
         16'had00, 16'had01, 16'had02, 16'had03, 16'had04, 16'had05, 16'had06, 16'had07 	:	val_out <= 16'h0daa;
         16'had08, 16'had09, 16'had0a, 16'had0b, 16'had0c, 16'had0d, 16'had0e, 16'had0f 	:	val_out <= 16'h0d9f;
         16'had10, 16'had11, 16'had12, 16'had13, 16'had14, 16'had15, 16'had16, 16'had17 	:	val_out <= 16'h0d94;
         16'had18, 16'had19, 16'had1a, 16'had1b, 16'had1c, 16'had1d, 16'had1e, 16'had1f 	:	val_out <= 16'h0d89;
         16'had20, 16'had21, 16'had22, 16'had23, 16'had24, 16'had25, 16'had26, 16'had27 	:	val_out <= 16'h0d7d;
         16'had28, 16'had29, 16'had2a, 16'had2b, 16'had2c, 16'had2d, 16'had2e, 16'had2f 	:	val_out <= 16'h0d72;
         16'had30, 16'had31, 16'had32, 16'had33, 16'had34, 16'had35, 16'had36, 16'had37 	:	val_out <= 16'h0d67;
         16'had38, 16'had39, 16'had3a, 16'had3b, 16'had3c, 16'had3d, 16'had3e, 16'had3f 	:	val_out <= 16'h0d5c;
         16'had40, 16'had41, 16'had42, 16'had43, 16'had44, 16'had45, 16'had46, 16'had47 	:	val_out <= 16'h0d50;
         16'had48, 16'had49, 16'had4a, 16'had4b, 16'had4c, 16'had4d, 16'had4e, 16'had4f 	:	val_out <= 16'h0d45;
         16'had50, 16'had51, 16'had52, 16'had53, 16'had54, 16'had55, 16'had56, 16'had57 	:	val_out <= 16'h0d3a;
         16'had58, 16'had59, 16'had5a, 16'had5b, 16'had5c, 16'had5d, 16'had5e, 16'had5f 	:	val_out <= 16'h0d2f;
         16'had60, 16'had61, 16'had62, 16'had63, 16'had64, 16'had65, 16'had66, 16'had67 	:	val_out <= 16'h0d24;
         16'had68, 16'had69, 16'had6a, 16'had6b, 16'had6c, 16'had6d, 16'had6e, 16'had6f 	:	val_out <= 16'h0d19;
         16'had70, 16'had71, 16'had72, 16'had73, 16'had74, 16'had75, 16'had76, 16'had77 	:	val_out <= 16'h0d0e;
         16'had78, 16'had79, 16'had7a, 16'had7b, 16'had7c, 16'had7d, 16'had7e, 16'had7f 	:	val_out <= 16'h0d03;
         16'had80, 16'had81, 16'had82, 16'had83, 16'had84, 16'had85, 16'had86, 16'had87 	:	val_out <= 16'h0cf8;
         16'had88, 16'had89, 16'had8a, 16'had8b, 16'had8c, 16'had8d, 16'had8e, 16'had8f 	:	val_out <= 16'h0ced;
         16'had90, 16'had91, 16'had92, 16'had93, 16'had94, 16'had95, 16'had96, 16'had97 	:	val_out <= 16'h0ce2;
         16'had98, 16'had99, 16'had9a, 16'had9b, 16'had9c, 16'had9d, 16'had9e, 16'had9f 	:	val_out <= 16'h0cd7;
         16'hada0, 16'hada1, 16'hada2, 16'hada3, 16'hada4, 16'hada5, 16'hada6, 16'hada7 	:	val_out <= 16'h0ccc;
         16'hada8, 16'hada9, 16'hadaa, 16'hadab, 16'hadac, 16'hadad, 16'hadae, 16'hadaf 	:	val_out <= 16'h0cc1;
         16'hadb0, 16'hadb1, 16'hadb2, 16'hadb3, 16'hadb4, 16'hadb5, 16'hadb6, 16'hadb7 	:	val_out <= 16'h0cb6;
         16'hadb8, 16'hadb9, 16'hadba, 16'hadbb, 16'hadbc, 16'hadbd, 16'hadbe, 16'hadbf 	:	val_out <= 16'h0cab;
         16'hadc0, 16'hadc1, 16'hadc2, 16'hadc3, 16'hadc4, 16'hadc5, 16'hadc6, 16'hadc7 	:	val_out <= 16'h0ca0;
         16'hadc8, 16'hadc9, 16'hadca, 16'hadcb, 16'hadcc, 16'hadcd, 16'hadce, 16'hadcf 	:	val_out <= 16'h0c95;
         16'hadd0, 16'hadd1, 16'hadd2, 16'hadd3, 16'hadd4, 16'hadd5, 16'hadd6, 16'hadd7 	:	val_out <= 16'h0c8a;
         16'hadd8, 16'hadd9, 16'hadda, 16'haddb, 16'haddc, 16'haddd, 16'hadde, 16'haddf 	:	val_out <= 16'h0c80;
         16'hade0, 16'hade1, 16'hade2, 16'hade3, 16'hade4, 16'hade5, 16'hade6, 16'hade7 	:	val_out <= 16'h0c75;
         16'hade8, 16'hade9, 16'hadea, 16'hadeb, 16'hadec, 16'haded, 16'hadee, 16'hadef 	:	val_out <= 16'h0c6a;
         16'hadf0, 16'hadf1, 16'hadf2, 16'hadf3, 16'hadf4, 16'hadf5, 16'hadf6, 16'hadf7 	:	val_out <= 16'h0c5f;
         16'hadf8, 16'hadf9, 16'hadfa, 16'hadfb, 16'hadfc, 16'hadfd, 16'hadfe, 16'hadff 	:	val_out <= 16'h0c54;
         16'hae00, 16'hae01, 16'hae02, 16'hae03, 16'hae04, 16'hae05, 16'hae06, 16'hae07 	:	val_out <= 16'h0c4a;
         16'hae08, 16'hae09, 16'hae0a, 16'hae0b, 16'hae0c, 16'hae0d, 16'hae0e, 16'hae0f 	:	val_out <= 16'h0c3f;
         16'hae10, 16'hae11, 16'hae12, 16'hae13, 16'hae14, 16'hae15, 16'hae16, 16'hae17 	:	val_out <= 16'h0c34;
         16'hae18, 16'hae19, 16'hae1a, 16'hae1b, 16'hae1c, 16'hae1d, 16'hae1e, 16'hae1f 	:	val_out <= 16'h0c29;
         16'hae20, 16'hae21, 16'hae22, 16'hae23, 16'hae24, 16'hae25, 16'hae26, 16'hae27 	:	val_out <= 16'h0c1f;
         16'hae28, 16'hae29, 16'hae2a, 16'hae2b, 16'hae2c, 16'hae2d, 16'hae2e, 16'hae2f 	:	val_out <= 16'h0c14;
         16'hae30, 16'hae31, 16'hae32, 16'hae33, 16'hae34, 16'hae35, 16'hae36, 16'hae37 	:	val_out <= 16'h0c09;
         16'hae38, 16'hae39, 16'hae3a, 16'hae3b, 16'hae3c, 16'hae3d, 16'hae3e, 16'hae3f 	:	val_out <= 16'h0bff;
         16'hae40, 16'hae41, 16'hae42, 16'hae43, 16'hae44, 16'hae45, 16'hae46, 16'hae47 	:	val_out <= 16'h0bf4;
         16'hae48, 16'hae49, 16'hae4a, 16'hae4b, 16'hae4c, 16'hae4d, 16'hae4e, 16'hae4f 	:	val_out <= 16'h0bea;
         16'hae50, 16'hae51, 16'hae52, 16'hae53, 16'hae54, 16'hae55, 16'hae56, 16'hae57 	:	val_out <= 16'h0bdf;
         16'hae58, 16'hae59, 16'hae5a, 16'hae5b, 16'hae5c, 16'hae5d, 16'hae5e, 16'hae5f 	:	val_out <= 16'h0bd4;
         16'hae60, 16'hae61, 16'hae62, 16'hae63, 16'hae64, 16'hae65, 16'hae66, 16'hae67 	:	val_out <= 16'h0bca;
         16'hae68, 16'hae69, 16'hae6a, 16'hae6b, 16'hae6c, 16'hae6d, 16'hae6e, 16'hae6f 	:	val_out <= 16'h0bbf;
         16'hae70, 16'hae71, 16'hae72, 16'hae73, 16'hae74, 16'hae75, 16'hae76, 16'hae77 	:	val_out <= 16'h0bb5;
         16'hae78, 16'hae79, 16'hae7a, 16'hae7b, 16'hae7c, 16'hae7d, 16'hae7e, 16'hae7f 	:	val_out <= 16'h0baa;
         16'hae80, 16'hae81, 16'hae82, 16'hae83, 16'hae84, 16'hae85, 16'hae86, 16'hae87 	:	val_out <= 16'h0ba0;
         16'hae88, 16'hae89, 16'hae8a, 16'hae8b, 16'hae8c, 16'hae8d, 16'hae8e, 16'hae8f 	:	val_out <= 16'h0b95;
         16'hae90, 16'hae91, 16'hae92, 16'hae93, 16'hae94, 16'hae95, 16'hae96, 16'hae97 	:	val_out <= 16'h0b8b;
         16'hae98, 16'hae99, 16'hae9a, 16'hae9b, 16'hae9c, 16'hae9d, 16'hae9e, 16'hae9f 	:	val_out <= 16'h0b81;
         16'haea0, 16'haea1, 16'haea2, 16'haea3, 16'haea4, 16'haea5, 16'haea6, 16'haea7 	:	val_out <= 16'h0b76;
         16'haea8, 16'haea9, 16'haeaa, 16'haeab, 16'haeac, 16'haead, 16'haeae, 16'haeaf 	:	val_out <= 16'h0b6c;
         16'haeb0, 16'haeb1, 16'haeb2, 16'haeb3, 16'haeb4, 16'haeb5, 16'haeb6, 16'haeb7 	:	val_out <= 16'h0b61;
         16'haeb8, 16'haeb9, 16'haeba, 16'haebb, 16'haebc, 16'haebd, 16'haebe, 16'haebf 	:	val_out <= 16'h0b57;
         16'haec0, 16'haec1, 16'haec2, 16'haec3, 16'haec4, 16'haec5, 16'haec6, 16'haec7 	:	val_out <= 16'h0b4d;
         16'haec8, 16'haec9, 16'haeca, 16'haecb, 16'haecc, 16'haecd, 16'haece, 16'haecf 	:	val_out <= 16'h0b42;
         16'haed0, 16'haed1, 16'haed2, 16'haed3, 16'haed4, 16'haed5, 16'haed6, 16'haed7 	:	val_out <= 16'h0b38;
         16'haed8, 16'haed9, 16'haeda, 16'haedb, 16'haedc, 16'haedd, 16'haede, 16'haedf 	:	val_out <= 16'h0b2e;
         16'haee0, 16'haee1, 16'haee2, 16'haee3, 16'haee4, 16'haee5, 16'haee6, 16'haee7 	:	val_out <= 16'h0b24;
         16'haee8, 16'haee9, 16'haeea, 16'haeeb, 16'haeec, 16'haeed, 16'haeee, 16'haeef 	:	val_out <= 16'h0b19;
         16'haef0, 16'haef1, 16'haef2, 16'haef3, 16'haef4, 16'haef5, 16'haef6, 16'haef7 	:	val_out <= 16'h0b0f;
         16'haef8, 16'haef9, 16'haefa, 16'haefb, 16'haefc, 16'haefd, 16'haefe, 16'haeff 	:	val_out <= 16'h0b05;
         16'haf00, 16'haf01, 16'haf02, 16'haf03, 16'haf04, 16'haf05, 16'haf06, 16'haf07 	:	val_out <= 16'h0afb;
         16'haf08, 16'haf09, 16'haf0a, 16'haf0b, 16'haf0c, 16'haf0d, 16'haf0e, 16'haf0f 	:	val_out <= 16'h0af0;
         16'haf10, 16'haf11, 16'haf12, 16'haf13, 16'haf14, 16'haf15, 16'haf16, 16'haf17 	:	val_out <= 16'h0ae6;
         16'haf18, 16'haf19, 16'haf1a, 16'haf1b, 16'haf1c, 16'haf1d, 16'haf1e, 16'haf1f 	:	val_out <= 16'h0adc;
         16'haf20, 16'haf21, 16'haf22, 16'haf23, 16'haf24, 16'haf25, 16'haf26, 16'haf27 	:	val_out <= 16'h0ad2;
         16'haf28, 16'haf29, 16'haf2a, 16'haf2b, 16'haf2c, 16'haf2d, 16'haf2e, 16'haf2f 	:	val_out <= 16'h0ac8;
         16'haf30, 16'haf31, 16'haf32, 16'haf33, 16'haf34, 16'haf35, 16'haf36, 16'haf37 	:	val_out <= 16'h0abe;
         16'haf38, 16'haf39, 16'haf3a, 16'haf3b, 16'haf3c, 16'haf3d, 16'haf3e, 16'haf3f 	:	val_out <= 16'h0ab4;
         16'haf40, 16'haf41, 16'haf42, 16'haf43, 16'haf44, 16'haf45, 16'haf46, 16'haf47 	:	val_out <= 16'h0aaa;
         16'haf48, 16'haf49, 16'haf4a, 16'haf4b, 16'haf4c, 16'haf4d, 16'haf4e, 16'haf4f 	:	val_out <= 16'h0aa0;
         16'haf50, 16'haf51, 16'haf52, 16'haf53, 16'haf54, 16'haf55, 16'haf56, 16'haf57 	:	val_out <= 16'h0a96;
         16'haf58, 16'haf59, 16'haf5a, 16'haf5b, 16'haf5c, 16'haf5d, 16'haf5e, 16'haf5f 	:	val_out <= 16'h0a8c;
         16'haf60, 16'haf61, 16'haf62, 16'haf63, 16'haf64, 16'haf65, 16'haf66, 16'haf67 	:	val_out <= 16'h0a82;
         16'haf68, 16'haf69, 16'haf6a, 16'haf6b, 16'haf6c, 16'haf6d, 16'haf6e, 16'haf6f 	:	val_out <= 16'h0a78;
         16'haf70, 16'haf71, 16'haf72, 16'haf73, 16'haf74, 16'haf75, 16'haf76, 16'haf77 	:	val_out <= 16'h0a6e;
         16'haf78, 16'haf79, 16'haf7a, 16'haf7b, 16'haf7c, 16'haf7d, 16'haf7e, 16'haf7f 	:	val_out <= 16'h0a64;
         16'haf80, 16'haf81, 16'haf82, 16'haf83, 16'haf84, 16'haf85, 16'haf86, 16'haf87 	:	val_out <= 16'h0a5a;
         16'haf88, 16'haf89, 16'haf8a, 16'haf8b, 16'haf8c, 16'haf8d, 16'haf8e, 16'haf8f 	:	val_out <= 16'h0a50;
         16'haf90, 16'haf91, 16'haf92, 16'haf93, 16'haf94, 16'haf95, 16'haf96, 16'haf97 	:	val_out <= 16'h0a46;
         16'haf98, 16'haf99, 16'haf9a, 16'haf9b, 16'haf9c, 16'haf9d, 16'haf9e, 16'haf9f 	:	val_out <= 16'h0a3c;
         16'hafa0, 16'hafa1, 16'hafa2, 16'hafa3, 16'hafa4, 16'hafa5, 16'hafa6, 16'hafa7 	:	val_out <= 16'h0a33;
         16'hafa8, 16'hafa9, 16'hafaa, 16'hafab, 16'hafac, 16'hafad, 16'hafae, 16'hafaf 	:	val_out <= 16'h0a29;
         16'hafb0, 16'hafb1, 16'hafb2, 16'hafb3, 16'hafb4, 16'hafb5, 16'hafb6, 16'hafb7 	:	val_out <= 16'h0a1f;
         16'hafb8, 16'hafb9, 16'hafba, 16'hafbb, 16'hafbc, 16'hafbd, 16'hafbe, 16'hafbf 	:	val_out <= 16'h0a15;
         16'hafc0, 16'hafc1, 16'hafc2, 16'hafc3, 16'hafc4, 16'hafc5, 16'hafc6, 16'hafc7 	:	val_out <= 16'h0a0b;
         16'hafc8, 16'hafc9, 16'hafca, 16'hafcb, 16'hafcc, 16'hafcd, 16'hafce, 16'hafcf 	:	val_out <= 16'h0a02;
         16'hafd0, 16'hafd1, 16'hafd2, 16'hafd3, 16'hafd4, 16'hafd5, 16'hafd6, 16'hafd7 	:	val_out <= 16'h09f8;
         16'hafd8, 16'hafd9, 16'hafda, 16'hafdb, 16'hafdc, 16'hafdd, 16'hafde, 16'hafdf 	:	val_out <= 16'h09ee;
         16'hafe0, 16'hafe1, 16'hafe2, 16'hafe3, 16'hafe4, 16'hafe5, 16'hafe6, 16'hafe7 	:	val_out <= 16'h09e4;
         16'hafe8, 16'hafe9, 16'hafea, 16'hafeb, 16'hafec, 16'hafed, 16'hafee, 16'hafef 	:	val_out <= 16'h09db;
         16'haff0, 16'haff1, 16'haff2, 16'haff3, 16'haff4, 16'haff5, 16'haff6, 16'haff7 	:	val_out <= 16'h09d1;
         16'haff8, 16'haff9, 16'haffa, 16'haffb, 16'haffc, 16'haffd, 16'haffe, 16'hafff 	:	val_out <= 16'h09c7;
         16'hb000, 16'hb001, 16'hb002, 16'hb003, 16'hb004, 16'hb005, 16'hb006, 16'hb007 	:	val_out <= 16'h09be;
         16'hb008, 16'hb009, 16'hb00a, 16'hb00b, 16'hb00c, 16'hb00d, 16'hb00e, 16'hb00f 	:	val_out <= 16'h09b4;
         16'hb010, 16'hb011, 16'hb012, 16'hb013, 16'hb014, 16'hb015, 16'hb016, 16'hb017 	:	val_out <= 16'h09ab;
         16'hb018, 16'hb019, 16'hb01a, 16'hb01b, 16'hb01c, 16'hb01d, 16'hb01e, 16'hb01f 	:	val_out <= 16'h09a1;
         16'hb020, 16'hb021, 16'hb022, 16'hb023, 16'hb024, 16'hb025, 16'hb026, 16'hb027 	:	val_out <= 16'h0997;
         16'hb028, 16'hb029, 16'hb02a, 16'hb02b, 16'hb02c, 16'hb02d, 16'hb02e, 16'hb02f 	:	val_out <= 16'h098e;
         16'hb030, 16'hb031, 16'hb032, 16'hb033, 16'hb034, 16'hb035, 16'hb036, 16'hb037 	:	val_out <= 16'h0984;
         16'hb038, 16'hb039, 16'hb03a, 16'hb03b, 16'hb03c, 16'hb03d, 16'hb03e, 16'hb03f 	:	val_out <= 16'h097b;
         16'hb040, 16'hb041, 16'hb042, 16'hb043, 16'hb044, 16'hb045, 16'hb046, 16'hb047 	:	val_out <= 16'h0971;
         16'hb048, 16'hb049, 16'hb04a, 16'hb04b, 16'hb04c, 16'hb04d, 16'hb04e, 16'hb04f 	:	val_out <= 16'h0968;
         16'hb050, 16'hb051, 16'hb052, 16'hb053, 16'hb054, 16'hb055, 16'hb056, 16'hb057 	:	val_out <= 16'h095f;
         16'hb058, 16'hb059, 16'hb05a, 16'hb05b, 16'hb05c, 16'hb05d, 16'hb05e, 16'hb05f 	:	val_out <= 16'h0955;
         16'hb060, 16'hb061, 16'hb062, 16'hb063, 16'hb064, 16'hb065, 16'hb066, 16'hb067 	:	val_out <= 16'h094c;
         16'hb068, 16'hb069, 16'hb06a, 16'hb06b, 16'hb06c, 16'hb06d, 16'hb06e, 16'hb06f 	:	val_out <= 16'h0942;
         16'hb070, 16'hb071, 16'hb072, 16'hb073, 16'hb074, 16'hb075, 16'hb076, 16'hb077 	:	val_out <= 16'h0939;
         16'hb078, 16'hb079, 16'hb07a, 16'hb07b, 16'hb07c, 16'hb07d, 16'hb07e, 16'hb07f 	:	val_out <= 16'h0930;
         16'hb080, 16'hb081, 16'hb082, 16'hb083, 16'hb084, 16'hb085, 16'hb086, 16'hb087 	:	val_out <= 16'h0926;
         16'hb088, 16'hb089, 16'hb08a, 16'hb08b, 16'hb08c, 16'hb08d, 16'hb08e, 16'hb08f 	:	val_out <= 16'h091d;
         16'hb090, 16'hb091, 16'hb092, 16'hb093, 16'hb094, 16'hb095, 16'hb096, 16'hb097 	:	val_out <= 16'h0914;
         16'hb098, 16'hb099, 16'hb09a, 16'hb09b, 16'hb09c, 16'hb09d, 16'hb09e, 16'hb09f 	:	val_out <= 16'h090a;
         16'hb0a0, 16'hb0a1, 16'hb0a2, 16'hb0a3, 16'hb0a4, 16'hb0a5, 16'hb0a6, 16'hb0a7 	:	val_out <= 16'h0901;
         16'hb0a8, 16'hb0a9, 16'hb0aa, 16'hb0ab, 16'hb0ac, 16'hb0ad, 16'hb0ae, 16'hb0af 	:	val_out <= 16'h08f8;
         16'hb0b0, 16'hb0b1, 16'hb0b2, 16'hb0b3, 16'hb0b4, 16'hb0b5, 16'hb0b6, 16'hb0b7 	:	val_out <= 16'h08ef;
         16'hb0b8, 16'hb0b9, 16'hb0ba, 16'hb0bb, 16'hb0bc, 16'hb0bd, 16'hb0be, 16'hb0bf 	:	val_out <= 16'h08e5;
         16'hb0c0, 16'hb0c1, 16'hb0c2, 16'hb0c3, 16'hb0c4, 16'hb0c5, 16'hb0c6, 16'hb0c7 	:	val_out <= 16'h08dc;
         16'hb0c8, 16'hb0c9, 16'hb0ca, 16'hb0cb, 16'hb0cc, 16'hb0cd, 16'hb0ce, 16'hb0cf 	:	val_out <= 16'h08d3;
         16'hb0d0, 16'hb0d1, 16'hb0d2, 16'hb0d3, 16'hb0d4, 16'hb0d5, 16'hb0d6, 16'hb0d7 	:	val_out <= 16'h08ca;
         16'hb0d8, 16'hb0d9, 16'hb0da, 16'hb0db, 16'hb0dc, 16'hb0dd, 16'hb0de, 16'hb0df 	:	val_out <= 16'h08c1;
         16'hb0e0, 16'hb0e1, 16'hb0e2, 16'hb0e3, 16'hb0e4, 16'hb0e5, 16'hb0e6, 16'hb0e7 	:	val_out <= 16'h08b8;
         16'hb0e8, 16'hb0e9, 16'hb0ea, 16'hb0eb, 16'hb0ec, 16'hb0ed, 16'hb0ee, 16'hb0ef 	:	val_out <= 16'h08ae;
         16'hb0f0, 16'hb0f1, 16'hb0f2, 16'hb0f3, 16'hb0f4, 16'hb0f5, 16'hb0f6, 16'hb0f7 	:	val_out <= 16'h08a5;
         16'hb0f8, 16'hb0f9, 16'hb0fa, 16'hb0fb, 16'hb0fc, 16'hb0fd, 16'hb0fe, 16'hb0ff 	:	val_out <= 16'h089c;
         16'hb100, 16'hb101, 16'hb102, 16'hb103, 16'hb104, 16'hb105, 16'hb106, 16'hb107 	:	val_out <= 16'h0893;
         16'hb108, 16'hb109, 16'hb10a, 16'hb10b, 16'hb10c, 16'hb10d, 16'hb10e, 16'hb10f 	:	val_out <= 16'h088a;
         16'hb110, 16'hb111, 16'hb112, 16'hb113, 16'hb114, 16'hb115, 16'hb116, 16'hb117 	:	val_out <= 16'h0881;
         16'hb118, 16'hb119, 16'hb11a, 16'hb11b, 16'hb11c, 16'hb11d, 16'hb11e, 16'hb11f 	:	val_out <= 16'h0878;
         16'hb120, 16'hb121, 16'hb122, 16'hb123, 16'hb124, 16'hb125, 16'hb126, 16'hb127 	:	val_out <= 16'h086f;
         16'hb128, 16'hb129, 16'hb12a, 16'hb12b, 16'hb12c, 16'hb12d, 16'hb12e, 16'hb12f 	:	val_out <= 16'h0866;
         16'hb130, 16'hb131, 16'hb132, 16'hb133, 16'hb134, 16'hb135, 16'hb136, 16'hb137 	:	val_out <= 16'h085d;
         16'hb138, 16'hb139, 16'hb13a, 16'hb13b, 16'hb13c, 16'hb13d, 16'hb13e, 16'hb13f 	:	val_out <= 16'h0854;
         16'hb140, 16'hb141, 16'hb142, 16'hb143, 16'hb144, 16'hb145, 16'hb146, 16'hb147 	:	val_out <= 16'h084b;
         16'hb148, 16'hb149, 16'hb14a, 16'hb14b, 16'hb14c, 16'hb14d, 16'hb14e, 16'hb14f 	:	val_out <= 16'h0843;
         16'hb150, 16'hb151, 16'hb152, 16'hb153, 16'hb154, 16'hb155, 16'hb156, 16'hb157 	:	val_out <= 16'h083a;
         16'hb158, 16'hb159, 16'hb15a, 16'hb15b, 16'hb15c, 16'hb15d, 16'hb15e, 16'hb15f 	:	val_out <= 16'h0831;
         16'hb160, 16'hb161, 16'hb162, 16'hb163, 16'hb164, 16'hb165, 16'hb166, 16'hb167 	:	val_out <= 16'h0828;
         16'hb168, 16'hb169, 16'hb16a, 16'hb16b, 16'hb16c, 16'hb16d, 16'hb16e, 16'hb16f 	:	val_out <= 16'h081f;
         16'hb170, 16'hb171, 16'hb172, 16'hb173, 16'hb174, 16'hb175, 16'hb176, 16'hb177 	:	val_out <= 16'h0816;
         16'hb178, 16'hb179, 16'hb17a, 16'hb17b, 16'hb17c, 16'hb17d, 16'hb17e, 16'hb17f 	:	val_out <= 16'h080e;
         16'hb180, 16'hb181, 16'hb182, 16'hb183, 16'hb184, 16'hb185, 16'hb186, 16'hb187 	:	val_out <= 16'h0805;
         16'hb188, 16'hb189, 16'hb18a, 16'hb18b, 16'hb18c, 16'hb18d, 16'hb18e, 16'hb18f 	:	val_out <= 16'h07fc;
         16'hb190, 16'hb191, 16'hb192, 16'hb193, 16'hb194, 16'hb195, 16'hb196, 16'hb197 	:	val_out <= 16'h07f3;
         16'hb198, 16'hb199, 16'hb19a, 16'hb19b, 16'hb19c, 16'hb19d, 16'hb19e, 16'hb19f 	:	val_out <= 16'h07eb;
         16'hb1a0, 16'hb1a1, 16'hb1a2, 16'hb1a3, 16'hb1a4, 16'hb1a5, 16'hb1a6, 16'hb1a7 	:	val_out <= 16'h07e2;
         16'hb1a8, 16'hb1a9, 16'hb1aa, 16'hb1ab, 16'hb1ac, 16'hb1ad, 16'hb1ae, 16'hb1af 	:	val_out <= 16'h07d9;
         16'hb1b0, 16'hb1b1, 16'hb1b2, 16'hb1b3, 16'hb1b4, 16'hb1b5, 16'hb1b6, 16'hb1b7 	:	val_out <= 16'h07d1;
         16'hb1b8, 16'hb1b9, 16'hb1ba, 16'hb1bb, 16'hb1bc, 16'hb1bd, 16'hb1be, 16'hb1bf 	:	val_out <= 16'h07c8;
         16'hb1c0, 16'hb1c1, 16'hb1c2, 16'hb1c3, 16'hb1c4, 16'hb1c5, 16'hb1c6, 16'hb1c7 	:	val_out <= 16'h07bf;
         16'hb1c8, 16'hb1c9, 16'hb1ca, 16'hb1cb, 16'hb1cc, 16'hb1cd, 16'hb1ce, 16'hb1cf 	:	val_out <= 16'h07b7;
         16'hb1d0, 16'hb1d1, 16'hb1d2, 16'hb1d3, 16'hb1d4, 16'hb1d5, 16'hb1d6, 16'hb1d7 	:	val_out <= 16'h07ae;
         16'hb1d8, 16'hb1d9, 16'hb1da, 16'hb1db, 16'hb1dc, 16'hb1dd, 16'hb1de, 16'hb1df 	:	val_out <= 16'h07a6;
         16'hb1e0, 16'hb1e1, 16'hb1e2, 16'hb1e3, 16'hb1e4, 16'hb1e5, 16'hb1e6, 16'hb1e7 	:	val_out <= 16'h079d;
         16'hb1e8, 16'hb1e9, 16'hb1ea, 16'hb1eb, 16'hb1ec, 16'hb1ed, 16'hb1ee, 16'hb1ef 	:	val_out <= 16'h0794;
         16'hb1f0, 16'hb1f1, 16'hb1f2, 16'hb1f3, 16'hb1f4, 16'hb1f5, 16'hb1f6, 16'hb1f7 	:	val_out <= 16'h078c;
         16'hb1f8, 16'hb1f9, 16'hb1fa, 16'hb1fb, 16'hb1fc, 16'hb1fd, 16'hb1fe, 16'hb1ff 	:	val_out <= 16'h0783;
         16'hb200, 16'hb201, 16'hb202, 16'hb203, 16'hb204, 16'hb205, 16'hb206, 16'hb207 	:	val_out <= 16'h077b;
         16'hb208, 16'hb209, 16'hb20a, 16'hb20b, 16'hb20c, 16'hb20d, 16'hb20e, 16'hb20f 	:	val_out <= 16'h0773;
         16'hb210, 16'hb211, 16'hb212, 16'hb213, 16'hb214, 16'hb215, 16'hb216, 16'hb217 	:	val_out <= 16'h076a;
         16'hb218, 16'hb219, 16'hb21a, 16'hb21b, 16'hb21c, 16'hb21d, 16'hb21e, 16'hb21f 	:	val_out <= 16'h0762;
         16'hb220, 16'hb221, 16'hb222, 16'hb223, 16'hb224, 16'hb225, 16'hb226, 16'hb227 	:	val_out <= 16'h0759;
         16'hb228, 16'hb229, 16'hb22a, 16'hb22b, 16'hb22c, 16'hb22d, 16'hb22e, 16'hb22f 	:	val_out <= 16'h0751;
         16'hb230, 16'hb231, 16'hb232, 16'hb233, 16'hb234, 16'hb235, 16'hb236, 16'hb237 	:	val_out <= 16'h0749;
         16'hb238, 16'hb239, 16'hb23a, 16'hb23b, 16'hb23c, 16'hb23d, 16'hb23e, 16'hb23f 	:	val_out <= 16'h0740;
         16'hb240, 16'hb241, 16'hb242, 16'hb243, 16'hb244, 16'hb245, 16'hb246, 16'hb247 	:	val_out <= 16'h0738;
         16'hb248, 16'hb249, 16'hb24a, 16'hb24b, 16'hb24c, 16'hb24d, 16'hb24e, 16'hb24f 	:	val_out <= 16'h0730;
         16'hb250, 16'hb251, 16'hb252, 16'hb253, 16'hb254, 16'hb255, 16'hb256, 16'hb257 	:	val_out <= 16'h0727;
         16'hb258, 16'hb259, 16'hb25a, 16'hb25b, 16'hb25c, 16'hb25d, 16'hb25e, 16'hb25f 	:	val_out <= 16'h071f;
         16'hb260, 16'hb261, 16'hb262, 16'hb263, 16'hb264, 16'hb265, 16'hb266, 16'hb267 	:	val_out <= 16'h0717;
         16'hb268, 16'hb269, 16'hb26a, 16'hb26b, 16'hb26c, 16'hb26d, 16'hb26e, 16'hb26f 	:	val_out <= 16'h070e;
         16'hb270, 16'hb271, 16'hb272, 16'hb273, 16'hb274, 16'hb275, 16'hb276, 16'hb277 	:	val_out <= 16'h0706;
         16'hb278, 16'hb279, 16'hb27a, 16'hb27b, 16'hb27c, 16'hb27d, 16'hb27e, 16'hb27f 	:	val_out <= 16'h06fe;
         16'hb280, 16'hb281, 16'hb282, 16'hb283, 16'hb284, 16'hb285, 16'hb286, 16'hb287 	:	val_out <= 16'h06f6;
         16'hb288, 16'hb289, 16'hb28a, 16'hb28b, 16'hb28c, 16'hb28d, 16'hb28e, 16'hb28f 	:	val_out <= 16'h06ee;
         16'hb290, 16'hb291, 16'hb292, 16'hb293, 16'hb294, 16'hb295, 16'hb296, 16'hb297 	:	val_out <= 16'h06e6;
         16'hb298, 16'hb299, 16'hb29a, 16'hb29b, 16'hb29c, 16'hb29d, 16'hb29e, 16'hb29f 	:	val_out <= 16'h06dd;
         16'hb2a0, 16'hb2a1, 16'hb2a2, 16'hb2a3, 16'hb2a4, 16'hb2a5, 16'hb2a6, 16'hb2a7 	:	val_out <= 16'h06d5;
         16'hb2a8, 16'hb2a9, 16'hb2aa, 16'hb2ab, 16'hb2ac, 16'hb2ad, 16'hb2ae, 16'hb2af 	:	val_out <= 16'h06cd;
         16'hb2b0, 16'hb2b1, 16'hb2b2, 16'hb2b3, 16'hb2b4, 16'hb2b5, 16'hb2b6, 16'hb2b7 	:	val_out <= 16'h06c5;
         16'hb2b8, 16'hb2b9, 16'hb2ba, 16'hb2bb, 16'hb2bc, 16'hb2bd, 16'hb2be, 16'hb2bf 	:	val_out <= 16'h06bd;
         16'hb2c0, 16'hb2c1, 16'hb2c2, 16'hb2c3, 16'hb2c4, 16'hb2c5, 16'hb2c6, 16'hb2c7 	:	val_out <= 16'h06b5;
         16'hb2c8, 16'hb2c9, 16'hb2ca, 16'hb2cb, 16'hb2cc, 16'hb2cd, 16'hb2ce, 16'hb2cf 	:	val_out <= 16'h06ad;
         16'hb2d0, 16'hb2d1, 16'hb2d2, 16'hb2d3, 16'hb2d4, 16'hb2d5, 16'hb2d6, 16'hb2d7 	:	val_out <= 16'h06a5;
         16'hb2d8, 16'hb2d9, 16'hb2da, 16'hb2db, 16'hb2dc, 16'hb2dd, 16'hb2de, 16'hb2df 	:	val_out <= 16'h069d;
         16'hb2e0, 16'hb2e1, 16'hb2e2, 16'hb2e3, 16'hb2e4, 16'hb2e5, 16'hb2e6, 16'hb2e7 	:	val_out <= 16'h0695;
         16'hb2e8, 16'hb2e9, 16'hb2ea, 16'hb2eb, 16'hb2ec, 16'hb2ed, 16'hb2ee, 16'hb2ef 	:	val_out <= 16'h068d;
         16'hb2f0, 16'hb2f1, 16'hb2f2, 16'hb2f3, 16'hb2f4, 16'hb2f5, 16'hb2f6, 16'hb2f7 	:	val_out <= 16'h0685;
         16'hb2f8, 16'hb2f9, 16'hb2fa, 16'hb2fb, 16'hb2fc, 16'hb2fd, 16'hb2fe, 16'hb2ff 	:	val_out <= 16'h067d;
         16'hb300, 16'hb301, 16'hb302, 16'hb303, 16'hb304, 16'hb305, 16'hb306, 16'hb307 	:	val_out <= 16'h0675;
         16'hb308, 16'hb309, 16'hb30a, 16'hb30b, 16'hb30c, 16'hb30d, 16'hb30e, 16'hb30f 	:	val_out <= 16'h066d;
         16'hb310, 16'hb311, 16'hb312, 16'hb313, 16'hb314, 16'hb315, 16'hb316, 16'hb317 	:	val_out <= 16'h0666;
         16'hb318, 16'hb319, 16'hb31a, 16'hb31b, 16'hb31c, 16'hb31d, 16'hb31e, 16'hb31f 	:	val_out <= 16'h065e;
         16'hb320, 16'hb321, 16'hb322, 16'hb323, 16'hb324, 16'hb325, 16'hb326, 16'hb327 	:	val_out <= 16'h0656;
         16'hb328, 16'hb329, 16'hb32a, 16'hb32b, 16'hb32c, 16'hb32d, 16'hb32e, 16'hb32f 	:	val_out <= 16'h064e;
         16'hb330, 16'hb331, 16'hb332, 16'hb333, 16'hb334, 16'hb335, 16'hb336, 16'hb337 	:	val_out <= 16'h0646;
         16'hb338, 16'hb339, 16'hb33a, 16'hb33b, 16'hb33c, 16'hb33d, 16'hb33e, 16'hb33f 	:	val_out <= 16'h063f;
         16'hb340, 16'hb341, 16'hb342, 16'hb343, 16'hb344, 16'hb345, 16'hb346, 16'hb347 	:	val_out <= 16'h0637;
         16'hb348, 16'hb349, 16'hb34a, 16'hb34b, 16'hb34c, 16'hb34d, 16'hb34e, 16'hb34f 	:	val_out <= 16'h062f;
         16'hb350, 16'hb351, 16'hb352, 16'hb353, 16'hb354, 16'hb355, 16'hb356, 16'hb357 	:	val_out <= 16'h0627;
         16'hb358, 16'hb359, 16'hb35a, 16'hb35b, 16'hb35c, 16'hb35d, 16'hb35e, 16'hb35f 	:	val_out <= 16'h0620;
         16'hb360, 16'hb361, 16'hb362, 16'hb363, 16'hb364, 16'hb365, 16'hb366, 16'hb367 	:	val_out <= 16'h0618;
         16'hb368, 16'hb369, 16'hb36a, 16'hb36b, 16'hb36c, 16'hb36d, 16'hb36e, 16'hb36f 	:	val_out <= 16'h0610;
         16'hb370, 16'hb371, 16'hb372, 16'hb373, 16'hb374, 16'hb375, 16'hb376, 16'hb377 	:	val_out <= 16'h0609;
         16'hb378, 16'hb379, 16'hb37a, 16'hb37b, 16'hb37c, 16'hb37d, 16'hb37e, 16'hb37f 	:	val_out <= 16'h0601;
         16'hb380, 16'hb381, 16'hb382, 16'hb383, 16'hb384, 16'hb385, 16'hb386, 16'hb387 	:	val_out <= 16'h05fa;
         16'hb388, 16'hb389, 16'hb38a, 16'hb38b, 16'hb38c, 16'hb38d, 16'hb38e, 16'hb38f 	:	val_out <= 16'h05f2;
         16'hb390, 16'hb391, 16'hb392, 16'hb393, 16'hb394, 16'hb395, 16'hb396, 16'hb397 	:	val_out <= 16'h05ea;
         16'hb398, 16'hb399, 16'hb39a, 16'hb39b, 16'hb39c, 16'hb39d, 16'hb39e, 16'hb39f 	:	val_out <= 16'h05e3;
         16'hb3a0, 16'hb3a1, 16'hb3a2, 16'hb3a3, 16'hb3a4, 16'hb3a5, 16'hb3a6, 16'hb3a7 	:	val_out <= 16'h05db;
         16'hb3a8, 16'hb3a9, 16'hb3aa, 16'hb3ab, 16'hb3ac, 16'hb3ad, 16'hb3ae, 16'hb3af 	:	val_out <= 16'h05d4;
         16'hb3b0, 16'hb3b1, 16'hb3b2, 16'hb3b3, 16'hb3b4, 16'hb3b5, 16'hb3b6, 16'hb3b7 	:	val_out <= 16'h05cc;
         16'hb3b8, 16'hb3b9, 16'hb3ba, 16'hb3bb, 16'hb3bc, 16'hb3bd, 16'hb3be, 16'hb3bf 	:	val_out <= 16'h05c5;
         16'hb3c0, 16'hb3c1, 16'hb3c2, 16'hb3c3, 16'hb3c4, 16'hb3c5, 16'hb3c6, 16'hb3c7 	:	val_out <= 16'h05bd;
         16'hb3c8, 16'hb3c9, 16'hb3ca, 16'hb3cb, 16'hb3cc, 16'hb3cd, 16'hb3ce, 16'hb3cf 	:	val_out <= 16'h05b6;
         16'hb3d0, 16'hb3d1, 16'hb3d2, 16'hb3d3, 16'hb3d4, 16'hb3d5, 16'hb3d6, 16'hb3d7 	:	val_out <= 16'h05af;
         16'hb3d8, 16'hb3d9, 16'hb3da, 16'hb3db, 16'hb3dc, 16'hb3dd, 16'hb3de, 16'hb3df 	:	val_out <= 16'h05a7;
         16'hb3e0, 16'hb3e1, 16'hb3e2, 16'hb3e3, 16'hb3e4, 16'hb3e5, 16'hb3e6, 16'hb3e7 	:	val_out <= 16'h05a0;
         16'hb3e8, 16'hb3e9, 16'hb3ea, 16'hb3eb, 16'hb3ec, 16'hb3ed, 16'hb3ee, 16'hb3ef 	:	val_out <= 16'h0598;
         16'hb3f0, 16'hb3f1, 16'hb3f2, 16'hb3f3, 16'hb3f4, 16'hb3f5, 16'hb3f6, 16'hb3f7 	:	val_out <= 16'h0591;
         16'hb3f8, 16'hb3f9, 16'hb3fa, 16'hb3fb, 16'hb3fc, 16'hb3fd, 16'hb3fe, 16'hb3ff 	:	val_out <= 16'h058a;
         16'hb400, 16'hb401, 16'hb402, 16'hb403, 16'hb404, 16'hb405, 16'hb406, 16'hb407 	:	val_out <= 16'h0582;
         16'hb408, 16'hb409, 16'hb40a, 16'hb40b, 16'hb40c, 16'hb40d, 16'hb40e, 16'hb40f 	:	val_out <= 16'h057b;
         16'hb410, 16'hb411, 16'hb412, 16'hb413, 16'hb414, 16'hb415, 16'hb416, 16'hb417 	:	val_out <= 16'h0574;
         16'hb418, 16'hb419, 16'hb41a, 16'hb41b, 16'hb41c, 16'hb41d, 16'hb41e, 16'hb41f 	:	val_out <= 16'h056d;
         16'hb420, 16'hb421, 16'hb422, 16'hb423, 16'hb424, 16'hb425, 16'hb426, 16'hb427 	:	val_out <= 16'h0565;
         16'hb428, 16'hb429, 16'hb42a, 16'hb42b, 16'hb42c, 16'hb42d, 16'hb42e, 16'hb42f 	:	val_out <= 16'h055e;
         16'hb430, 16'hb431, 16'hb432, 16'hb433, 16'hb434, 16'hb435, 16'hb436, 16'hb437 	:	val_out <= 16'h0557;
         16'hb438, 16'hb439, 16'hb43a, 16'hb43b, 16'hb43c, 16'hb43d, 16'hb43e, 16'hb43f 	:	val_out <= 16'h0550;
         16'hb440, 16'hb441, 16'hb442, 16'hb443, 16'hb444, 16'hb445, 16'hb446, 16'hb447 	:	val_out <= 16'h0549;
         16'hb448, 16'hb449, 16'hb44a, 16'hb44b, 16'hb44c, 16'hb44d, 16'hb44e, 16'hb44f 	:	val_out <= 16'h0542;
         16'hb450, 16'hb451, 16'hb452, 16'hb453, 16'hb454, 16'hb455, 16'hb456, 16'hb457 	:	val_out <= 16'h053a;
         16'hb458, 16'hb459, 16'hb45a, 16'hb45b, 16'hb45c, 16'hb45d, 16'hb45e, 16'hb45f 	:	val_out <= 16'h0533;
         16'hb460, 16'hb461, 16'hb462, 16'hb463, 16'hb464, 16'hb465, 16'hb466, 16'hb467 	:	val_out <= 16'h052c;
         16'hb468, 16'hb469, 16'hb46a, 16'hb46b, 16'hb46c, 16'hb46d, 16'hb46e, 16'hb46f 	:	val_out <= 16'h0525;
         16'hb470, 16'hb471, 16'hb472, 16'hb473, 16'hb474, 16'hb475, 16'hb476, 16'hb477 	:	val_out <= 16'h051e;
         16'hb478, 16'hb479, 16'hb47a, 16'hb47b, 16'hb47c, 16'hb47d, 16'hb47e, 16'hb47f 	:	val_out <= 16'h0517;
         16'hb480, 16'hb481, 16'hb482, 16'hb483, 16'hb484, 16'hb485, 16'hb486, 16'hb487 	:	val_out <= 16'h0510;
         16'hb488, 16'hb489, 16'hb48a, 16'hb48b, 16'hb48c, 16'hb48d, 16'hb48e, 16'hb48f 	:	val_out <= 16'h0509;
         16'hb490, 16'hb491, 16'hb492, 16'hb493, 16'hb494, 16'hb495, 16'hb496, 16'hb497 	:	val_out <= 16'h0502;
         16'hb498, 16'hb499, 16'hb49a, 16'hb49b, 16'hb49c, 16'hb49d, 16'hb49e, 16'hb49f 	:	val_out <= 16'h04fb;
         16'hb4a0, 16'hb4a1, 16'hb4a2, 16'hb4a3, 16'hb4a4, 16'hb4a5, 16'hb4a6, 16'hb4a7 	:	val_out <= 16'h04f4;
         16'hb4a8, 16'hb4a9, 16'hb4aa, 16'hb4ab, 16'hb4ac, 16'hb4ad, 16'hb4ae, 16'hb4af 	:	val_out <= 16'h04ed;
         16'hb4b0, 16'hb4b1, 16'hb4b2, 16'hb4b3, 16'hb4b4, 16'hb4b5, 16'hb4b6, 16'hb4b7 	:	val_out <= 16'h04e6;
         16'hb4b8, 16'hb4b9, 16'hb4ba, 16'hb4bb, 16'hb4bc, 16'hb4bd, 16'hb4be, 16'hb4bf 	:	val_out <= 16'h04e0;
         16'hb4c0, 16'hb4c1, 16'hb4c2, 16'hb4c3, 16'hb4c4, 16'hb4c5, 16'hb4c6, 16'hb4c7 	:	val_out <= 16'h04d9;
         16'hb4c8, 16'hb4c9, 16'hb4ca, 16'hb4cb, 16'hb4cc, 16'hb4cd, 16'hb4ce, 16'hb4cf 	:	val_out <= 16'h04d2;
         16'hb4d0, 16'hb4d1, 16'hb4d2, 16'hb4d3, 16'hb4d4, 16'hb4d5, 16'hb4d6, 16'hb4d7 	:	val_out <= 16'h04cb;
         16'hb4d8, 16'hb4d9, 16'hb4da, 16'hb4db, 16'hb4dc, 16'hb4dd, 16'hb4de, 16'hb4df 	:	val_out <= 16'h04c4;
         16'hb4e0, 16'hb4e1, 16'hb4e2, 16'hb4e3, 16'hb4e4, 16'hb4e5, 16'hb4e6, 16'hb4e7 	:	val_out <= 16'h04bd;
         16'hb4e8, 16'hb4e9, 16'hb4ea, 16'hb4eb, 16'hb4ec, 16'hb4ed, 16'hb4ee, 16'hb4ef 	:	val_out <= 16'h04b7;
         16'hb4f0, 16'hb4f1, 16'hb4f2, 16'hb4f3, 16'hb4f4, 16'hb4f5, 16'hb4f6, 16'hb4f7 	:	val_out <= 16'h04b0;
         16'hb4f8, 16'hb4f9, 16'hb4fa, 16'hb4fb, 16'hb4fc, 16'hb4fd, 16'hb4fe, 16'hb4ff 	:	val_out <= 16'h04a9;
         16'hb500, 16'hb501, 16'hb502, 16'hb503, 16'hb504, 16'hb505, 16'hb506, 16'hb507 	:	val_out <= 16'h04a2;
         16'hb508, 16'hb509, 16'hb50a, 16'hb50b, 16'hb50c, 16'hb50d, 16'hb50e, 16'hb50f 	:	val_out <= 16'h049c;
         16'hb510, 16'hb511, 16'hb512, 16'hb513, 16'hb514, 16'hb515, 16'hb516, 16'hb517 	:	val_out <= 16'h0495;
         16'hb518, 16'hb519, 16'hb51a, 16'hb51b, 16'hb51c, 16'hb51d, 16'hb51e, 16'hb51f 	:	val_out <= 16'h048e;
         16'hb520, 16'hb521, 16'hb522, 16'hb523, 16'hb524, 16'hb525, 16'hb526, 16'hb527 	:	val_out <= 16'h0488;
         16'hb528, 16'hb529, 16'hb52a, 16'hb52b, 16'hb52c, 16'hb52d, 16'hb52e, 16'hb52f 	:	val_out <= 16'h0481;
         16'hb530, 16'hb531, 16'hb532, 16'hb533, 16'hb534, 16'hb535, 16'hb536, 16'hb537 	:	val_out <= 16'h047b;
         16'hb538, 16'hb539, 16'hb53a, 16'hb53b, 16'hb53c, 16'hb53d, 16'hb53e, 16'hb53f 	:	val_out <= 16'h0474;
         16'hb540, 16'hb541, 16'hb542, 16'hb543, 16'hb544, 16'hb545, 16'hb546, 16'hb547 	:	val_out <= 16'h046d;
         16'hb548, 16'hb549, 16'hb54a, 16'hb54b, 16'hb54c, 16'hb54d, 16'hb54e, 16'hb54f 	:	val_out <= 16'h0467;
         16'hb550, 16'hb551, 16'hb552, 16'hb553, 16'hb554, 16'hb555, 16'hb556, 16'hb557 	:	val_out <= 16'h0460;
         16'hb558, 16'hb559, 16'hb55a, 16'hb55b, 16'hb55c, 16'hb55d, 16'hb55e, 16'hb55f 	:	val_out <= 16'h045a;
         16'hb560, 16'hb561, 16'hb562, 16'hb563, 16'hb564, 16'hb565, 16'hb566, 16'hb567 	:	val_out <= 16'h0453;
         16'hb568, 16'hb569, 16'hb56a, 16'hb56b, 16'hb56c, 16'hb56d, 16'hb56e, 16'hb56f 	:	val_out <= 16'h044d;
         16'hb570, 16'hb571, 16'hb572, 16'hb573, 16'hb574, 16'hb575, 16'hb576, 16'hb577 	:	val_out <= 16'h0446;
         16'hb578, 16'hb579, 16'hb57a, 16'hb57b, 16'hb57c, 16'hb57d, 16'hb57e, 16'hb57f 	:	val_out <= 16'h0440;
         16'hb580, 16'hb581, 16'hb582, 16'hb583, 16'hb584, 16'hb585, 16'hb586, 16'hb587 	:	val_out <= 16'h043a;
         16'hb588, 16'hb589, 16'hb58a, 16'hb58b, 16'hb58c, 16'hb58d, 16'hb58e, 16'hb58f 	:	val_out <= 16'h0433;
         16'hb590, 16'hb591, 16'hb592, 16'hb593, 16'hb594, 16'hb595, 16'hb596, 16'hb597 	:	val_out <= 16'h042d;
         16'hb598, 16'hb599, 16'hb59a, 16'hb59b, 16'hb59c, 16'hb59d, 16'hb59e, 16'hb59f 	:	val_out <= 16'h0426;
         16'hb5a0, 16'hb5a1, 16'hb5a2, 16'hb5a3, 16'hb5a4, 16'hb5a5, 16'hb5a6, 16'hb5a7 	:	val_out <= 16'h0420;
         16'hb5a8, 16'hb5a9, 16'hb5aa, 16'hb5ab, 16'hb5ac, 16'hb5ad, 16'hb5ae, 16'hb5af 	:	val_out <= 16'h041a;
         16'hb5b0, 16'hb5b1, 16'hb5b2, 16'hb5b3, 16'hb5b4, 16'hb5b5, 16'hb5b6, 16'hb5b7 	:	val_out <= 16'h0414;
         16'hb5b8, 16'hb5b9, 16'hb5ba, 16'hb5bb, 16'hb5bc, 16'hb5bd, 16'hb5be, 16'hb5bf 	:	val_out <= 16'h040d;
         16'hb5c0, 16'hb5c1, 16'hb5c2, 16'hb5c3, 16'hb5c4, 16'hb5c5, 16'hb5c6, 16'hb5c7 	:	val_out <= 16'h0407;
         16'hb5c8, 16'hb5c9, 16'hb5ca, 16'hb5cb, 16'hb5cc, 16'hb5cd, 16'hb5ce, 16'hb5cf 	:	val_out <= 16'h0401;
         16'hb5d0, 16'hb5d1, 16'hb5d2, 16'hb5d3, 16'hb5d4, 16'hb5d5, 16'hb5d6, 16'hb5d7 	:	val_out <= 16'h03fa;
         16'hb5d8, 16'hb5d9, 16'hb5da, 16'hb5db, 16'hb5dc, 16'hb5dd, 16'hb5de, 16'hb5df 	:	val_out <= 16'h03f4;
         16'hb5e0, 16'hb5e1, 16'hb5e2, 16'hb5e3, 16'hb5e4, 16'hb5e5, 16'hb5e6, 16'hb5e7 	:	val_out <= 16'h03ee;
         16'hb5e8, 16'hb5e9, 16'hb5ea, 16'hb5eb, 16'hb5ec, 16'hb5ed, 16'hb5ee, 16'hb5ef 	:	val_out <= 16'h03e8;
         16'hb5f0, 16'hb5f1, 16'hb5f2, 16'hb5f3, 16'hb5f4, 16'hb5f5, 16'hb5f6, 16'hb5f7 	:	val_out <= 16'h03e2;
         16'hb5f8, 16'hb5f9, 16'hb5fa, 16'hb5fb, 16'hb5fc, 16'hb5fd, 16'hb5fe, 16'hb5ff 	:	val_out <= 16'h03dc;
         16'hb600, 16'hb601, 16'hb602, 16'hb603, 16'hb604, 16'hb605, 16'hb606, 16'hb607 	:	val_out <= 16'h03d6;
         16'hb608, 16'hb609, 16'hb60a, 16'hb60b, 16'hb60c, 16'hb60d, 16'hb60e, 16'hb60f 	:	val_out <= 16'h03cf;
         16'hb610, 16'hb611, 16'hb612, 16'hb613, 16'hb614, 16'hb615, 16'hb616, 16'hb617 	:	val_out <= 16'h03c9;
         16'hb618, 16'hb619, 16'hb61a, 16'hb61b, 16'hb61c, 16'hb61d, 16'hb61e, 16'hb61f 	:	val_out <= 16'h03c3;
         16'hb620, 16'hb621, 16'hb622, 16'hb623, 16'hb624, 16'hb625, 16'hb626, 16'hb627 	:	val_out <= 16'h03bd;
         16'hb628, 16'hb629, 16'hb62a, 16'hb62b, 16'hb62c, 16'hb62d, 16'hb62e, 16'hb62f 	:	val_out <= 16'h03b7;
         16'hb630, 16'hb631, 16'hb632, 16'hb633, 16'hb634, 16'hb635, 16'hb636, 16'hb637 	:	val_out <= 16'h03b1;
         16'hb638, 16'hb639, 16'hb63a, 16'hb63b, 16'hb63c, 16'hb63d, 16'hb63e, 16'hb63f 	:	val_out <= 16'h03ab;
         16'hb640, 16'hb641, 16'hb642, 16'hb643, 16'hb644, 16'hb645, 16'hb646, 16'hb647 	:	val_out <= 16'h03a5;
         16'hb648, 16'hb649, 16'hb64a, 16'hb64b, 16'hb64c, 16'hb64d, 16'hb64e, 16'hb64f 	:	val_out <= 16'h039f;
         16'hb650, 16'hb651, 16'hb652, 16'hb653, 16'hb654, 16'hb655, 16'hb656, 16'hb657 	:	val_out <= 16'h0399;
         16'hb658, 16'hb659, 16'hb65a, 16'hb65b, 16'hb65c, 16'hb65d, 16'hb65e, 16'hb65f 	:	val_out <= 16'h0393;
         16'hb660, 16'hb661, 16'hb662, 16'hb663, 16'hb664, 16'hb665, 16'hb666, 16'hb667 	:	val_out <= 16'h038e;
         16'hb668, 16'hb669, 16'hb66a, 16'hb66b, 16'hb66c, 16'hb66d, 16'hb66e, 16'hb66f 	:	val_out <= 16'h0388;
         16'hb670, 16'hb671, 16'hb672, 16'hb673, 16'hb674, 16'hb675, 16'hb676, 16'hb677 	:	val_out <= 16'h0382;
         16'hb678, 16'hb679, 16'hb67a, 16'hb67b, 16'hb67c, 16'hb67d, 16'hb67e, 16'hb67f 	:	val_out <= 16'h037c;
         16'hb680, 16'hb681, 16'hb682, 16'hb683, 16'hb684, 16'hb685, 16'hb686, 16'hb687 	:	val_out <= 16'h0376;
         16'hb688, 16'hb689, 16'hb68a, 16'hb68b, 16'hb68c, 16'hb68d, 16'hb68e, 16'hb68f 	:	val_out <= 16'h0370;
         16'hb690, 16'hb691, 16'hb692, 16'hb693, 16'hb694, 16'hb695, 16'hb696, 16'hb697 	:	val_out <= 16'h036b;
         16'hb698, 16'hb699, 16'hb69a, 16'hb69b, 16'hb69c, 16'hb69d, 16'hb69e, 16'hb69f 	:	val_out <= 16'h0365;
         16'hb6a0, 16'hb6a1, 16'hb6a2, 16'hb6a3, 16'hb6a4, 16'hb6a5, 16'hb6a6, 16'hb6a7 	:	val_out <= 16'h035f;
         16'hb6a8, 16'hb6a9, 16'hb6aa, 16'hb6ab, 16'hb6ac, 16'hb6ad, 16'hb6ae, 16'hb6af 	:	val_out <= 16'h0359;
         16'hb6b0, 16'hb6b1, 16'hb6b2, 16'hb6b3, 16'hb6b4, 16'hb6b5, 16'hb6b6, 16'hb6b7 	:	val_out <= 16'h0354;
         16'hb6b8, 16'hb6b9, 16'hb6ba, 16'hb6bb, 16'hb6bc, 16'hb6bd, 16'hb6be, 16'hb6bf 	:	val_out <= 16'h034e;
         16'hb6c0, 16'hb6c1, 16'hb6c2, 16'hb6c3, 16'hb6c4, 16'hb6c5, 16'hb6c6, 16'hb6c7 	:	val_out <= 16'h0348;
         16'hb6c8, 16'hb6c9, 16'hb6ca, 16'hb6cb, 16'hb6cc, 16'hb6cd, 16'hb6ce, 16'hb6cf 	:	val_out <= 16'h0343;
         16'hb6d0, 16'hb6d1, 16'hb6d2, 16'hb6d3, 16'hb6d4, 16'hb6d5, 16'hb6d6, 16'hb6d7 	:	val_out <= 16'h033d;
         16'hb6d8, 16'hb6d9, 16'hb6da, 16'hb6db, 16'hb6dc, 16'hb6dd, 16'hb6de, 16'hb6df 	:	val_out <= 16'h0337;
         16'hb6e0, 16'hb6e1, 16'hb6e2, 16'hb6e3, 16'hb6e4, 16'hb6e5, 16'hb6e6, 16'hb6e7 	:	val_out <= 16'h0332;
         16'hb6e8, 16'hb6e9, 16'hb6ea, 16'hb6eb, 16'hb6ec, 16'hb6ed, 16'hb6ee, 16'hb6ef 	:	val_out <= 16'h032c;
         16'hb6f0, 16'hb6f1, 16'hb6f2, 16'hb6f3, 16'hb6f4, 16'hb6f5, 16'hb6f6, 16'hb6f7 	:	val_out <= 16'h0327;
         16'hb6f8, 16'hb6f9, 16'hb6fa, 16'hb6fb, 16'hb6fc, 16'hb6fd, 16'hb6fe, 16'hb6ff 	:	val_out <= 16'h0321;
         16'hb700, 16'hb701, 16'hb702, 16'hb703, 16'hb704, 16'hb705, 16'hb706, 16'hb707 	:	val_out <= 16'h031c;
         16'hb708, 16'hb709, 16'hb70a, 16'hb70b, 16'hb70c, 16'hb70d, 16'hb70e, 16'hb70f 	:	val_out <= 16'h0316;
         16'hb710, 16'hb711, 16'hb712, 16'hb713, 16'hb714, 16'hb715, 16'hb716, 16'hb717 	:	val_out <= 16'h0311;
         16'hb718, 16'hb719, 16'hb71a, 16'hb71b, 16'hb71c, 16'hb71d, 16'hb71e, 16'hb71f 	:	val_out <= 16'h030b;
         16'hb720, 16'hb721, 16'hb722, 16'hb723, 16'hb724, 16'hb725, 16'hb726, 16'hb727 	:	val_out <= 16'h0306;
         16'hb728, 16'hb729, 16'hb72a, 16'hb72b, 16'hb72c, 16'hb72d, 16'hb72e, 16'hb72f 	:	val_out <= 16'h0300;
         16'hb730, 16'hb731, 16'hb732, 16'hb733, 16'hb734, 16'hb735, 16'hb736, 16'hb737 	:	val_out <= 16'h02fb;
         16'hb738, 16'hb739, 16'hb73a, 16'hb73b, 16'hb73c, 16'hb73d, 16'hb73e, 16'hb73f 	:	val_out <= 16'h02f6;
         16'hb740, 16'hb741, 16'hb742, 16'hb743, 16'hb744, 16'hb745, 16'hb746, 16'hb747 	:	val_out <= 16'h02f0;
         16'hb748, 16'hb749, 16'hb74a, 16'hb74b, 16'hb74c, 16'hb74d, 16'hb74e, 16'hb74f 	:	val_out <= 16'h02eb;
         16'hb750, 16'hb751, 16'hb752, 16'hb753, 16'hb754, 16'hb755, 16'hb756, 16'hb757 	:	val_out <= 16'h02e6;
         16'hb758, 16'hb759, 16'hb75a, 16'hb75b, 16'hb75c, 16'hb75d, 16'hb75e, 16'hb75f 	:	val_out <= 16'h02e0;
         16'hb760, 16'hb761, 16'hb762, 16'hb763, 16'hb764, 16'hb765, 16'hb766, 16'hb767 	:	val_out <= 16'h02db;
         16'hb768, 16'hb769, 16'hb76a, 16'hb76b, 16'hb76c, 16'hb76d, 16'hb76e, 16'hb76f 	:	val_out <= 16'h02d6;
         16'hb770, 16'hb771, 16'hb772, 16'hb773, 16'hb774, 16'hb775, 16'hb776, 16'hb777 	:	val_out <= 16'h02d0;
         16'hb778, 16'hb779, 16'hb77a, 16'hb77b, 16'hb77c, 16'hb77d, 16'hb77e, 16'hb77f 	:	val_out <= 16'h02cb;
         16'hb780, 16'hb781, 16'hb782, 16'hb783, 16'hb784, 16'hb785, 16'hb786, 16'hb787 	:	val_out <= 16'h02c6;
         16'hb788, 16'hb789, 16'hb78a, 16'hb78b, 16'hb78c, 16'hb78d, 16'hb78e, 16'hb78f 	:	val_out <= 16'h02c1;
         16'hb790, 16'hb791, 16'hb792, 16'hb793, 16'hb794, 16'hb795, 16'hb796, 16'hb797 	:	val_out <= 16'h02bc;
         16'hb798, 16'hb799, 16'hb79a, 16'hb79b, 16'hb79c, 16'hb79d, 16'hb79e, 16'hb79f 	:	val_out <= 16'h02b6;
         16'hb7a0, 16'hb7a1, 16'hb7a2, 16'hb7a3, 16'hb7a4, 16'hb7a5, 16'hb7a6, 16'hb7a7 	:	val_out <= 16'h02b1;
         16'hb7a8, 16'hb7a9, 16'hb7aa, 16'hb7ab, 16'hb7ac, 16'hb7ad, 16'hb7ae, 16'hb7af 	:	val_out <= 16'h02ac;
         16'hb7b0, 16'hb7b1, 16'hb7b2, 16'hb7b3, 16'hb7b4, 16'hb7b5, 16'hb7b6, 16'hb7b7 	:	val_out <= 16'h02a7;
         16'hb7b8, 16'hb7b9, 16'hb7ba, 16'hb7bb, 16'hb7bc, 16'hb7bd, 16'hb7be, 16'hb7bf 	:	val_out <= 16'h02a2;
         16'hb7c0, 16'hb7c1, 16'hb7c2, 16'hb7c3, 16'hb7c4, 16'hb7c5, 16'hb7c6, 16'hb7c7 	:	val_out <= 16'h029d;
         16'hb7c8, 16'hb7c9, 16'hb7ca, 16'hb7cb, 16'hb7cc, 16'hb7cd, 16'hb7ce, 16'hb7cf 	:	val_out <= 16'h0298;
         16'hb7d0, 16'hb7d1, 16'hb7d2, 16'hb7d3, 16'hb7d4, 16'hb7d5, 16'hb7d6, 16'hb7d7 	:	val_out <= 16'h0293;
         16'hb7d8, 16'hb7d9, 16'hb7da, 16'hb7db, 16'hb7dc, 16'hb7dd, 16'hb7de, 16'hb7df 	:	val_out <= 16'h028e;
         16'hb7e0, 16'hb7e1, 16'hb7e2, 16'hb7e3, 16'hb7e4, 16'hb7e5, 16'hb7e6, 16'hb7e7 	:	val_out <= 16'h0289;
         16'hb7e8, 16'hb7e9, 16'hb7ea, 16'hb7eb, 16'hb7ec, 16'hb7ed, 16'hb7ee, 16'hb7ef 	:	val_out <= 16'h0284;
         16'hb7f0, 16'hb7f1, 16'hb7f2, 16'hb7f3, 16'hb7f4, 16'hb7f5, 16'hb7f6, 16'hb7f7 	:	val_out <= 16'h027f;
         16'hb7f8, 16'hb7f9, 16'hb7fa, 16'hb7fb, 16'hb7fc, 16'hb7fd, 16'hb7fe, 16'hb7ff 	:	val_out <= 16'h027a;
         16'hb800, 16'hb801, 16'hb802, 16'hb803, 16'hb804, 16'hb805, 16'hb806, 16'hb807 	:	val_out <= 16'h0275;
         16'hb808, 16'hb809, 16'hb80a, 16'hb80b, 16'hb80c, 16'hb80d, 16'hb80e, 16'hb80f 	:	val_out <= 16'h0270;
         16'hb810, 16'hb811, 16'hb812, 16'hb813, 16'hb814, 16'hb815, 16'hb816, 16'hb817 	:	val_out <= 16'h026b;
         16'hb818, 16'hb819, 16'hb81a, 16'hb81b, 16'hb81c, 16'hb81d, 16'hb81e, 16'hb81f 	:	val_out <= 16'h0267;
         16'hb820, 16'hb821, 16'hb822, 16'hb823, 16'hb824, 16'hb825, 16'hb826, 16'hb827 	:	val_out <= 16'h0262;
         16'hb828, 16'hb829, 16'hb82a, 16'hb82b, 16'hb82c, 16'hb82d, 16'hb82e, 16'hb82f 	:	val_out <= 16'h025d;
         16'hb830, 16'hb831, 16'hb832, 16'hb833, 16'hb834, 16'hb835, 16'hb836, 16'hb837 	:	val_out <= 16'h0258;
         16'hb838, 16'hb839, 16'hb83a, 16'hb83b, 16'hb83c, 16'hb83d, 16'hb83e, 16'hb83f 	:	val_out <= 16'h0253;
         16'hb840, 16'hb841, 16'hb842, 16'hb843, 16'hb844, 16'hb845, 16'hb846, 16'hb847 	:	val_out <= 16'h024f;
         16'hb848, 16'hb849, 16'hb84a, 16'hb84b, 16'hb84c, 16'hb84d, 16'hb84e, 16'hb84f 	:	val_out <= 16'h024a;
         16'hb850, 16'hb851, 16'hb852, 16'hb853, 16'hb854, 16'hb855, 16'hb856, 16'hb857 	:	val_out <= 16'h0245;
         16'hb858, 16'hb859, 16'hb85a, 16'hb85b, 16'hb85c, 16'hb85d, 16'hb85e, 16'hb85f 	:	val_out <= 16'h0240;
         16'hb860, 16'hb861, 16'hb862, 16'hb863, 16'hb864, 16'hb865, 16'hb866, 16'hb867 	:	val_out <= 16'h023c;
         16'hb868, 16'hb869, 16'hb86a, 16'hb86b, 16'hb86c, 16'hb86d, 16'hb86e, 16'hb86f 	:	val_out <= 16'h0237;
         16'hb870, 16'hb871, 16'hb872, 16'hb873, 16'hb874, 16'hb875, 16'hb876, 16'hb877 	:	val_out <= 16'h0232;
         16'hb878, 16'hb879, 16'hb87a, 16'hb87b, 16'hb87c, 16'hb87d, 16'hb87e, 16'hb87f 	:	val_out <= 16'h022e;
         16'hb880, 16'hb881, 16'hb882, 16'hb883, 16'hb884, 16'hb885, 16'hb886, 16'hb887 	:	val_out <= 16'h0229;
         16'hb888, 16'hb889, 16'hb88a, 16'hb88b, 16'hb88c, 16'hb88d, 16'hb88e, 16'hb88f 	:	val_out <= 16'h0225;
         16'hb890, 16'hb891, 16'hb892, 16'hb893, 16'hb894, 16'hb895, 16'hb896, 16'hb897 	:	val_out <= 16'h0220;
         16'hb898, 16'hb899, 16'hb89a, 16'hb89b, 16'hb89c, 16'hb89d, 16'hb89e, 16'hb89f 	:	val_out <= 16'h021b;
         16'hb8a0, 16'hb8a1, 16'hb8a2, 16'hb8a3, 16'hb8a4, 16'hb8a5, 16'hb8a6, 16'hb8a7 	:	val_out <= 16'h0217;
         16'hb8a8, 16'hb8a9, 16'hb8aa, 16'hb8ab, 16'hb8ac, 16'hb8ad, 16'hb8ae, 16'hb8af 	:	val_out <= 16'h0212;
         16'hb8b0, 16'hb8b1, 16'hb8b2, 16'hb8b3, 16'hb8b4, 16'hb8b5, 16'hb8b6, 16'hb8b7 	:	val_out <= 16'h020e;
         16'hb8b8, 16'hb8b9, 16'hb8ba, 16'hb8bb, 16'hb8bc, 16'hb8bd, 16'hb8be, 16'hb8bf 	:	val_out <= 16'h0209;
         16'hb8c0, 16'hb8c1, 16'hb8c2, 16'hb8c3, 16'hb8c4, 16'hb8c5, 16'hb8c6, 16'hb8c7 	:	val_out <= 16'h0205;
         16'hb8c8, 16'hb8c9, 16'hb8ca, 16'hb8cb, 16'hb8cc, 16'hb8cd, 16'hb8ce, 16'hb8cf 	:	val_out <= 16'h0200;
         16'hb8d0, 16'hb8d1, 16'hb8d2, 16'hb8d3, 16'hb8d4, 16'hb8d5, 16'hb8d6, 16'hb8d7 	:	val_out <= 16'h01fc;
         16'hb8d8, 16'hb8d9, 16'hb8da, 16'hb8db, 16'hb8dc, 16'hb8dd, 16'hb8de, 16'hb8df 	:	val_out <= 16'h01f8;
         16'hb8e0, 16'hb8e1, 16'hb8e2, 16'hb8e3, 16'hb8e4, 16'hb8e5, 16'hb8e6, 16'hb8e7 	:	val_out <= 16'h01f3;
         16'hb8e8, 16'hb8e9, 16'hb8ea, 16'hb8eb, 16'hb8ec, 16'hb8ed, 16'hb8ee, 16'hb8ef 	:	val_out <= 16'h01ef;
         16'hb8f0, 16'hb8f1, 16'hb8f2, 16'hb8f3, 16'hb8f4, 16'hb8f5, 16'hb8f6, 16'hb8f7 	:	val_out <= 16'h01eb;
         16'hb8f8, 16'hb8f9, 16'hb8fa, 16'hb8fb, 16'hb8fc, 16'hb8fd, 16'hb8fe, 16'hb8ff 	:	val_out <= 16'h01e6;
         16'hb900, 16'hb901, 16'hb902, 16'hb903, 16'hb904, 16'hb905, 16'hb906, 16'hb907 	:	val_out <= 16'h01e2;
         16'hb908, 16'hb909, 16'hb90a, 16'hb90b, 16'hb90c, 16'hb90d, 16'hb90e, 16'hb90f 	:	val_out <= 16'h01de;
         16'hb910, 16'hb911, 16'hb912, 16'hb913, 16'hb914, 16'hb915, 16'hb916, 16'hb917 	:	val_out <= 16'h01d9;
         16'hb918, 16'hb919, 16'hb91a, 16'hb91b, 16'hb91c, 16'hb91d, 16'hb91e, 16'hb91f 	:	val_out <= 16'h01d5;
         16'hb920, 16'hb921, 16'hb922, 16'hb923, 16'hb924, 16'hb925, 16'hb926, 16'hb927 	:	val_out <= 16'h01d1;
         16'hb928, 16'hb929, 16'hb92a, 16'hb92b, 16'hb92c, 16'hb92d, 16'hb92e, 16'hb92f 	:	val_out <= 16'h01cd;
         16'hb930, 16'hb931, 16'hb932, 16'hb933, 16'hb934, 16'hb935, 16'hb936, 16'hb937 	:	val_out <= 16'h01c8;
         16'hb938, 16'hb939, 16'hb93a, 16'hb93b, 16'hb93c, 16'hb93d, 16'hb93e, 16'hb93f 	:	val_out <= 16'h01c4;
         16'hb940, 16'hb941, 16'hb942, 16'hb943, 16'hb944, 16'hb945, 16'hb946, 16'hb947 	:	val_out <= 16'h01c0;
         16'hb948, 16'hb949, 16'hb94a, 16'hb94b, 16'hb94c, 16'hb94d, 16'hb94e, 16'hb94f 	:	val_out <= 16'h01bc;
         16'hb950, 16'hb951, 16'hb952, 16'hb953, 16'hb954, 16'hb955, 16'hb956, 16'hb957 	:	val_out <= 16'h01b8;
         16'hb958, 16'hb959, 16'hb95a, 16'hb95b, 16'hb95c, 16'hb95d, 16'hb95e, 16'hb95f 	:	val_out <= 16'h01b4;
         16'hb960, 16'hb961, 16'hb962, 16'hb963, 16'hb964, 16'hb965, 16'hb966, 16'hb967 	:	val_out <= 16'h01b0;
         16'hb968, 16'hb969, 16'hb96a, 16'hb96b, 16'hb96c, 16'hb96d, 16'hb96e, 16'hb96f 	:	val_out <= 16'h01ac;
         16'hb970, 16'hb971, 16'hb972, 16'hb973, 16'hb974, 16'hb975, 16'hb976, 16'hb977 	:	val_out <= 16'h01a8;
         16'hb978, 16'hb979, 16'hb97a, 16'hb97b, 16'hb97c, 16'hb97d, 16'hb97e, 16'hb97f 	:	val_out <= 16'h01a4;
         16'hb980, 16'hb981, 16'hb982, 16'hb983, 16'hb984, 16'hb985, 16'hb986, 16'hb987 	:	val_out <= 16'h01a0;
         16'hb988, 16'hb989, 16'hb98a, 16'hb98b, 16'hb98c, 16'hb98d, 16'hb98e, 16'hb98f 	:	val_out <= 16'h019c;
         16'hb990, 16'hb991, 16'hb992, 16'hb993, 16'hb994, 16'hb995, 16'hb996, 16'hb997 	:	val_out <= 16'h0198;
         16'hb998, 16'hb999, 16'hb99a, 16'hb99b, 16'hb99c, 16'hb99d, 16'hb99e, 16'hb99f 	:	val_out <= 16'h0194;
         16'hb9a0, 16'hb9a1, 16'hb9a2, 16'hb9a3, 16'hb9a4, 16'hb9a5, 16'hb9a6, 16'hb9a7 	:	val_out <= 16'h0190;
         16'hb9a8, 16'hb9a9, 16'hb9aa, 16'hb9ab, 16'hb9ac, 16'hb9ad, 16'hb9ae, 16'hb9af 	:	val_out <= 16'h018c;
         16'hb9b0, 16'hb9b1, 16'hb9b2, 16'hb9b3, 16'hb9b4, 16'hb9b5, 16'hb9b6, 16'hb9b7 	:	val_out <= 16'h0188;
         16'hb9b8, 16'hb9b9, 16'hb9ba, 16'hb9bb, 16'hb9bc, 16'hb9bd, 16'hb9be, 16'hb9bf 	:	val_out <= 16'h0184;
         16'hb9c0, 16'hb9c1, 16'hb9c2, 16'hb9c3, 16'hb9c4, 16'hb9c5, 16'hb9c6, 16'hb9c7 	:	val_out <= 16'h0180;
         16'hb9c8, 16'hb9c9, 16'hb9ca, 16'hb9cb, 16'hb9cc, 16'hb9cd, 16'hb9ce, 16'hb9cf 	:	val_out <= 16'h017c;
         16'hb9d0, 16'hb9d1, 16'hb9d2, 16'hb9d3, 16'hb9d4, 16'hb9d5, 16'hb9d6, 16'hb9d7 	:	val_out <= 16'h0179;
         16'hb9d8, 16'hb9d9, 16'hb9da, 16'hb9db, 16'hb9dc, 16'hb9dd, 16'hb9de, 16'hb9df 	:	val_out <= 16'h0175;
         16'hb9e0, 16'hb9e1, 16'hb9e2, 16'hb9e3, 16'hb9e4, 16'hb9e5, 16'hb9e6, 16'hb9e7 	:	val_out <= 16'h0171;
         16'hb9e8, 16'hb9e9, 16'hb9ea, 16'hb9eb, 16'hb9ec, 16'hb9ed, 16'hb9ee, 16'hb9ef 	:	val_out <= 16'h016d;
         16'hb9f0, 16'hb9f1, 16'hb9f2, 16'hb9f3, 16'hb9f4, 16'hb9f5, 16'hb9f6, 16'hb9f7 	:	val_out <= 16'h016a;
         16'hb9f8, 16'hb9f9, 16'hb9fa, 16'hb9fb, 16'hb9fc, 16'hb9fd, 16'hb9fe, 16'hb9ff 	:	val_out <= 16'h0166;
         16'hba00, 16'hba01, 16'hba02, 16'hba03, 16'hba04, 16'hba05, 16'hba06, 16'hba07 	:	val_out <= 16'h0162;
         16'hba08, 16'hba09, 16'hba0a, 16'hba0b, 16'hba0c, 16'hba0d, 16'hba0e, 16'hba0f 	:	val_out <= 16'h015e;
         16'hba10, 16'hba11, 16'hba12, 16'hba13, 16'hba14, 16'hba15, 16'hba16, 16'hba17 	:	val_out <= 16'h015b;
         16'hba18, 16'hba19, 16'hba1a, 16'hba1b, 16'hba1c, 16'hba1d, 16'hba1e, 16'hba1f 	:	val_out <= 16'h0157;
         16'hba20, 16'hba21, 16'hba22, 16'hba23, 16'hba24, 16'hba25, 16'hba26, 16'hba27 	:	val_out <= 16'h0154;
         16'hba28, 16'hba29, 16'hba2a, 16'hba2b, 16'hba2c, 16'hba2d, 16'hba2e, 16'hba2f 	:	val_out <= 16'h0150;
         16'hba30, 16'hba31, 16'hba32, 16'hba33, 16'hba34, 16'hba35, 16'hba36, 16'hba37 	:	val_out <= 16'h014c;
         16'hba38, 16'hba39, 16'hba3a, 16'hba3b, 16'hba3c, 16'hba3d, 16'hba3e, 16'hba3f 	:	val_out <= 16'h0149;
         16'hba40, 16'hba41, 16'hba42, 16'hba43, 16'hba44, 16'hba45, 16'hba46, 16'hba47 	:	val_out <= 16'h0145;
         16'hba48, 16'hba49, 16'hba4a, 16'hba4b, 16'hba4c, 16'hba4d, 16'hba4e, 16'hba4f 	:	val_out <= 16'h0142;
         16'hba50, 16'hba51, 16'hba52, 16'hba53, 16'hba54, 16'hba55, 16'hba56, 16'hba57 	:	val_out <= 16'h013e;
         16'hba58, 16'hba59, 16'hba5a, 16'hba5b, 16'hba5c, 16'hba5d, 16'hba5e, 16'hba5f 	:	val_out <= 16'h013b;
         16'hba60, 16'hba61, 16'hba62, 16'hba63, 16'hba64, 16'hba65, 16'hba66, 16'hba67 	:	val_out <= 16'h0137;
         16'hba68, 16'hba69, 16'hba6a, 16'hba6b, 16'hba6c, 16'hba6d, 16'hba6e, 16'hba6f 	:	val_out <= 16'h0134;
         16'hba70, 16'hba71, 16'hba72, 16'hba73, 16'hba74, 16'hba75, 16'hba76, 16'hba77 	:	val_out <= 16'h0130;
         16'hba78, 16'hba79, 16'hba7a, 16'hba7b, 16'hba7c, 16'hba7d, 16'hba7e, 16'hba7f 	:	val_out <= 16'h012d;
         16'hba80, 16'hba81, 16'hba82, 16'hba83, 16'hba84, 16'hba85, 16'hba86, 16'hba87 	:	val_out <= 16'h012a;
         16'hba88, 16'hba89, 16'hba8a, 16'hba8b, 16'hba8c, 16'hba8d, 16'hba8e, 16'hba8f 	:	val_out <= 16'h0126;
         16'hba90, 16'hba91, 16'hba92, 16'hba93, 16'hba94, 16'hba95, 16'hba96, 16'hba97 	:	val_out <= 16'h0123;
         16'hba98, 16'hba99, 16'hba9a, 16'hba9b, 16'hba9c, 16'hba9d, 16'hba9e, 16'hba9f 	:	val_out <= 16'h0120;
         16'hbaa0, 16'hbaa1, 16'hbaa2, 16'hbaa3, 16'hbaa4, 16'hbaa5, 16'hbaa6, 16'hbaa7 	:	val_out <= 16'h011c;
         16'hbaa8, 16'hbaa9, 16'hbaaa, 16'hbaab, 16'hbaac, 16'hbaad, 16'hbaae, 16'hbaaf 	:	val_out <= 16'h0119;
         16'hbab0, 16'hbab1, 16'hbab2, 16'hbab3, 16'hbab4, 16'hbab5, 16'hbab6, 16'hbab7 	:	val_out <= 16'h0116;
         16'hbab8, 16'hbab9, 16'hbaba, 16'hbabb, 16'hbabc, 16'hbabd, 16'hbabe, 16'hbabf 	:	val_out <= 16'h0112;
         16'hbac0, 16'hbac1, 16'hbac2, 16'hbac3, 16'hbac4, 16'hbac5, 16'hbac6, 16'hbac7 	:	val_out <= 16'h010f;
         16'hbac8, 16'hbac9, 16'hbaca, 16'hbacb, 16'hbacc, 16'hbacd, 16'hbace, 16'hbacf 	:	val_out <= 16'h010c;
         16'hbad0, 16'hbad1, 16'hbad2, 16'hbad3, 16'hbad4, 16'hbad5, 16'hbad6, 16'hbad7 	:	val_out <= 16'h0109;
         16'hbad8, 16'hbad9, 16'hbada, 16'hbadb, 16'hbadc, 16'hbadd, 16'hbade, 16'hbadf 	:	val_out <= 16'h0106;
         16'hbae0, 16'hbae1, 16'hbae2, 16'hbae3, 16'hbae4, 16'hbae5, 16'hbae6, 16'hbae7 	:	val_out <= 16'h0102;
         16'hbae8, 16'hbae9, 16'hbaea, 16'hbaeb, 16'hbaec, 16'hbaed, 16'hbaee, 16'hbaef 	:	val_out <= 16'h00ff;
         16'hbaf0, 16'hbaf1, 16'hbaf2, 16'hbaf3, 16'hbaf4, 16'hbaf5, 16'hbaf6, 16'hbaf7 	:	val_out <= 16'h00fc;
         16'hbaf8, 16'hbaf9, 16'hbafa, 16'hbafb, 16'hbafc, 16'hbafd, 16'hbafe, 16'hbaff 	:	val_out <= 16'h00f9;
         16'hbb00, 16'hbb01, 16'hbb02, 16'hbb03, 16'hbb04, 16'hbb05, 16'hbb06, 16'hbb07 	:	val_out <= 16'h00f6;
         16'hbb08, 16'hbb09, 16'hbb0a, 16'hbb0b, 16'hbb0c, 16'hbb0d, 16'hbb0e, 16'hbb0f 	:	val_out <= 16'h00f3;
         16'hbb10, 16'hbb11, 16'hbb12, 16'hbb13, 16'hbb14, 16'hbb15, 16'hbb16, 16'hbb17 	:	val_out <= 16'h00f0;
         16'hbb18, 16'hbb19, 16'hbb1a, 16'hbb1b, 16'hbb1c, 16'hbb1d, 16'hbb1e, 16'hbb1f 	:	val_out <= 16'h00ed;
         16'hbb20, 16'hbb21, 16'hbb22, 16'hbb23, 16'hbb24, 16'hbb25, 16'hbb26, 16'hbb27 	:	val_out <= 16'h00ea;
         16'hbb28, 16'hbb29, 16'hbb2a, 16'hbb2b, 16'hbb2c, 16'hbb2d, 16'hbb2e, 16'hbb2f 	:	val_out <= 16'h00e7;
         16'hbb30, 16'hbb31, 16'hbb32, 16'hbb33, 16'hbb34, 16'hbb35, 16'hbb36, 16'hbb37 	:	val_out <= 16'h00e4;
         16'hbb38, 16'hbb39, 16'hbb3a, 16'hbb3b, 16'hbb3c, 16'hbb3d, 16'hbb3e, 16'hbb3f 	:	val_out <= 16'h00e1;
         16'hbb40, 16'hbb41, 16'hbb42, 16'hbb43, 16'hbb44, 16'hbb45, 16'hbb46, 16'hbb47 	:	val_out <= 16'h00de;
         16'hbb48, 16'hbb49, 16'hbb4a, 16'hbb4b, 16'hbb4c, 16'hbb4d, 16'hbb4e, 16'hbb4f 	:	val_out <= 16'h00db;
         16'hbb50, 16'hbb51, 16'hbb52, 16'hbb53, 16'hbb54, 16'hbb55, 16'hbb56, 16'hbb57 	:	val_out <= 16'h00d8;
         16'hbb58, 16'hbb59, 16'hbb5a, 16'hbb5b, 16'hbb5c, 16'hbb5d, 16'hbb5e, 16'hbb5f 	:	val_out <= 16'h00d5;
         16'hbb60, 16'hbb61, 16'hbb62, 16'hbb63, 16'hbb64, 16'hbb65, 16'hbb66, 16'hbb67 	:	val_out <= 16'h00d2;
         16'hbb68, 16'hbb69, 16'hbb6a, 16'hbb6b, 16'hbb6c, 16'hbb6d, 16'hbb6e, 16'hbb6f 	:	val_out <= 16'h00d0;
         16'hbb70, 16'hbb71, 16'hbb72, 16'hbb73, 16'hbb74, 16'hbb75, 16'hbb76, 16'hbb77 	:	val_out <= 16'h00cd;
         16'hbb78, 16'hbb79, 16'hbb7a, 16'hbb7b, 16'hbb7c, 16'hbb7d, 16'hbb7e, 16'hbb7f 	:	val_out <= 16'h00ca;
         16'hbb80, 16'hbb81, 16'hbb82, 16'hbb83, 16'hbb84, 16'hbb85, 16'hbb86, 16'hbb87 	:	val_out <= 16'h00c7;
         16'hbb88, 16'hbb89, 16'hbb8a, 16'hbb8b, 16'hbb8c, 16'hbb8d, 16'hbb8e, 16'hbb8f 	:	val_out <= 16'h00c4;
         16'hbb90, 16'hbb91, 16'hbb92, 16'hbb93, 16'hbb94, 16'hbb95, 16'hbb96, 16'hbb97 	:	val_out <= 16'h00c2;
         16'hbb98, 16'hbb99, 16'hbb9a, 16'hbb9b, 16'hbb9c, 16'hbb9d, 16'hbb9e, 16'hbb9f 	:	val_out <= 16'h00bf;
         16'hbba0, 16'hbba1, 16'hbba2, 16'hbba3, 16'hbba4, 16'hbba5, 16'hbba6, 16'hbba7 	:	val_out <= 16'h00bc;
         16'hbba8, 16'hbba9, 16'hbbaa, 16'hbbab, 16'hbbac, 16'hbbad, 16'hbbae, 16'hbbaf 	:	val_out <= 16'h00ba;
         16'hbbb0, 16'hbbb1, 16'hbbb2, 16'hbbb3, 16'hbbb4, 16'hbbb5, 16'hbbb6, 16'hbbb7 	:	val_out <= 16'h00b7;
         16'hbbb8, 16'hbbb9, 16'hbbba, 16'hbbbb, 16'hbbbc, 16'hbbbd, 16'hbbbe, 16'hbbbf 	:	val_out <= 16'h00b4;
         16'hbbc0, 16'hbbc1, 16'hbbc2, 16'hbbc3, 16'hbbc4, 16'hbbc5, 16'hbbc6, 16'hbbc7 	:	val_out <= 16'h00b2;
         16'hbbc8, 16'hbbc9, 16'hbbca, 16'hbbcb, 16'hbbcc, 16'hbbcd, 16'hbbce, 16'hbbcf 	:	val_out <= 16'h00af;
         16'hbbd0, 16'hbbd1, 16'hbbd2, 16'hbbd3, 16'hbbd4, 16'hbbd5, 16'hbbd6, 16'hbbd7 	:	val_out <= 16'h00ac;
         16'hbbd8, 16'hbbd9, 16'hbbda, 16'hbbdb, 16'hbbdc, 16'hbbdd, 16'hbbde, 16'hbbdf 	:	val_out <= 16'h00aa;
         16'hbbe0, 16'hbbe1, 16'hbbe2, 16'hbbe3, 16'hbbe4, 16'hbbe5, 16'hbbe6, 16'hbbe7 	:	val_out <= 16'h00a7;
         16'hbbe8, 16'hbbe9, 16'hbbea, 16'hbbeb, 16'hbbec, 16'hbbed, 16'hbbee, 16'hbbef 	:	val_out <= 16'h00a5;
         16'hbbf0, 16'hbbf1, 16'hbbf2, 16'hbbf3, 16'hbbf4, 16'hbbf5, 16'hbbf6, 16'hbbf7 	:	val_out <= 16'h00a2;
         16'hbbf8, 16'hbbf9, 16'hbbfa, 16'hbbfb, 16'hbbfc, 16'hbbfd, 16'hbbfe, 16'hbbff 	:	val_out <= 16'h00a0;
         16'hbc00, 16'hbc01, 16'hbc02, 16'hbc03, 16'hbc04, 16'hbc05, 16'hbc06, 16'hbc07 	:	val_out <= 16'h009d;
         16'hbc08, 16'hbc09, 16'hbc0a, 16'hbc0b, 16'hbc0c, 16'hbc0d, 16'hbc0e, 16'hbc0f 	:	val_out <= 16'h009b;
         16'hbc10, 16'hbc11, 16'hbc12, 16'hbc13, 16'hbc14, 16'hbc15, 16'hbc16, 16'hbc17 	:	val_out <= 16'h0098;
         16'hbc18, 16'hbc19, 16'hbc1a, 16'hbc1b, 16'hbc1c, 16'hbc1d, 16'hbc1e, 16'hbc1f 	:	val_out <= 16'h0096;
         16'hbc20, 16'hbc21, 16'hbc22, 16'hbc23, 16'hbc24, 16'hbc25, 16'hbc26, 16'hbc27 	:	val_out <= 16'h0094;
         16'hbc28, 16'hbc29, 16'hbc2a, 16'hbc2b, 16'hbc2c, 16'hbc2d, 16'hbc2e, 16'hbc2f 	:	val_out <= 16'h0091;
         16'hbc30, 16'hbc31, 16'hbc32, 16'hbc33, 16'hbc34, 16'hbc35, 16'hbc36, 16'hbc37 	:	val_out <= 16'h008f;
         16'hbc38, 16'hbc39, 16'hbc3a, 16'hbc3b, 16'hbc3c, 16'hbc3d, 16'hbc3e, 16'hbc3f 	:	val_out <= 16'h008d;
         16'hbc40, 16'hbc41, 16'hbc42, 16'hbc43, 16'hbc44, 16'hbc45, 16'hbc46, 16'hbc47 	:	val_out <= 16'h008a;
         16'hbc48, 16'hbc49, 16'hbc4a, 16'hbc4b, 16'hbc4c, 16'hbc4d, 16'hbc4e, 16'hbc4f 	:	val_out <= 16'h0088;
         16'hbc50, 16'hbc51, 16'hbc52, 16'hbc53, 16'hbc54, 16'hbc55, 16'hbc56, 16'hbc57 	:	val_out <= 16'h0086;
         16'hbc58, 16'hbc59, 16'hbc5a, 16'hbc5b, 16'hbc5c, 16'hbc5d, 16'hbc5e, 16'hbc5f 	:	val_out <= 16'h0083;
         16'hbc60, 16'hbc61, 16'hbc62, 16'hbc63, 16'hbc64, 16'hbc65, 16'hbc66, 16'hbc67 	:	val_out <= 16'h0081;
         16'hbc68, 16'hbc69, 16'hbc6a, 16'hbc6b, 16'hbc6c, 16'hbc6d, 16'hbc6e, 16'hbc6f 	:	val_out <= 16'h007f;
         16'hbc70, 16'hbc71, 16'hbc72, 16'hbc73, 16'hbc74, 16'hbc75, 16'hbc76, 16'hbc77 	:	val_out <= 16'h007d;
         16'hbc78, 16'hbc79, 16'hbc7a, 16'hbc7b, 16'hbc7c, 16'hbc7d, 16'hbc7e, 16'hbc7f 	:	val_out <= 16'h007a;
         16'hbc80, 16'hbc81, 16'hbc82, 16'hbc83, 16'hbc84, 16'hbc85, 16'hbc86, 16'hbc87 	:	val_out <= 16'h0078;
         16'hbc88, 16'hbc89, 16'hbc8a, 16'hbc8b, 16'hbc8c, 16'hbc8d, 16'hbc8e, 16'hbc8f 	:	val_out <= 16'h0076;
         16'hbc90, 16'hbc91, 16'hbc92, 16'hbc93, 16'hbc94, 16'hbc95, 16'hbc96, 16'hbc97 	:	val_out <= 16'h0074;
         16'hbc98, 16'hbc99, 16'hbc9a, 16'hbc9b, 16'hbc9c, 16'hbc9d, 16'hbc9e, 16'hbc9f 	:	val_out <= 16'h0072;
         16'hbca0, 16'hbca1, 16'hbca2, 16'hbca3, 16'hbca4, 16'hbca5, 16'hbca6, 16'hbca7 	:	val_out <= 16'h0070;
         16'hbca8, 16'hbca9, 16'hbcaa, 16'hbcab, 16'hbcac, 16'hbcad, 16'hbcae, 16'hbcaf 	:	val_out <= 16'h006e;
         16'hbcb0, 16'hbcb1, 16'hbcb2, 16'hbcb3, 16'hbcb4, 16'hbcb5, 16'hbcb6, 16'hbcb7 	:	val_out <= 16'h006c;
         16'hbcb8, 16'hbcb9, 16'hbcba, 16'hbcbb, 16'hbcbc, 16'hbcbd, 16'hbcbe, 16'hbcbf 	:	val_out <= 16'h006a;
         16'hbcc0, 16'hbcc1, 16'hbcc2, 16'hbcc3, 16'hbcc4, 16'hbcc5, 16'hbcc6, 16'hbcc7 	:	val_out <= 16'h0068;
         16'hbcc8, 16'hbcc9, 16'hbcca, 16'hbccb, 16'hbccc, 16'hbccd, 16'hbcce, 16'hbccf 	:	val_out <= 16'h0066;
         16'hbcd0, 16'hbcd1, 16'hbcd2, 16'hbcd3, 16'hbcd4, 16'hbcd5, 16'hbcd6, 16'hbcd7 	:	val_out <= 16'h0064;
         16'hbcd8, 16'hbcd9, 16'hbcda, 16'hbcdb, 16'hbcdc, 16'hbcdd, 16'hbcde, 16'hbcdf 	:	val_out <= 16'h0062;
         16'hbce0, 16'hbce1, 16'hbce2, 16'hbce3, 16'hbce4, 16'hbce5, 16'hbce6, 16'hbce7 	:	val_out <= 16'h0060;
         16'hbce8, 16'hbce9, 16'hbcea, 16'hbceb, 16'hbcec, 16'hbced, 16'hbcee, 16'hbcef 	:	val_out <= 16'h005e;
         16'hbcf0, 16'hbcf1, 16'hbcf2, 16'hbcf3, 16'hbcf4, 16'hbcf5, 16'hbcf6, 16'hbcf7 	:	val_out <= 16'h005c;
         16'hbcf8, 16'hbcf9, 16'hbcfa, 16'hbcfb, 16'hbcfc, 16'hbcfd, 16'hbcfe, 16'hbcff 	:	val_out <= 16'h005a;
         16'hbd00, 16'hbd01, 16'hbd02, 16'hbd03, 16'hbd04, 16'hbd05, 16'hbd06, 16'hbd07 	:	val_out <= 16'h0058;
         16'hbd08, 16'hbd09, 16'hbd0a, 16'hbd0b, 16'hbd0c, 16'hbd0d, 16'hbd0e, 16'hbd0f 	:	val_out <= 16'h0056;
         16'hbd10, 16'hbd11, 16'hbd12, 16'hbd13, 16'hbd14, 16'hbd15, 16'hbd16, 16'hbd17 	:	val_out <= 16'h0055;
         16'hbd18, 16'hbd19, 16'hbd1a, 16'hbd1b, 16'hbd1c, 16'hbd1d, 16'hbd1e, 16'hbd1f 	:	val_out <= 16'h0053;
         16'hbd20, 16'hbd21, 16'hbd22, 16'hbd23, 16'hbd24, 16'hbd25, 16'hbd26, 16'hbd27 	:	val_out <= 16'h0051;
         16'hbd28, 16'hbd29, 16'hbd2a, 16'hbd2b, 16'hbd2c, 16'hbd2d, 16'hbd2e, 16'hbd2f 	:	val_out <= 16'h004f;
         16'hbd30, 16'hbd31, 16'hbd32, 16'hbd33, 16'hbd34, 16'hbd35, 16'hbd36, 16'hbd37 	:	val_out <= 16'h004e;
         16'hbd38, 16'hbd39, 16'hbd3a, 16'hbd3b, 16'hbd3c, 16'hbd3d, 16'hbd3e, 16'hbd3f 	:	val_out <= 16'h004c;
         16'hbd40, 16'hbd41, 16'hbd42, 16'hbd43, 16'hbd44, 16'hbd45, 16'hbd46, 16'hbd47 	:	val_out <= 16'h004a;
         16'hbd48, 16'hbd49, 16'hbd4a, 16'hbd4b, 16'hbd4c, 16'hbd4d, 16'hbd4e, 16'hbd4f 	:	val_out <= 16'h0048;
         16'hbd50, 16'hbd51, 16'hbd52, 16'hbd53, 16'hbd54, 16'hbd55, 16'hbd56, 16'hbd57 	:	val_out <= 16'h0047;
         16'hbd58, 16'hbd59, 16'hbd5a, 16'hbd5b, 16'hbd5c, 16'hbd5d, 16'hbd5e, 16'hbd5f 	:	val_out <= 16'h0045;
         16'hbd60, 16'hbd61, 16'hbd62, 16'hbd63, 16'hbd64, 16'hbd65, 16'hbd66, 16'hbd67 	:	val_out <= 16'h0043;
         16'hbd68, 16'hbd69, 16'hbd6a, 16'hbd6b, 16'hbd6c, 16'hbd6d, 16'hbd6e, 16'hbd6f 	:	val_out <= 16'h0042;
         16'hbd70, 16'hbd71, 16'hbd72, 16'hbd73, 16'hbd74, 16'hbd75, 16'hbd76, 16'hbd77 	:	val_out <= 16'h0040;
         16'hbd78, 16'hbd79, 16'hbd7a, 16'hbd7b, 16'hbd7c, 16'hbd7d, 16'hbd7e, 16'hbd7f 	:	val_out <= 16'h003f;
         16'hbd80, 16'hbd81, 16'hbd82, 16'hbd83, 16'hbd84, 16'hbd85, 16'hbd86, 16'hbd87 	:	val_out <= 16'h003d;
         16'hbd88, 16'hbd89, 16'hbd8a, 16'hbd8b, 16'hbd8c, 16'hbd8d, 16'hbd8e, 16'hbd8f 	:	val_out <= 16'h003c;
         16'hbd90, 16'hbd91, 16'hbd92, 16'hbd93, 16'hbd94, 16'hbd95, 16'hbd96, 16'hbd97 	:	val_out <= 16'h003a;
         16'hbd98, 16'hbd99, 16'hbd9a, 16'hbd9b, 16'hbd9c, 16'hbd9d, 16'hbd9e, 16'hbd9f 	:	val_out <= 16'h0039;
         16'hbda0, 16'hbda1, 16'hbda2, 16'hbda3, 16'hbda4, 16'hbda5, 16'hbda6, 16'hbda7 	:	val_out <= 16'h0037;
         16'hbda8, 16'hbda9, 16'hbdaa, 16'hbdab, 16'hbdac, 16'hbdad, 16'hbdae, 16'hbdaf 	:	val_out <= 16'h0036;
         16'hbdb0, 16'hbdb1, 16'hbdb2, 16'hbdb3, 16'hbdb4, 16'hbdb5, 16'hbdb6, 16'hbdb7 	:	val_out <= 16'h0034;
         16'hbdb8, 16'hbdb9, 16'hbdba, 16'hbdbb, 16'hbdbc, 16'hbdbd, 16'hbdbe, 16'hbdbf 	:	val_out <= 16'h0033;
         16'hbdc0, 16'hbdc1, 16'hbdc2, 16'hbdc3, 16'hbdc4, 16'hbdc5, 16'hbdc6, 16'hbdc7 	:	val_out <= 16'h0031;
         16'hbdc8, 16'hbdc9, 16'hbdca, 16'hbdcb, 16'hbdcc, 16'hbdcd, 16'hbdce, 16'hbdcf 	:	val_out <= 16'h0030;
         16'hbdd0, 16'hbdd1, 16'hbdd2, 16'hbdd3, 16'hbdd4, 16'hbdd5, 16'hbdd6, 16'hbdd7 	:	val_out <= 16'h002f;
         16'hbdd8, 16'hbdd9, 16'hbdda, 16'hbddb, 16'hbddc, 16'hbddd, 16'hbdde, 16'hbddf 	:	val_out <= 16'h002d;
         16'hbde0, 16'hbde1, 16'hbde2, 16'hbde3, 16'hbde4, 16'hbde5, 16'hbde6, 16'hbde7 	:	val_out <= 16'h002c;
         16'hbde8, 16'hbde9, 16'hbdea, 16'hbdeb, 16'hbdec, 16'hbded, 16'hbdee, 16'hbdef 	:	val_out <= 16'h002b;
         16'hbdf0, 16'hbdf1, 16'hbdf2, 16'hbdf3, 16'hbdf4, 16'hbdf5, 16'hbdf6, 16'hbdf7 	:	val_out <= 16'h0029;
         16'hbdf8, 16'hbdf9, 16'hbdfa, 16'hbdfb, 16'hbdfc, 16'hbdfd, 16'hbdfe, 16'hbdff 	:	val_out <= 16'h0028;
         16'hbe00, 16'hbe01, 16'hbe02, 16'hbe03, 16'hbe04, 16'hbe05, 16'hbe06, 16'hbe07 	:	val_out <= 16'h0027;
         16'hbe08, 16'hbe09, 16'hbe0a, 16'hbe0b, 16'hbe0c, 16'hbe0d, 16'hbe0e, 16'hbe0f 	:	val_out <= 16'h0026;
         16'hbe10, 16'hbe11, 16'hbe12, 16'hbe13, 16'hbe14, 16'hbe15, 16'hbe16, 16'hbe17 	:	val_out <= 16'h0025;
         16'hbe18, 16'hbe19, 16'hbe1a, 16'hbe1b, 16'hbe1c, 16'hbe1d, 16'hbe1e, 16'hbe1f 	:	val_out <= 16'h0023;
         16'hbe20, 16'hbe21, 16'hbe22, 16'hbe23, 16'hbe24, 16'hbe25, 16'hbe26, 16'hbe27 	:	val_out <= 16'h0022;
         16'hbe28, 16'hbe29, 16'hbe2a, 16'hbe2b, 16'hbe2c, 16'hbe2d, 16'hbe2e, 16'hbe2f 	:	val_out <= 16'h0021;
         16'hbe30, 16'hbe31, 16'hbe32, 16'hbe33, 16'hbe34, 16'hbe35, 16'hbe36, 16'hbe37 	:	val_out <= 16'h0020;
         16'hbe38, 16'hbe39, 16'hbe3a, 16'hbe3b, 16'hbe3c, 16'hbe3d, 16'hbe3e, 16'hbe3f 	:	val_out <= 16'h001f;
         16'hbe40, 16'hbe41, 16'hbe42, 16'hbe43, 16'hbe44, 16'hbe45, 16'hbe46, 16'hbe47 	:	val_out <= 16'h001e;
         16'hbe48, 16'hbe49, 16'hbe4a, 16'hbe4b, 16'hbe4c, 16'hbe4d, 16'hbe4e, 16'hbe4f 	:	val_out <= 16'h001d;
         16'hbe50, 16'hbe51, 16'hbe52, 16'hbe53, 16'hbe54, 16'hbe55, 16'hbe56, 16'hbe57 	:	val_out <= 16'h001c;
         16'hbe58, 16'hbe59, 16'hbe5a, 16'hbe5b, 16'hbe5c, 16'hbe5d, 16'hbe5e, 16'hbe5f 	:	val_out <= 16'h001b;
         16'hbe60, 16'hbe61, 16'hbe62, 16'hbe63, 16'hbe64, 16'hbe65, 16'hbe66, 16'hbe67 	:	val_out <= 16'h001a;
         16'hbe68, 16'hbe69, 16'hbe6a, 16'hbe6b, 16'hbe6c, 16'hbe6d, 16'hbe6e, 16'hbe6f 	:	val_out <= 16'h0019;
         16'hbe70, 16'hbe71, 16'hbe72, 16'hbe73, 16'hbe74, 16'hbe75, 16'hbe76, 16'hbe77 	:	val_out <= 16'h0018;
         16'hbe78, 16'hbe79, 16'hbe7a, 16'hbe7b, 16'hbe7c, 16'hbe7d, 16'hbe7e, 16'hbe7f 	:	val_out <= 16'h0017;
         16'hbe80, 16'hbe81, 16'hbe82, 16'hbe83, 16'hbe84, 16'hbe85, 16'hbe86, 16'hbe87 	:	val_out <= 16'h0016;
         16'hbe88, 16'hbe89, 16'hbe8a, 16'hbe8b, 16'hbe8c, 16'hbe8d, 16'hbe8e, 16'hbe8f 	:	val_out <= 16'h0015;
         16'hbe90, 16'hbe91, 16'hbe92, 16'hbe93, 16'hbe94, 16'hbe95, 16'hbe96, 16'hbe97 	:	val_out <= 16'h0014;
         16'hbe98, 16'hbe99, 16'hbe9a, 16'hbe9b, 16'hbe9c, 16'hbe9d, 16'hbe9e, 16'hbe9f 	:	val_out <= 16'h0013;
         16'hbea0, 16'hbea1, 16'hbea2, 16'hbea3, 16'hbea4, 16'hbea5, 16'hbea6, 16'hbea7 	:	val_out <= 16'h0012;
         16'hbea8, 16'hbea9, 16'hbeaa, 16'hbeab, 16'hbeac, 16'hbead, 16'hbeae, 16'hbeaf 	:	val_out <= 16'h0011;
         16'hbeb0, 16'hbeb1, 16'hbeb2, 16'hbeb3, 16'hbeb4, 16'hbeb5, 16'hbeb6, 16'hbeb7 	:	val_out <= 16'h0011;
         16'hbeb8, 16'hbeb9, 16'hbeba, 16'hbebb, 16'hbebc, 16'hbebd, 16'hbebe, 16'hbebf 	:	val_out <= 16'h0010;
         16'hbec0, 16'hbec1, 16'hbec2, 16'hbec3, 16'hbec4, 16'hbec5, 16'hbec6, 16'hbec7 	:	val_out <= 16'h000f;
         16'hbec8, 16'hbec9, 16'hbeca, 16'hbecb, 16'hbecc, 16'hbecd, 16'hbece, 16'hbecf 	:	val_out <= 16'h000e;
         16'hbed0, 16'hbed1, 16'hbed2, 16'hbed3, 16'hbed4, 16'hbed5, 16'hbed6, 16'hbed7 	:	val_out <= 16'h000d;
         16'hbed8, 16'hbed9, 16'hbeda, 16'hbedb, 16'hbedc, 16'hbedd, 16'hbede, 16'hbedf 	:	val_out <= 16'h000d;
         16'hbee0, 16'hbee1, 16'hbee2, 16'hbee3, 16'hbee4, 16'hbee5, 16'hbee6, 16'hbee7 	:	val_out <= 16'h000c;
         16'hbee8, 16'hbee9, 16'hbeea, 16'hbeeb, 16'hbeec, 16'hbeed, 16'hbeee, 16'hbeef 	:	val_out <= 16'h000b;
         16'hbef0, 16'hbef1, 16'hbef2, 16'hbef3, 16'hbef4, 16'hbef5, 16'hbef6, 16'hbef7 	:	val_out <= 16'h000b;
         16'hbef8, 16'hbef9, 16'hbefa, 16'hbefb, 16'hbefc, 16'hbefd, 16'hbefe, 16'hbeff 	:	val_out <= 16'h000a;
         16'hbf00, 16'hbf01, 16'hbf02, 16'hbf03, 16'hbf04, 16'hbf05, 16'hbf06, 16'hbf07 	:	val_out <= 16'h0009;
         16'hbf08, 16'hbf09, 16'hbf0a, 16'hbf0b, 16'hbf0c, 16'hbf0d, 16'hbf0e, 16'hbf0f 	:	val_out <= 16'h0009;
         16'hbf10, 16'hbf11, 16'hbf12, 16'hbf13, 16'hbf14, 16'hbf15, 16'hbf16, 16'hbf17 	:	val_out <= 16'h0008;
         16'hbf18, 16'hbf19, 16'hbf1a, 16'hbf1b, 16'hbf1c, 16'hbf1d, 16'hbf1e, 16'hbf1f 	:	val_out <= 16'h0008;
         16'hbf20, 16'hbf21, 16'hbf22, 16'hbf23, 16'hbf24, 16'hbf25, 16'hbf26, 16'hbf27 	:	val_out <= 16'h0007;
         16'hbf28, 16'hbf29, 16'hbf2a, 16'hbf2b, 16'hbf2c, 16'hbf2d, 16'hbf2e, 16'hbf2f 	:	val_out <= 16'h0007;
         16'hbf30, 16'hbf31, 16'hbf32, 16'hbf33, 16'hbf34, 16'hbf35, 16'hbf36, 16'hbf37 	:	val_out <= 16'h0006;
         16'hbf38, 16'hbf39, 16'hbf3a, 16'hbf3b, 16'hbf3c, 16'hbf3d, 16'hbf3e, 16'hbf3f 	:	val_out <= 16'h0006;
         16'hbf40, 16'hbf41, 16'hbf42, 16'hbf43, 16'hbf44, 16'hbf45, 16'hbf46, 16'hbf47 	:	val_out <= 16'h0005;
         16'hbf48, 16'hbf49, 16'hbf4a, 16'hbf4b, 16'hbf4c, 16'hbf4d, 16'hbf4e, 16'hbf4f 	:	val_out <= 16'h0005;
         16'hbf50, 16'hbf51, 16'hbf52, 16'hbf53, 16'hbf54, 16'hbf55, 16'hbf56, 16'hbf57 	:	val_out <= 16'h0004;
         16'hbf58, 16'hbf59, 16'hbf5a, 16'hbf5b, 16'hbf5c, 16'hbf5d, 16'hbf5e, 16'hbf5f 	:	val_out <= 16'h0004;
         16'hbf60, 16'hbf61, 16'hbf62, 16'hbf63, 16'hbf64, 16'hbf65, 16'hbf66, 16'hbf67 	:	val_out <= 16'h0003;
         16'hbf68, 16'hbf69, 16'hbf6a, 16'hbf6b, 16'hbf6c, 16'hbf6d, 16'hbf6e, 16'hbf6f 	:	val_out <= 16'h0003;
         16'hbf70, 16'hbf71, 16'hbf72, 16'hbf73, 16'hbf74, 16'hbf75, 16'hbf76, 16'hbf77 	:	val_out <= 16'h0003;
         16'hbf78, 16'hbf79, 16'hbf7a, 16'hbf7b, 16'hbf7c, 16'hbf7d, 16'hbf7e, 16'hbf7f 	:	val_out <= 16'h0002;
         16'hbf80, 16'hbf81, 16'hbf82, 16'hbf83, 16'hbf84, 16'hbf85, 16'hbf86, 16'hbf87 	:	val_out <= 16'h0002;
         16'hbf88, 16'hbf89, 16'hbf8a, 16'hbf8b, 16'hbf8c, 16'hbf8d, 16'hbf8e, 16'hbf8f 	:	val_out <= 16'h0002;
         16'hbf90, 16'hbf91, 16'hbf92, 16'hbf93, 16'hbf94, 16'hbf95, 16'hbf96, 16'hbf97 	:	val_out <= 16'h0001;
         16'hbf98, 16'hbf99, 16'hbf9a, 16'hbf9b, 16'hbf9c, 16'hbf9d, 16'hbf9e, 16'hbf9f 	:	val_out <= 16'h0001;
         16'hbfa0, 16'hbfa1, 16'hbfa2, 16'hbfa3, 16'hbfa4, 16'hbfa5, 16'hbfa6, 16'hbfa7 	:	val_out <= 16'h0001;
         16'hbfa8, 16'hbfa9, 16'hbfaa, 16'hbfab, 16'hbfac, 16'hbfad, 16'hbfae, 16'hbfaf 	:	val_out <= 16'h0001;
         16'hbfb0, 16'hbfb1, 16'hbfb2, 16'hbfb3, 16'hbfb4, 16'hbfb5, 16'hbfb6, 16'hbfb7 	:	val_out <= 16'h0000;
         16'hbfb8, 16'hbfb9, 16'hbfba, 16'hbfbb, 16'hbfbc, 16'hbfbd, 16'hbfbe, 16'hbfbf 	:	val_out <= 16'h0000;
         16'hbfc0, 16'hbfc1, 16'hbfc2, 16'hbfc3, 16'hbfc4, 16'hbfc5, 16'hbfc6, 16'hbfc7 	:	val_out <= 16'h0000;
         16'hbfc8, 16'hbfc9, 16'hbfca, 16'hbfcb, 16'hbfcc, 16'hbfcd, 16'hbfce, 16'hbfcf 	:	val_out <= 16'h0000;
         16'hbfd0, 16'hbfd1, 16'hbfd2, 16'hbfd3, 16'hbfd4, 16'hbfd5, 16'hbfd6, 16'hbfd7 	:	val_out <= 16'h0000;
         16'hbfd8, 16'hbfd9, 16'hbfda, 16'hbfdb, 16'hbfdc, 16'hbfdd, 16'hbfde, 16'hbfdf 	:	val_out <= 16'h0000;
         16'hbfe0, 16'hbfe1, 16'hbfe2, 16'hbfe3, 16'hbfe4, 16'hbfe5, 16'hbfe6, 16'hbfe7 	:	val_out <= 16'h0000;
         16'hbfe8, 16'hbfe9, 16'hbfea, 16'hbfeb, 16'hbfec, 16'hbfed, 16'hbfee, 16'hbfef 	:	val_out <= 16'h0000;
         16'hbff0, 16'hbff1, 16'hbff2, 16'hbff3, 16'hbff4, 16'hbff5, 16'hbff6, 16'hbff7 	:	val_out <= 16'h0000;
         16'hbff8, 16'hbff9, 16'hbffa, 16'hbffb, 16'hbffc, 16'hbffd, 16'hbffe, 16'hbfff 	:	val_out <= 16'h0000;
         16'hc000, 16'hc001, 16'hc002, 16'hc003, 16'hc004, 16'hc005, 16'hc006, 16'hc007 	:	val_out <= 16'h0000;
         16'hc008, 16'hc009, 16'hc00a, 16'hc00b, 16'hc00c, 16'hc00d, 16'hc00e, 16'hc00f 	:	val_out <= 16'h0000;
         16'hc010, 16'hc011, 16'hc012, 16'hc013, 16'hc014, 16'hc015, 16'hc016, 16'hc017 	:	val_out <= 16'h0000;
         16'hc018, 16'hc019, 16'hc01a, 16'hc01b, 16'hc01c, 16'hc01d, 16'hc01e, 16'hc01f 	:	val_out <= 16'h0000;
         16'hc020, 16'hc021, 16'hc022, 16'hc023, 16'hc024, 16'hc025, 16'hc026, 16'hc027 	:	val_out <= 16'h0000;
         16'hc028, 16'hc029, 16'hc02a, 16'hc02b, 16'hc02c, 16'hc02d, 16'hc02e, 16'hc02f 	:	val_out <= 16'h0000;
         16'hc030, 16'hc031, 16'hc032, 16'hc033, 16'hc034, 16'hc035, 16'hc036, 16'hc037 	:	val_out <= 16'h0000;
         16'hc038, 16'hc039, 16'hc03a, 16'hc03b, 16'hc03c, 16'hc03d, 16'hc03e, 16'hc03f 	:	val_out <= 16'h0000;
         16'hc040, 16'hc041, 16'hc042, 16'hc043, 16'hc044, 16'hc045, 16'hc046, 16'hc047 	:	val_out <= 16'h0000;
         16'hc048, 16'hc049, 16'hc04a, 16'hc04b, 16'hc04c, 16'hc04d, 16'hc04e, 16'hc04f 	:	val_out <= 16'h0000;
         16'hc050, 16'hc051, 16'hc052, 16'hc053, 16'hc054, 16'hc055, 16'hc056, 16'hc057 	:	val_out <= 16'h0000;
         16'hc058, 16'hc059, 16'hc05a, 16'hc05b, 16'hc05c, 16'hc05d, 16'hc05e, 16'hc05f 	:	val_out <= 16'h0001;
         16'hc060, 16'hc061, 16'hc062, 16'hc063, 16'hc064, 16'hc065, 16'hc066, 16'hc067 	:	val_out <= 16'h0001;
         16'hc068, 16'hc069, 16'hc06a, 16'hc06b, 16'hc06c, 16'hc06d, 16'hc06e, 16'hc06f 	:	val_out <= 16'h0001;
         16'hc070, 16'hc071, 16'hc072, 16'hc073, 16'hc074, 16'hc075, 16'hc076, 16'hc077 	:	val_out <= 16'h0001;
         16'hc078, 16'hc079, 16'hc07a, 16'hc07b, 16'hc07c, 16'hc07d, 16'hc07e, 16'hc07f 	:	val_out <= 16'h0002;
         16'hc080, 16'hc081, 16'hc082, 16'hc083, 16'hc084, 16'hc085, 16'hc086, 16'hc087 	:	val_out <= 16'h0002;
         16'hc088, 16'hc089, 16'hc08a, 16'hc08b, 16'hc08c, 16'hc08d, 16'hc08e, 16'hc08f 	:	val_out <= 16'h0002;
         16'hc090, 16'hc091, 16'hc092, 16'hc093, 16'hc094, 16'hc095, 16'hc096, 16'hc097 	:	val_out <= 16'h0003;
         16'hc098, 16'hc099, 16'hc09a, 16'hc09b, 16'hc09c, 16'hc09d, 16'hc09e, 16'hc09f 	:	val_out <= 16'h0003;
         16'hc0a0, 16'hc0a1, 16'hc0a2, 16'hc0a3, 16'hc0a4, 16'hc0a5, 16'hc0a6, 16'hc0a7 	:	val_out <= 16'h0003;
         16'hc0a8, 16'hc0a9, 16'hc0aa, 16'hc0ab, 16'hc0ac, 16'hc0ad, 16'hc0ae, 16'hc0af 	:	val_out <= 16'h0004;
         16'hc0b0, 16'hc0b1, 16'hc0b2, 16'hc0b3, 16'hc0b4, 16'hc0b5, 16'hc0b6, 16'hc0b7 	:	val_out <= 16'h0004;
         16'hc0b8, 16'hc0b9, 16'hc0ba, 16'hc0bb, 16'hc0bc, 16'hc0bd, 16'hc0be, 16'hc0bf 	:	val_out <= 16'h0005;
         16'hc0c0, 16'hc0c1, 16'hc0c2, 16'hc0c3, 16'hc0c4, 16'hc0c5, 16'hc0c6, 16'hc0c7 	:	val_out <= 16'h0005;
         16'hc0c8, 16'hc0c9, 16'hc0ca, 16'hc0cb, 16'hc0cc, 16'hc0cd, 16'hc0ce, 16'hc0cf 	:	val_out <= 16'h0006;
         16'hc0d0, 16'hc0d1, 16'hc0d2, 16'hc0d3, 16'hc0d4, 16'hc0d5, 16'hc0d6, 16'hc0d7 	:	val_out <= 16'h0006;
         16'hc0d8, 16'hc0d9, 16'hc0da, 16'hc0db, 16'hc0dc, 16'hc0dd, 16'hc0de, 16'hc0df 	:	val_out <= 16'h0007;
         16'hc0e0, 16'hc0e1, 16'hc0e2, 16'hc0e3, 16'hc0e4, 16'hc0e5, 16'hc0e6, 16'hc0e7 	:	val_out <= 16'h0007;
         16'hc0e8, 16'hc0e9, 16'hc0ea, 16'hc0eb, 16'hc0ec, 16'hc0ed, 16'hc0ee, 16'hc0ef 	:	val_out <= 16'h0008;
         16'hc0f0, 16'hc0f1, 16'hc0f2, 16'hc0f3, 16'hc0f4, 16'hc0f5, 16'hc0f6, 16'hc0f7 	:	val_out <= 16'h0008;
         16'hc0f8, 16'hc0f9, 16'hc0fa, 16'hc0fb, 16'hc0fc, 16'hc0fd, 16'hc0fe, 16'hc0ff 	:	val_out <= 16'h0009;
         16'hc100, 16'hc101, 16'hc102, 16'hc103, 16'hc104, 16'hc105, 16'hc106, 16'hc107 	:	val_out <= 16'h0009;
         16'hc108, 16'hc109, 16'hc10a, 16'hc10b, 16'hc10c, 16'hc10d, 16'hc10e, 16'hc10f 	:	val_out <= 16'h000a;
         16'hc110, 16'hc111, 16'hc112, 16'hc113, 16'hc114, 16'hc115, 16'hc116, 16'hc117 	:	val_out <= 16'h000b;
         16'hc118, 16'hc119, 16'hc11a, 16'hc11b, 16'hc11c, 16'hc11d, 16'hc11e, 16'hc11f 	:	val_out <= 16'h000b;
         16'hc120, 16'hc121, 16'hc122, 16'hc123, 16'hc124, 16'hc125, 16'hc126, 16'hc127 	:	val_out <= 16'h000c;
         16'hc128, 16'hc129, 16'hc12a, 16'hc12b, 16'hc12c, 16'hc12d, 16'hc12e, 16'hc12f 	:	val_out <= 16'h000d;
         16'hc130, 16'hc131, 16'hc132, 16'hc133, 16'hc134, 16'hc135, 16'hc136, 16'hc137 	:	val_out <= 16'h000d;
         16'hc138, 16'hc139, 16'hc13a, 16'hc13b, 16'hc13c, 16'hc13d, 16'hc13e, 16'hc13f 	:	val_out <= 16'h000e;
         16'hc140, 16'hc141, 16'hc142, 16'hc143, 16'hc144, 16'hc145, 16'hc146, 16'hc147 	:	val_out <= 16'h000f;
         16'hc148, 16'hc149, 16'hc14a, 16'hc14b, 16'hc14c, 16'hc14d, 16'hc14e, 16'hc14f 	:	val_out <= 16'h0010;
         16'hc150, 16'hc151, 16'hc152, 16'hc153, 16'hc154, 16'hc155, 16'hc156, 16'hc157 	:	val_out <= 16'h0011;
         16'hc158, 16'hc159, 16'hc15a, 16'hc15b, 16'hc15c, 16'hc15d, 16'hc15e, 16'hc15f 	:	val_out <= 16'h0011;
         16'hc160, 16'hc161, 16'hc162, 16'hc163, 16'hc164, 16'hc165, 16'hc166, 16'hc167 	:	val_out <= 16'h0012;
         16'hc168, 16'hc169, 16'hc16a, 16'hc16b, 16'hc16c, 16'hc16d, 16'hc16e, 16'hc16f 	:	val_out <= 16'h0013;
         16'hc170, 16'hc171, 16'hc172, 16'hc173, 16'hc174, 16'hc175, 16'hc176, 16'hc177 	:	val_out <= 16'h0014;
         16'hc178, 16'hc179, 16'hc17a, 16'hc17b, 16'hc17c, 16'hc17d, 16'hc17e, 16'hc17f 	:	val_out <= 16'h0015;
         16'hc180, 16'hc181, 16'hc182, 16'hc183, 16'hc184, 16'hc185, 16'hc186, 16'hc187 	:	val_out <= 16'h0016;
         16'hc188, 16'hc189, 16'hc18a, 16'hc18b, 16'hc18c, 16'hc18d, 16'hc18e, 16'hc18f 	:	val_out <= 16'h0017;
         16'hc190, 16'hc191, 16'hc192, 16'hc193, 16'hc194, 16'hc195, 16'hc196, 16'hc197 	:	val_out <= 16'h0018;
         16'hc198, 16'hc199, 16'hc19a, 16'hc19b, 16'hc19c, 16'hc19d, 16'hc19e, 16'hc19f 	:	val_out <= 16'h0019;
         16'hc1a0, 16'hc1a1, 16'hc1a2, 16'hc1a3, 16'hc1a4, 16'hc1a5, 16'hc1a6, 16'hc1a7 	:	val_out <= 16'h001a;
         16'hc1a8, 16'hc1a9, 16'hc1aa, 16'hc1ab, 16'hc1ac, 16'hc1ad, 16'hc1ae, 16'hc1af 	:	val_out <= 16'h001b;
         16'hc1b0, 16'hc1b1, 16'hc1b2, 16'hc1b3, 16'hc1b4, 16'hc1b5, 16'hc1b6, 16'hc1b7 	:	val_out <= 16'h001c;
         16'hc1b8, 16'hc1b9, 16'hc1ba, 16'hc1bb, 16'hc1bc, 16'hc1bd, 16'hc1be, 16'hc1bf 	:	val_out <= 16'h001d;
         16'hc1c0, 16'hc1c1, 16'hc1c2, 16'hc1c3, 16'hc1c4, 16'hc1c5, 16'hc1c6, 16'hc1c7 	:	val_out <= 16'h001e;
         16'hc1c8, 16'hc1c9, 16'hc1ca, 16'hc1cb, 16'hc1cc, 16'hc1cd, 16'hc1ce, 16'hc1cf 	:	val_out <= 16'h001f;
         16'hc1d0, 16'hc1d1, 16'hc1d2, 16'hc1d3, 16'hc1d4, 16'hc1d5, 16'hc1d6, 16'hc1d7 	:	val_out <= 16'h0020;
         16'hc1d8, 16'hc1d9, 16'hc1da, 16'hc1db, 16'hc1dc, 16'hc1dd, 16'hc1de, 16'hc1df 	:	val_out <= 16'h0021;
         16'hc1e0, 16'hc1e1, 16'hc1e2, 16'hc1e3, 16'hc1e4, 16'hc1e5, 16'hc1e6, 16'hc1e7 	:	val_out <= 16'h0022;
         16'hc1e8, 16'hc1e9, 16'hc1ea, 16'hc1eb, 16'hc1ec, 16'hc1ed, 16'hc1ee, 16'hc1ef 	:	val_out <= 16'h0023;
         16'hc1f0, 16'hc1f1, 16'hc1f2, 16'hc1f3, 16'hc1f4, 16'hc1f5, 16'hc1f6, 16'hc1f7 	:	val_out <= 16'h0025;
         16'hc1f8, 16'hc1f9, 16'hc1fa, 16'hc1fb, 16'hc1fc, 16'hc1fd, 16'hc1fe, 16'hc1ff 	:	val_out <= 16'h0026;
         16'hc200, 16'hc201, 16'hc202, 16'hc203, 16'hc204, 16'hc205, 16'hc206, 16'hc207 	:	val_out <= 16'h0027;
         16'hc208, 16'hc209, 16'hc20a, 16'hc20b, 16'hc20c, 16'hc20d, 16'hc20e, 16'hc20f 	:	val_out <= 16'h0028;
         16'hc210, 16'hc211, 16'hc212, 16'hc213, 16'hc214, 16'hc215, 16'hc216, 16'hc217 	:	val_out <= 16'h0029;
         16'hc218, 16'hc219, 16'hc21a, 16'hc21b, 16'hc21c, 16'hc21d, 16'hc21e, 16'hc21f 	:	val_out <= 16'h002b;
         16'hc220, 16'hc221, 16'hc222, 16'hc223, 16'hc224, 16'hc225, 16'hc226, 16'hc227 	:	val_out <= 16'h002c;
         16'hc228, 16'hc229, 16'hc22a, 16'hc22b, 16'hc22c, 16'hc22d, 16'hc22e, 16'hc22f 	:	val_out <= 16'h002d;
         16'hc230, 16'hc231, 16'hc232, 16'hc233, 16'hc234, 16'hc235, 16'hc236, 16'hc237 	:	val_out <= 16'h002f;
         16'hc238, 16'hc239, 16'hc23a, 16'hc23b, 16'hc23c, 16'hc23d, 16'hc23e, 16'hc23f 	:	val_out <= 16'h0030;
         16'hc240, 16'hc241, 16'hc242, 16'hc243, 16'hc244, 16'hc245, 16'hc246, 16'hc247 	:	val_out <= 16'h0031;
         16'hc248, 16'hc249, 16'hc24a, 16'hc24b, 16'hc24c, 16'hc24d, 16'hc24e, 16'hc24f 	:	val_out <= 16'h0033;
         16'hc250, 16'hc251, 16'hc252, 16'hc253, 16'hc254, 16'hc255, 16'hc256, 16'hc257 	:	val_out <= 16'h0034;
         16'hc258, 16'hc259, 16'hc25a, 16'hc25b, 16'hc25c, 16'hc25d, 16'hc25e, 16'hc25f 	:	val_out <= 16'h0036;
         16'hc260, 16'hc261, 16'hc262, 16'hc263, 16'hc264, 16'hc265, 16'hc266, 16'hc267 	:	val_out <= 16'h0037;
         16'hc268, 16'hc269, 16'hc26a, 16'hc26b, 16'hc26c, 16'hc26d, 16'hc26e, 16'hc26f 	:	val_out <= 16'h0039;
         16'hc270, 16'hc271, 16'hc272, 16'hc273, 16'hc274, 16'hc275, 16'hc276, 16'hc277 	:	val_out <= 16'h003a;
         16'hc278, 16'hc279, 16'hc27a, 16'hc27b, 16'hc27c, 16'hc27d, 16'hc27e, 16'hc27f 	:	val_out <= 16'h003c;
         16'hc280, 16'hc281, 16'hc282, 16'hc283, 16'hc284, 16'hc285, 16'hc286, 16'hc287 	:	val_out <= 16'h003d;
         16'hc288, 16'hc289, 16'hc28a, 16'hc28b, 16'hc28c, 16'hc28d, 16'hc28e, 16'hc28f 	:	val_out <= 16'h003f;
         16'hc290, 16'hc291, 16'hc292, 16'hc293, 16'hc294, 16'hc295, 16'hc296, 16'hc297 	:	val_out <= 16'h0040;
         16'hc298, 16'hc299, 16'hc29a, 16'hc29b, 16'hc29c, 16'hc29d, 16'hc29e, 16'hc29f 	:	val_out <= 16'h0042;
         16'hc2a0, 16'hc2a1, 16'hc2a2, 16'hc2a3, 16'hc2a4, 16'hc2a5, 16'hc2a6, 16'hc2a7 	:	val_out <= 16'h0043;
         16'hc2a8, 16'hc2a9, 16'hc2aa, 16'hc2ab, 16'hc2ac, 16'hc2ad, 16'hc2ae, 16'hc2af 	:	val_out <= 16'h0045;
         16'hc2b0, 16'hc2b1, 16'hc2b2, 16'hc2b3, 16'hc2b4, 16'hc2b5, 16'hc2b6, 16'hc2b7 	:	val_out <= 16'h0047;
         16'hc2b8, 16'hc2b9, 16'hc2ba, 16'hc2bb, 16'hc2bc, 16'hc2bd, 16'hc2be, 16'hc2bf 	:	val_out <= 16'h0048;
         16'hc2c0, 16'hc2c1, 16'hc2c2, 16'hc2c3, 16'hc2c4, 16'hc2c5, 16'hc2c6, 16'hc2c7 	:	val_out <= 16'h004a;
         16'hc2c8, 16'hc2c9, 16'hc2ca, 16'hc2cb, 16'hc2cc, 16'hc2cd, 16'hc2ce, 16'hc2cf 	:	val_out <= 16'h004c;
         16'hc2d0, 16'hc2d1, 16'hc2d2, 16'hc2d3, 16'hc2d4, 16'hc2d5, 16'hc2d6, 16'hc2d7 	:	val_out <= 16'h004e;
         16'hc2d8, 16'hc2d9, 16'hc2da, 16'hc2db, 16'hc2dc, 16'hc2dd, 16'hc2de, 16'hc2df 	:	val_out <= 16'h004f;
         16'hc2e0, 16'hc2e1, 16'hc2e2, 16'hc2e3, 16'hc2e4, 16'hc2e5, 16'hc2e6, 16'hc2e7 	:	val_out <= 16'h0051;
         16'hc2e8, 16'hc2e9, 16'hc2ea, 16'hc2eb, 16'hc2ec, 16'hc2ed, 16'hc2ee, 16'hc2ef 	:	val_out <= 16'h0053;
         16'hc2f0, 16'hc2f1, 16'hc2f2, 16'hc2f3, 16'hc2f4, 16'hc2f5, 16'hc2f6, 16'hc2f7 	:	val_out <= 16'h0055;
         16'hc2f8, 16'hc2f9, 16'hc2fa, 16'hc2fb, 16'hc2fc, 16'hc2fd, 16'hc2fe, 16'hc2ff 	:	val_out <= 16'h0056;
         16'hc300, 16'hc301, 16'hc302, 16'hc303, 16'hc304, 16'hc305, 16'hc306, 16'hc307 	:	val_out <= 16'h0058;
         16'hc308, 16'hc309, 16'hc30a, 16'hc30b, 16'hc30c, 16'hc30d, 16'hc30e, 16'hc30f 	:	val_out <= 16'h005a;
         16'hc310, 16'hc311, 16'hc312, 16'hc313, 16'hc314, 16'hc315, 16'hc316, 16'hc317 	:	val_out <= 16'h005c;
         16'hc318, 16'hc319, 16'hc31a, 16'hc31b, 16'hc31c, 16'hc31d, 16'hc31e, 16'hc31f 	:	val_out <= 16'h005e;
         16'hc320, 16'hc321, 16'hc322, 16'hc323, 16'hc324, 16'hc325, 16'hc326, 16'hc327 	:	val_out <= 16'h0060;
         16'hc328, 16'hc329, 16'hc32a, 16'hc32b, 16'hc32c, 16'hc32d, 16'hc32e, 16'hc32f 	:	val_out <= 16'h0062;
         16'hc330, 16'hc331, 16'hc332, 16'hc333, 16'hc334, 16'hc335, 16'hc336, 16'hc337 	:	val_out <= 16'h0064;
         16'hc338, 16'hc339, 16'hc33a, 16'hc33b, 16'hc33c, 16'hc33d, 16'hc33e, 16'hc33f 	:	val_out <= 16'h0066;
         16'hc340, 16'hc341, 16'hc342, 16'hc343, 16'hc344, 16'hc345, 16'hc346, 16'hc347 	:	val_out <= 16'h0068;
         16'hc348, 16'hc349, 16'hc34a, 16'hc34b, 16'hc34c, 16'hc34d, 16'hc34e, 16'hc34f 	:	val_out <= 16'h006a;
         16'hc350, 16'hc351, 16'hc352, 16'hc353, 16'hc354, 16'hc355, 16'hc356, 16'hc357 	:	val_out <= 16'h006c;
         16'hc358, 16'hc359, 16'hc35a, 16'hc35b, 16'hc35c, 16'hc35d, 16'hc35e, 16'hc35f 	:	val_out <= 16'h006e;
         16'hc360, 16'hc361, 16'hc362, 16'hc363, 16'hc364, 16'hc365, 16'hc366, 16'hc367 	:	val_out <= 16'h0070;
         16'hc368, 16'hc369, 16'hc36a, 16'hc36b, 16'hc36c, 16'hc36d, 16'hc36e, 16'hc36f 	:	val_out <= 16'h0072;
         16'hc370, 16'hc371, 16'hc372, 16'hc373, 16'hc374, 16'hc375, 16'hc376, 16'hc377 	:	val_out <= 16'h0074;
         16'hc378, 16'hc379, 16'hc37a, 16'hc37b, 16'hc37c, 16'hc37d, 16'hc37e, 16'hc37f 	:	val_out <= 16'h0076;
         16'hc380, 16'hc381, 16'hc382, 16'hc383, 16'hc384, 16'hc385, 16'hc386, 16'hc387 	:	val_out <= 16'h0078;
         16'hc388, 16'hc389, 16'hc38a, 16'hc38b, 16'hc38c, 16'hc38d, 16'hc38e, 16'hc38f 	:	val_out <= 16'h007a;
         16'hc390, 16'hc391, 16'hc392, 16'hc393, 16'hc394, 16'hc395, 16'hc396, 16'hc397 	:	val_out <= 16'h007d;
         16'hc398, 16'hc399, 16'hc39a, 16'hc39b, 16'hc39c, 16'hc39d, 16'hc39e, 16'hc39f 	:	val_out <= 16'h007f;
         16'hc3a0, 16'hc3a1, 16'hc3a2, 16'hc3a3, 16'hc3a4, 16'hc3a5, 16'hc3a6, 16'hc3a7 	:	val_out <= 16'h0081;
         16'hc3a8, 16'hc3a9, 16'hc3aa, 16'hc3ab, 16'hc3ac, 16'hc3ad, 16'hc3ae, 16'hc3af 	:	val_out <= 16'h0083;
         16'hc3b0, 16'hc3b1, 16'hc3b2, 16'hc3b3, 16'hc3b4, 16'hc3b5, 16'hc3b6, 16'hc3b7 	:	val_out <= 16'h0086;
         16'hc3b8, 16'hc3b9, 16'hc3ba, 16'hc3bb, 16'hc3bc, 16'hc3bd, 16'hc3be, 16'hc3bf 	:	val_out <= 16'h0088;
         16'hc3c0, 16'hc3c1, 16'hc3c2, 16'hc3c3, 16'hc3c4, 16'hc3c5, 16'hc3c6, 16'hc3c7 	:	val_out <= 16'h008a;
         16'hc3c8, 16'hc3c9, 16'hc3ca, 16'hc3cb, 16'hc3cc, 16'hc3cd, 16'hc3ce, 16'hc3cf 	:	val_out <= 16'h008d;
         16'hc3d0, 16'hc3d1, 16'hc3d2, 16'hc3d3, 16'hc3d4, 16'hc3d5, 16'hc3d6, 16'hc3d7 	:	val_out <= 16'h008f;
         16'hc3d8, 16'hc3d9, 16'hc3da, 16'hc3db, 16'hc3dc, 16'hc3dd, 16'hc3de, 16'hc3df 	:	val_out <= 16'h0091;
         16'hc3e0, 16'hc3e1, 16'hc3e2, 16'hc3e3, 16'hc3e4, 16'hc3e5, 16'hc3e6, 16'hc3e7 	:	val_out <= 16'h0094;
         16'hc3e8, 16'hc3e9, 16'hc3ea, 16'hc3eb, 16'hc3ec, 16'hc3ed, 16'hc3ee, 16'hc3ef 	:	val_out <= 16'h0096;
         16'hc3f0, 16'hc3f1, 16'hc3f2, 16'hc3f3, 16'hc3f4, 16'hc3f5, 16'hc3f6, 16'hc3f7 	:	val_out <= 16'h0098;
         16'hc3f8, 16'hc3f9, 16'hc3fa, 16'hc3fb, 16'hc3fc, 16'hc3fd, 16'hc3fe, 16'hc3ff 	:	val_out <= 16'h009b;
         16'hc400, 16'hc401, 16'hc402, 16'hc403, 16'hc404, 16'hc405, 16'hc406, 16'hc407 	:	val_out <= 16'h009d;
         16'hc408, 16'hc409, 16'hc40a, 16'hc40b, 16'hc40c, 16'hc40d, 16'hc40e, 16'hc40f 	:	val_out <= 16'h00a0;
         16'hc410, 16'hc411, 16'hc412, 16'hc413, 16'hc414, 16'hc415, 16'hc416, 16'hc417 	:	val_out <= 16'h00a2;
         16'hc418, 16'hc419, 16'hc41a, 16'hc41b, 16'hc41c, 16'hc41d, 16'hc41e, 16'hc41f 	:	val_out <= 16'h00a5;
         16'hc420, 16'hc421, 16'hc422, 16'hc423, 16'hc424, 16'hc425, 16'hc426, 16'hc427 	:	val_out <= 16'h00a7;
         16'hc428, 16'hc429, 16'hc42a, 16'hc42b, 16'hc42c, 16'hc42d, 16'hc42e, 16'hc42f 	:	val_out <= 16'h00aa;
         16'hc430, 16'hc431, 16'hc432, 16'hc433, 16'hc434, 16'hc435, 16'hc436, 16'hc437 	:	val_out <= 16'h00ac;
         16'hc438, 16'hc439, 16'hc43a, 16'hc43b, 16'hc43c, 16'hc43d, 16'hc43e, 16'hc43f 	:	val_out <= 16'h00af;
         16'hc440, 16'hc441, 16'hc442, 16'hc443, 16'hc444, 16'hc445, 16'hc446, 16'hc447 	:	val_out <= 16'h00b2;
         16'hc448, 16'hc449, 16'hc44a, 16'hc44b, 16'hc44c, 16'hc44d, 16'hc44e, 16'hc44f 	:	val_out <= 16'h00b4;
         16'hc450, 16'hc451, 16'hc452, 16'hc453, 16'hc454, 16'hc455, 16'hc456, 16'hc457 	:	val_out <= 16'h00b7;
         16'hc458, 16'hc459, 16'hc45a, 16'hc45b, 16'hc45c, 16'hc45d, 16'hc45e, 16'hc45f 	:	val_out <= 16'h00ba;
         16'hc460, 16'hc461, 16'hc462, 16'hc463, 16'hc464, 16'hc465, 16'hc466, 16'hc467 	:	val_out <= 16'h00bc;
         16'hc468, 16'hc469, 16'hc46a, 16'hc46b, 16'hc46c, 16'hc46d, 16'hc46e, 16'hc46f 	:	val_out <= 16'h00bf;
         16'hc470, 16'hc471, 16'hc472, 16'hc473, 16'hc474, 16'hc475, 16'hc476, 16'hc477 	:	val_out <= 16'h00c2;
         16'hc478, 16'hc479, 16'hc47a, 16'hc47b, 16'hc47c, 16'hc47d, 16'hc47e, 16'hc47f 	:	val_out <= 16'h00c4;
         16'hc480, 16'hc481, 16'hc482, 16'hc483, 16'hc484, 16'hc485, 16'hc486, 16'hc487 	:	val_out <= 16'h00c7;
         16'hc488, 16'hc489, 16'hc48a, 16'hc48b, 16'hc48c, 16'hc48d, 16'hc48e, 16'hc48f 	:	val_out <= 16'h00ca;
         16'hc490, 16'hc491, 16'hc492, 16'hc493, 16'hc494, 16'hc495, 16'hc496, 16'hc497 	:	val_out <= 16'h00cd;
         16'hc498, 16'hc499, 16'hc49a, 16'hc49b, 16'hc49c, 16'hc49d, 16'hc49e, 16'hc49f 	:	val_out <= 16'h00d0;
         16'hc4a0, 16'hc4a1, 16'hc4a2, 16'hc4a3, 16'hc4a4, 16'hc4a5, 16'hc4a6, 16'hc4a7 	:	val_out <= 16'h00d2;
         16'hc4a8, 16'hc4a9, 16'hc4aa, 16'hc4ab, 16'hc4ac, 16'hc4ad, 16'hc4ae, 16'hc4af 	:	val_out <= 16'h00d5;
         16'hc4b0, 16'hc4b1, 16'hc4b2, 16'hc4b3, 16'hc4b4, 16'hc4b5, 16'hc4b6, 16'hc4b7 	:	val_out <= 16'h00d8;
         16'hc4b8, 16'hc4b9, 16'hc4ba, 16'hc4bb, 16'hc4bc, 16'hc4bd, 16'hc4be, 16'hc4bf 	:	val_out <= 16'h00db;
         16'hc4c0, 16'hc4c1, 16'hc4c2, 16'hc4c3, 16'hc4c4, 16'hc4c5, 16'hc4c6, 16'hc4c7 	:	val_out <= 16'h00de;
         16'hc4c8, 16'hc4c9, 16'hc4ca, 16'hc4cb, 16'hc4cc, 16'hc4cd, 16'hc4ce, 16'hc4cf 	:	val_out <= 16'h00e1;
         16'hc4d0, 16'hc4d1, 16'hc4d2, 16'hc4d3, 16'hc4d4, 16'hc4d5, 16'hc4d6, 16'hc4d7 	:	val_out <= 16'h00e4;
         16'hc4d8, 16'hc4d9, 16'hc4da, 16'hc4db, 16'hc4dc, 16'hc4dd, 16'hc4de, 16'hc4df 	:	val_out <= 16'h00e7;
         16'hc4e0, 16'hc4e1, 16'hc4e2, 16'hc4e3, 16'hc4e4, 16'hc4e5, 16'hc4e6, 16'hc4e7 	:	val_out <= 16'h00ea;
         16'hc4e8, 16'hc4e9, 16'hc4ea, 16'hc4eb, 16'hc4ec, 16'hc4ed, 16'hc4ee, 16'hc4ef 	:	val_out <= 16'h00ed;
         16'hc4f0, 16'hc4f1, 16'hc4f2, 16'hc4f3, 16'hc4f4, 16'hc4f5, 16'hc4f6, 16'hc4f7 	:	val_out <= 16'h00f0;
         16'hc4f8, 16'hc4f9, 16'hc4fa, 16'hc4fb, 16'hc4fc, 16'hc4fd, 16'hc4fe, 16'hc4ff 	:	val_out <= 16'h00f3;
         16'hc500, 16'hc501, 16'hc502, 16'hc503, 16'hc504, 16'hc505, 16'hc506, 16'hc507 	:	val_out <= 16'h00f6;
         16'hc508, 16'hc509, 16'hc50a, 16'hc50b, 16'hc50c, 16'hc50d, 16'hc50e, 16'hc50f 	:	val_out <= 16'h00f9;
         16'hc510, 16'hc511, 16'hc512, 16'hc513, 16'hc514, 16'hc515, 16'hc516, 16'hc517 	:	val_out <= 16'h00fc;
         16'hc518, 16'hc519, 16'hc51a, 16'hc51b, 16'hc51c, 16'hc51d, 16'hc51e, 16'hc51f 	:	val_out <= 16'h00ff;
         16'hc520, 16'hc521, 16'hc522, 16'hc523, 16'hc524, 16'hc525, 16'hc526, 16'hc527 	:	val_out <= 16'h0102;
         16'hc528, 16'hc529, 16'hc52a, 16'hc52b, 16'hc52c, 16'hc52d, 16'hc52e, 16'hc52f 	:	val_out <= 16'h0106;
         16'hc530, 16'hc531, 16'hc532, 16'hc533, 16'hc534, 16'hc535, 16'hc536, 16'hc537 	:	val_out <= 16'h0109;
         16'hc538, 16'hc539, 16'hc53a, 16'hc53b, 16'hc53c, 16'hc53d, 16'hc53e, 16'hc53f 	:	val_out <= 16'h010c;
         16'hc540, 16'hc541, 16'hc542, 16'hc543, 16'hc544, 16'hc545, 16'hc546, 16'hc547 	:	val_out <= 16'h010f;
         16'hc548, 16'hc549, 16'hc54a, 16'hc54b, 16'hc54c, 16'hc54d, 16'hc54e, 16'hc54f 	:	val_out <= 16'h0112;
         16'hc550, 16'hc551, 16'hc552, 16'hc553, 16'hc554, 16'hc555, 16'hc556, 16'hc557 	:	val_out <= 16'h0116;
         16'hc558, 16'hc559, 16'hc55a, 16'hc55b, 16'hc55c, 16'hc55d, 16'hc55e, 16'hc55f 	:	val_out <= 16'h0119;
         16'hc560, 16'hc561, 16'hc562, 16'hc563, 16'hc564, 16'hc565, 16'hc566, 16'hc567 	:	val_out <= 16'h011c;
         16'hc568, 16'hc569, 16'hc56a, 16'hc56b, 16'hc56c, 16'hc56d, 16'hc56e, 16'hc56f 	:	val_out <= 16'h0120;
         16'hc570, 16'hc571, 16'hc572, 16'hc573, 16'hc574, 16'hc575, 16'hc576, 16'hc577 	:	val_out <= 16'h0123;
         16'hc578, 16'hc579, 16'hc57a, 16'hc57b, 16'hc57c, 16'hc57d, 16'hc57e, 16'hc57f 	:	val_out <= 16'h0126;
         16'hc580, 16'hc581, 16'hc582, 16'hc583, 16'hc584, 16'hc585, 16'hc586, 16'hc587 	:	val_out <= 16'h012a;
         16'hc588, 16'hc589, 16'hc58a, 16'hc58b, 16'hc58c, 16'hc58d, 16'hc58e, 16'hc58f 	:	val_out <= 16'h012d;
         16'hc590, 16'hc591, 16'hc592, 16'hc593, 16'hc594, 16'hc595, 16'hc596, 16'hc597 	:	val_out <= 16'h0130;
         16'hc598, 16'hc599, 16'hc59a, 16'hc59b, 16'hc59c, 16'hc59d, 16'hc59e, 16'hc59f 	:	val_out <= 16'h0134;
         16'hc5a0, 16'hc5a1, 16'hc5a2, 16'hc5a3, 16'hc5a4, 16'hc5a5, 16'hc5a6, 16'hc5a7 	:	val_out <= 16'h0137;
         16'hc5a8, 16'hc5a9, 16'hc5aa, 16'hc5ab, 16'hc5ac, 16'hc5ad, 16'hc5ae, 16'hc5af 	:	val_out <= 16'h013b;
         16'hc5b0, 16'hc5b1, 16'hc5b2, 16'hc5b3, 16'hc5b4, 16'hc5b5, 16'hc5b6, 16'hc5b7 	:	val_out <= 16'h013e;
         16'hc5b8, 16'hc5b9, 16'hc5ba, 16'hc5bb, 16'hc5bc, 16'hc5bd, 16'hc5be, 16'hc5bf 	:	val_out <= 16'h0142;
         16'hc5c0, 16'hc5c1, 16'hc5c2, 16'hc5c3, 16'hc5c4, 16'hc5c5, 16'hc5c6, 16'hc5c7 	:	val_out <= 16'h0145;
         16'hc5c8, 16'hc5c9, 16'hc5ca, 16'hc5cb, 16'hc5cc, 16'hc5cd, 16'hc5ce, 16'hc5cf 	:	val_out <= 16'h0149;
         16'hc5d0, 16'hc5d1, 16'hc5d2, 16'hc5d3, 16'hc5d4, 16'hc5d5, 16'hc5d6, 16'hc5d7 	:	val_out <= 16'h014c;
         16'hc5d8, 16'hc5d9, 16'hc5da, 16'hc5db, 16'hc5dc, 16'hc5dd, 16'hc5de, 16'hc5df 	:	val_out <= 16'h0150;
         16'hc5e0, 16'hc5e1, 16'hc5e2, 16'hc5e3, 16'hc5e4, 16'hc5e5, 16'hc5e6, 16'hc5e7 	:	val_out <= 16'h0154;
         16'hc5e8, 16'hc5e9, 16'hc5ea, 16'hc5eb, 16'hc5ec, 16'hc5ed, 16'hc5ee, 16'hc5ef 	:	val_out <= 16'h0157;
         16'hc5f0, 16'hc5f1, 16'hc5f2, 16'hc5f3, 16'hc5f4, 16'hc5f5, 16'hc5f6, 16'hc5f7 	:	val_out <= 16'h015b;
         16'hc5f8, 16'hc5f9, 16'hc5fa, 16'hc5fb, 16'hc5fc, 16'hc5fd, 16'hc5fe, 16'hc5ff 	:	val_out <= 16'h015e;
         16'hc600, 16'hc601, 16'hc602, 16'hc603, 16'hc604, 16'hc605, 16'hc606, 16'hc607 	:	val_out <= 16'h0162;
         16'hc608, 16'hc609, 16'hc60a, 16'hc60b, 16'hc60c, 16'hc60d, 16'hc60e, 16'hc60f 	:	val_out <= 16'h0166;
         16'hc610, 16'hc611, 16'hc612, 16'hc613, 16'hc614, 16'hc615, 16'hc616, 16'hc617 	:	val_out <= 16'h016a;
         16'hc618, 16'hc619, 16'hc61a, 16'hc61b, 16'hc61c, 16'hc61d, 16'hc61e, 16'hc61f 	:	val_out <= 16'h016d;
         16'hc620, 16'hc621, 16'hc622, 16'hc623, 16'hc624, 16'hc625, 16'hc626, 16'hc627 	:	val_out <= 16'h0171;
         16'hc628, 16'hc629, 16'hc62a, 16'hc62b, 16'hc62c, 16'hc62d, 16'hc62e, 16'hc62f 	:	val_out <= 16'h0175;
         16'hc630, 16'hc631, 16'hc632, 16'hc633, 16'hc634, 16'hc635, 16'hc636, 16'hc637 	:	val_out <= 16'h0179;
         16'hc638, 16'hc639, 16'hc63a, 16'hc63b, 16'hc63c, 16'hc63d, 16'hc63e, 16'hc63f 	:	val_out <= 16'h017c;
         16'hc640, 16'hc641, 16'hc642, 16'hc643, 16'hc644, 16'hc645, 16'hc646, 16'hc647 	:	val_out <= 16'h0180;
         16'hc648, 16'hc649, 16'hc64a, 16'hc64b, 16'hc64c, 16'hc64d, 16'hc64e, 16'hc64f 	:	val_out <= 16'h0184;
         16'hc650, 16'hc651, 16'hc652, 16'hc653, 16'hc654, 16'hc655, 16'hc656, 16'hc657 	:	val_out <= 16'h0188;
         16'hc658, 16'hc659, 16'hc65a, 16'hc65b, 16'hc65c, 16'hc65d, 16'hc65e, 16'hc65f 	:	val_out <= 16'h018c;
         16'hc660, 16'hc661, 16'hc662, 16'hc663, 16'hc664, 16'hc665, 16'hc666, 16'hc667 	:	val_out <= 16'h0190;
         16'hc668, 16'hc669, 16'hc66a, 16'hc66b, 16'hc66c, 16'hc66d, 16'hc66e, 16'hc66f 	:	val_out <= 16'h0194;
         16'hc670, 16'hc671, 16'hc672, 16'hc673, 16'hc674, 16'hc675, 16'hc676, 16'hc677 	:	val_out <= 16'h0198;
         16'hc678, 16'hc679, 16'hc67a, 16'hc67b, 16'hc67c, 16'hc67d, 16'hc67e, 16'hc67f 	:	val_out <= 16'h019c;
         16'hc680, 16'hc681, 16'hc682, 16'hc683, 16'hc684, 16'hc685, 16'hc686, 16'hc687 	:	val_out <= 16'h01a0;
         16'hc688, 16'hc689, 16'hc68a, 16'hc68b, 16'hc68c, 16'hc68d, 16'hc68e, 16'hc68f 	:	val_out <= 16'h01a4;
         16'hc690, 16'hc691, 16'hc692, 16'hc693, 16'hc694, 16'hc695, 16'hc696, 16'hc697 	:	val_out <= 16'h01a8;
         16'hc698, 16'hc699, 16'hc69a, 16'hc69b, 16'hc69c, 16'hc69d, 16'hc69e, 16'hc69f 	:	val_out <= 16'h01ac;
         16'hc6a0, 16'hc6a1, 16'hc6a2, 16'hc6a3, 16'hc6a4, 16'hc6a5, 16'hc6a6, 16'hc6a7 	:	val_out <= 16'h01b0;
         16'hc6a8, 16'hc6a9, 16'hc6aa, 16'hc6ab, 16'hc6ac, 16'hc6ad, 16'hc6ae, 16'hc6af 	:	val_out <= 16'h01b4;
         16'hc6b0, 16'hc6b1, 16'hc6b2, 16'hc6b3, 16'hc6b4, 16'hc6b5, 16'hc6b6, 16'hc6b7 	:	val_out <= 16'h01b8;
         16'hc6b8, 16'hc6b9, 16'hc6ba, 16'hc6bb, 16'hc6bc, 16'hc6bd, 16'hc6be, 16'hc6bf 	:	val_out <= 16'h01bc;
         16'hc6c0, 16'hc6c1, 16'hc6c2, 16'hc6c3, 16'hc6c4, 16'hc6c5, 16'hc6c6, 16'hc6c7 	:	val_out <= 16'h01c0;
         16'hc6c8, 16'hc6c9, 16'hc6ca, 16'hc6cb, 16'hc6cc, 16'hc6cd, 16'hc6ce, 16'hc6cf 	:	val_out <= 16'h01c4;
         16'hc6d0, 16'hc6d1, 16'hc6d2, 16'hc6d3, 16'hc6d4, 16'hc6d5, 16'hc6d6, 16'hc6d7 	:	val_out <= 16'h01c8;
         16'hc6d8, 16'hc6d9, 16'hc6da, 16'hc6db, 16'hc6dc, 16'hc6dd, 16'hc6de, 16'hc6df 	:	val_out <= 16'h01cd;
         16'hc6e0, 16'hc6e1, 16'hc6e2, 16'hc6e3, 16'hc6e4, 16'hc6e5, 16'hc6e6, 16'hc6e7 	:	val_out <= 16'h01d1;
         16'hc6e8, 16'hc6e9, 16'hc6ea, 16'hc6eb, 16'hc6ec, 16'hc6ed, 16'hc6ee, 16'hc6ef 	:	val_out <= 16'h01d5;
         16'hc6f0, 16'hc6f1, 16'hc6f2, 16'hc6f3, 16'hc6f4, 16'hc6f5, 16'hc6f6, 16'hc6f7 	:	val_out <= 16'h01d9;
         16'hc6f8, 16'hc6f9, 16'hc6fa, 16'hc6fb, 16'hc6fc, 16'hc6fd, 16'hc6fe, 16'hc6ff 	:	val_out <= 16'h01de;
         16'hc700, 16'hc701, 16'hc702, 16'hc703, 16'hc704, 16'hc705, 16'hc706, 16'hc707 	:	val_out <= 16'h01e2;
         16'hc708, 16'hc709, 16'hc70a, 16'hc70b, 16'hc70c, 16'hc70d, 16'hc70e, 16'hc70f 	:	val_out <= 16'h01e6;
         16'hc710, 16'hc711, 16'hc712, 16'hc713, 16'hc714, 16'hc715, 16'hc716, 16'hc717 	:	val_out <= 16'h01eb;
         16'hc718, 16'hc719, 16'hc71a, 16'hc71b, 16'hc71c, 16'hc71d, 16'hc71e, 16'hc71f 	:	val_out <= 16'h01ef;
         16'hc720, 16'hc721, 16'hc722, 16'hc723, 16'hc724, 16'hc725, 16'hc726, 16'hc727 	:	val_out <= 16'h01f3;
         16'hc728, 16'hc729, 16'hc72a, 16'hc72b, 16'hc72c, 16'hc72d, 16'hc72e, 16'hc72f 	:	val_out <= 16'h01f8;
         16'hc730, 16'hc731, 16'hc732, 16'hc733, 16'hc734, 16'hc735, 16'hc736, 16'hc737 	:	val_out <= 16'h01fc;
         16'hc738, 16'hc739, 16'hc73a, 16'hc73b, 16'hc73c, 16'hc73d, 16'hc73e, 16'hc73f 	:	val_out <= 16'h0200;
         16'hc740, 16'hc741, 16'hc742, 16'hc743, 16'hc744, 16'hc745, 16'hc746, 16'hc747 	:	val_out <= 16'h0205;
         16'hc748, 16'hc749, 16'hc74a, 16'hc74b, 16'hc74c, 16'hc74d, 16'hc74e, 16'hc74f 	:	val_out <= 16'h0209;
         16'hc750, 16'hc751, 16'hc752, 16'hc753, 16'hc754, 16'hc755, 16'hc756, 16'hc757 	:	val_out <= 16'h020e;
         16'hc758, 16'hc759, 16'hc75a, 16'hc75b, 16'hc75c, 16'hc75d, 16'hc75e, 16'hc75f 	:	val_out <= 16'h0212;
         16'hc760, 16'hc761, 16'hc762, 16'hc763, 16'hc764, 16'hc765, 16'hc766, 16'hc767 	:	val_out <= 16'h0217;
         16'hc768, 16'hc769, 16'hc76a, 16'hc76b, 16'hc76c, 16'hc76d, 16'hc76e, 16'hc76f 	:	val_out <= 16'h021b;
         16'hc770, 16'hc771, 16'hc772, 16'hc773, 16'hc774, 16'hc775, 16'hc776, 16'hc777 	:	val_out <= 16'h0220;
         16'hc778, 16'hc779, 16'hc77a, 16'hc77b, 16'hc77c, 16'hc77d, 16'hc77e, 16'hc77f 	:	val_out <= 16'h0225;
         16'hc780, 16'hc781, 16'hc782, 16'hc783, 16'hc784, 16'hc785, 16'hc786, 16'hc787 	:	val_out <= 16'h0229;
         16'hc788, 16'hc789, 16'hc78a, 16'hc78b, 16'hc78c, 16'hc78d, 16'hc78e, 16'hc78f 	:	val_out <= 16'h022e;
         16'hc790, 16'hc791, 16'hc792, 16'hc793, 16'hc794, 16'hc795, 16'hc796, 16'hc797 	:	val_out <= 16'h0232;
         16'hc798, 16'hc799, 16'hc79a, 16'hc79b, 16'hc79c, 16'hc79d, 16'hc79e, 16'hc79f 	:	val_out <= 16'h0237;
         16'hc7a0, 16'hc7a1, 16'hc7a2, 16'hc7a3, 16'hc7a4, 16'hc7a5, 16'hc7a6, 16'hc7a7 	:	val_out <= 16'h023c;
         16'hc7a8, 16'hc7a9, 16'hc7aa, 16'hc7ab, 16'hc7ac, 16'hc7ad, 16'hc7ae, 16'hc7af 	:	val_out <= 16'h0240;
         16'hc7b0, 16'hc7b1, 16'hc7b2, 16'hc7b3, 16'hc7b4, 16'hc7b5, 16'hc7b6, 16'hc7b7 	:	val_out <= 16'h0245;
         16'hc7b8, 16'hc7b9, 16'hc7ba, 16'hc7bb, 16'hc7bc, 16'hc7bd, 16'hc7be, 16'hc7bf 	:	val_out <= 16'h024a;
         16'hc7c0, 16'hc7c1, 16'hc7c2, 16'hc7c3, 16'hc7c4, 16'hc7c5, 16'hc7c6, 16'hc7c7 	:	val_out <= 16'h024f;
         16'hc7c8, 16'hc7c9, 16'hc7ca, 16'hc7cb, 16'hc7cc, 16'hc7cd, 16'hc7ce, 16'hc7cf 	:	val_out <= 16'h0253;
         16'hc7d0, 16'hc7d1, 16'hc7d2, 16'hc7d3, 16'hc7d4, 16'hc7d5, 16'hc7d6, 16'hc7d7 	:	val_out <= 16'h0258;
         16'hc7d8, 16'hc7d9, 16'hc7da, 16'hc7db, 16'hc7dc, 16'hc7dd, 16'hc7de, 16'hc7df 	:	val_out <= 16'h025d;
         16'hc7e0, 16'hc7e1, 16'hc7e2, 16'hc7e3, 16'hc7e4, 16'hc7e5, 16'hc7e6, 16'hc7e7 	:	val_out <= 16'h0262;
         16'hc7e8, 16'hc7e9, 16'hc7ea, 16'hc7eb, 16'hc7ec, 16'hc7ed, 16'hc7ee, 16'hc7ef 	:	val_out <= 16'h0267;
         16'hc7f0, 16'hc7f1, 16'hc7f2, 16'hc7f3, 16'hc7f4, 16'hc7f5, 16'hc7f6, 16'hc7f7 	:	val_out <= 16'h026b;
         16'hc7f8, 16'hc7f9, 16'hc7fa, 16'hc7fb, 16'hc7fc, 16'hc7fd, 16'hc7fe, 16'hc7ff 	:	val_out <= 16'h0270;
         16'hc800, 16'hc801, 16'hc802, 16'hc803, 16'hc804, 16'hc805, 16'hc806, 16'hc807 	:	val_out <= 16'h0275;
         16'hc808, 16'hc809, 16'hc80a, 16'hc80b, 16'hc80c, 16'hc80d, 16'hc80e, 16'hc80f 	:	val_out <= 16'h027a;
         16'hc810, 16'hc811, 16'hc812, 16'hc813, 16'hc814, 16'hc815, 16'hc816, 16'hc817 	:	val_out <= 16'h027f;
         16'hc818, 16'hc819, 16'hc81a, 16'hc81b, 16'hc81c, 16'hc81d, 16'hc81e, 16'hc81f 	:	val_out <= 16'h0284;
         16'hc820, 16'hc821, 16'hc822, 16'hc823, 16'hc824, 16'hc825, 16'hc826, 16'hc827 	:	val_out <= 16'h0289;
         16'hc828, 16'hc829, 16'hc82a, 16'hc82b, 16'hc82c, 16'hc82d, 16'hc82e, 16'hc82f 	:	val_out <= 16'h028e;
         16'hc830, 16'hc831, 16'hc832, 16'hc833, 16'hc834, 16'hc835, 16'hc836, 16'hc837 	:	val_out <= 16'h0293;
         16'hc838, 16'hc839, 16'hc83a, 16'hc83b, 16'hc83c, 16'hc83d, 16'hc83e, 16'hc83f 	:	val_out <= 16'h0298;
         16'hc840, 16'hc841, 16'hc842, 16'hc843, 16'hc844, 16'hc845, 16'hc846, 16'hc847 	:	val_out <= 16'h029d;
         16'hc848, 16'hc849, 16'hc84a, 16'hc84b, 16'hc84c, 16'hc84d, 16'hc84e, 16'hc84f 	:	val_out <= 16'h02a2;
         16'hc850, 16'hc851, 16'hc852, 16'hc853, 16'hc854, 16'hc855, 16'hc856, 16'hc857 	:	val_out <= 16'h02a7;
         16'hc858, 16'hc859, 16'hc85a, 16'hc85b, 16'hc85c, 16'hc85d, 16'hc85e, 16'hc85f 	:	val_out <= 16'h02ac;
         16'hc860, 16'hc861, 16'hc862, 16'hc863, 16'hc864, 16'hc865, 16'hc866, 16'hc867 	:	val_out <= 16'h02b1;
         16'hc868, 16'hc869, 16'hc86a, 16'hc86b, 16'hc86c, 16'hc86d, 16'hc86e, 16'hc86f 	:	val_out <= 16'h02b6;
         16'hc870, 16'hc871, 16'hc872, 16'hc873, 16'hc874, 16'hc875, 16'hc876, 16'hc877 	:	val_out <= 16'h02bc;
         16'hc878, 16'hc879, 16'hc87a, 16'hc87b, 16'hc87c, 16'hc87d, 16'hc87e, 16'hc87f 	:	val_out <= 16'h02c1;
         16'hc880, 16'hc881, 16'hc882, 16'hc883, 16'hc884, 16'hc885, 16'hc886, 16'hc887 	:	val_out <= 16'h02c6;
         16'hc888, 16'hc889, 16'hc88a, 16'hc88b, 16'hc88c, 16'hc88d, 16'hc88e, 16'hc88f 	:	val_out <= 16'h02cb;
         16'hc890, 16'hc891, 16'hc892, 16'hc893, 16'hc894, 16'hc895, 16'hc896, 16'hc897 	:	val_out <= 16'h02d0;
         16'hc898, 16'hc899, 16'hc89a, 16'hc89b, 16'hc89c, 16'hc89d, 16'hc89e, 16'hc89f 	:	val_out <= 16'h02d6;
         16'hc8a0, 16'hc8a1, 16'hc8a2, 16'hc8a3, 16'hc8a4, 16'hc8a5, 16'hc8a6, 16'hc8a7 	:	val_out <= 16'h02db;
         16'hc8a8, 16'hc8a9, 16'hc8aa, 16'hc8ab, 16'hc8ac, 16'hc8ad, 16'hc8ae, 16'hc8af 	:	val_out <= 16'h02e0;
         16'hc8b0, 16'hc8b1, 16'hc8b2, 16'hc8b3, 16'hc8b4, 16'hc8b5, 16'hc8b6, 16'hc8b7 	:	val_out <= 16'h02e6;
         16'hc8b8, 16'hc8b9, 16'hc8ba, 16'hc8bb, 16'hc8bc, 16'hc8bd, 16'hc8be, 16'hc8bf 	:	val_out <= 16'h02eb;
         16'hc8c0, 16'hc8c1, 16'hc8c2, 16'hc8c3, 16'hc8c4, 16'hc8c5, 16'hc8c6, 16'hc8c7 	:	val_out <= 16'h02f0;
         16'hc8c8, 16'hc8c9, 16'hc8ca, 16'hc8cb, 16'hc8cc, 16'hc8cd, 16'hc8ce, 16'hc8cf 	:	val_out <= 16'h02f6;
         16'hc8d0, 16'hc8d1, 16'hc8d2, 16'hc8d3, 16'hc8d4, 16'hc8d5, 16'hc8d6, 16'hc8d7 	:	val_out <= 16'h02fb;
         16'hc8d8, 16'hc8d9, 16'hc8da, 16'hc8db, 16'hc8dc, 16'hc8dd, 16'hc8de, 16'hc8df 	:	val_out <= 16'h0300;
         16'hc8e0, 16'hc8e1, 16'hc8e2, 16'hc8e3, 16'hc8e4, 16'hc8e5, 16'hc8e6, 16'hc8e7 	:	val_out <= 16'h0306;
         16'hc8e8, 16'hc8e9, 16'hc8ea, 16'hc8eb, 16'hc8ec, 16'hc8ed, 16'hc8ee, 16'hc8ef 	:	val_out <= 16'h030b;
         16'hc8f0, 16'hc8f1, 16'hc8f2, 16'hc8f3, 16'hc8f4, 16'hc8f5, 16'hc8f6, 16'hc8f7 	:	val_out <= 16'h0311;
         16'hc8f8, 16'hc8f9, 16'hc8fa, 16'hc8fb, 16'hc8fc, 16'hc8fd, 16'hc8fe, 16'hc8ff 	:	val_out <= 16'h0316;
         16'hc900, 16'hc901, 16'hc902, 16'hc903, 16'hc904, 16'hc905, 16'hc906, 16'hc907 	:	val_out <= 16'h031c;
         16'hc908, 16'hc909, 16'hc90a, 16'hc90b, 16'hc90c, 16'hc90d, 16'hc90e, 16'hc90f 	:	val_out <= 16'h0321;
         16'hc910, 16'hc911, 16'hc912, 16'hc913, 16'hc914, 16'hc915, 16'hc916, 16'hc917 	:	val_out <= 16'h0327;
         16'hc918, 16'hc919, 16'hc91a, 16'hc91b, 16'hc91c, 16'hc91d, 16'hc91e, 16'hc91f 	:	val_out <= 16'h032c;
         16'hc920, 16'hc921, 16'hc922, 16'hc923, 16'hc924, 16'hc925, 16'hc926, 16'hc927 	:	val_out <= 16'h0332;
         16'hc928, 16'hc929, 16'hc92a, 16'hc92b, 16'hc92c, 16'hc92d, 16'hc92e, 16'hc92f 	:	val_out <= 16'h0337;
         16'hc930, 16'hc931, 16'hc932, 16'hc933, 16'hc934, 16'hc935, 16'hc936, 16'hc937 	:	val_out <= 16'h033d;
         16'hc938, 16'hc939, 16'hc93a, 16'hc93b, 16'hc93c, 16'hc93d, 16'hc93e, 16'hc93f 	:	val_out <= 16'h0343;
         16'hc940, 16'hc941, 16'hc942, 16'hc943, 16'hc944, 16'hc945, 16'hc946, 16'hc947 	:	val_out <= 16'h0348;
         16'hc948, 16'hc949, 16'hc94a, 16'hc94b, 16'hc94c, 16'hc94d, 16'hc94e, 16'hc94f 	:	val_out <= 16'h034e;
         16'hc950, 16'hc951, 16'hc952, 16'hc953, 16'hc954, 16'hc955, 16'hc956, 16'hc957 	:	val_out <= 16'h0354;
         16'hc958, 16'hc959, 16'hc95a, 16'hc95b, 16'hc95c, 16'hc95d, 16'hc95e, 16'hc95f 	:	val_out <= 16'h0359;
         16'hc960, 16'hc961, 16'hc962, 16'hc963, 16'hc964, 16'hc965, 16'hc966, 16'hc967 	:	val_out <= 16'h035f;
         16'hc968, 16'hc969, 16'hc96a, 16'hc96b, 16'hc96c, 16'hc96d, 16'hc96e, 16'hc96f 	:	val_out <= 16'h0365;
         16'hc970, 16'hc971, 16'hc972, 16'hc973, 16'hc974, 16'hc975, 16'hc976, 16'hc977 	:	val_out <= 16'h036b;
         16'hc978, 16'hc979, 16'hc97a, 16'hc97b, 16'hc97c, 16'hc97d, 16'hc97e, 16'hc97f 	:	val_out <= 16'h0370;
         16'hc980, 16'hc981, 16'hc982, 16'hc983, 16'hc984, 16'hc985, 16'hc986, 16'hc987 	:	val_out <= 16'h0376;
         16'hc988, 16'hc989, 16'hc98a, 16'hc98b, 16'hc98c, 16'hc98d, 16'hc98e, 16'hc98f 	:	val_out <= 16'h037c;
         16'hc990, 16'hc991, 16'hc992, 16'hc993, 16'hc994, 16'hc995, 16'hc996, 16'hc997 	:	val_out <= 16'h0382;
         16'hc998, 16'hc999, 16'hc99a, 16'hc99b, 16'hc99c, 16'hc99d, 16'hc99e, 16'hc99f 	:	val_out <= 16'h0388;
         16'hc9a0, 16'hc9a1, 16'hc9a2, 16'hc9a3, 16'hc9a4, 16'hc9a5, 16'hc9a6, 16'hc9a7 	:	val_out <= 16'h038e;
         16'hc9a8, 16'hc9a9, 16'hc9aa, 16'hc9ab, 16'hc9ac, 16'hc9ad, 16'hc9ae, 16'hc9af 	:	val_out <= 16'h0393;
         16'hc9b0, 16'hc9b1, 16'hc9b2, 16'hc9b3, 16'hc9b4, 16'hc9b5, 16'hc9b6, 16'hc9b7 	:	val_out <= 16'h0399;
         16'hc9b8, 16'hc9b9, 16'hc9ba, 16'hc9bb, 16'hc9bc, 16'hc9bd, 16'hc9be, 16'hc9bf 	:	val_out <= 16'h039f;
         16'hc9c0, 16'hc9c1, 16'hc9c2, 16'hc9c3, 16'hc9c4, 16'hc9c5, 16'hc9c6, 16'hc9c7 	:	val_out <= 16'h03a5;
         16'hc9c8, 16'hc9c9, 16'hc9ca, 16'hc9cb, 16'hc9cc, 16'hc9cd, 16'hc9ce, 16'hc9cf 	:	val_out <= 16'h03ab;
         16'hc9d0, 16'hc9d1, 16'hc9d2, 16'hc9d3, 16'hc9d4, 16'hc9d5, 16'hc9d6, 16'hc9d7 	:	val_out <= 16'h03b1;
         16'hc9d8, 16'hc9d9, 16'hc9da, 16'hc9db, 16'hc9dc, 16'hc9dd, 16'hc9de, 16'hc9df 	:	val_out <= 16'h03b7;
         16'hc9e0, 16'hc9e1, 16'hc9e2, 16'hc9e3, 16'hc9e4, 16'hc9e5, 16'hc9e6, 16'hc9e7 	:	val_out <= 16'h03bd;
         16'hc9e8, 16'hc9e9, 16'hc9ea, 16'hc9eb, 16'hc9ec, 16'hc9ed, 16'hc9ee, 16'hc9ef 	:	val_out <= 16'h03c3;
         16'hc9f0, 16'hc9f1, 16'hc9f2, 16'hc9f3, 16'hc9f4, 16'hc9f5, 16'hc9f6, 16'hc9f7 	:	val_out <= 16'h03c9;
         16'hc9f8, 16'hc9f9, 16'hc9fa, 16'hc9fb, 16'hc9fc, 16'hc9fd, 16'hc9fe, 16'hc9ff 	:	val_out <= 16'h03cf;
         16'hca00, 16'hca01, 16'hca02, 16'hca03, 16'hca04, 16'hca05, 16'hca06, 16'hca07 	:	val_out <= 16'h03d6;
         16'hca08, 16'hca09, 16'hca0a, 16'hca0b, 16'hca0c, 16'hca0d, 16'hca0e, 16'hca0f 	:	val_out <= 16'h03dc;
         16'hca10, 16'hca11, 16'hca12, 16'hca13, 16'hca14, 16'hca15, 16'hca16, 16'hca17 	:	val_out <= 16'h03e2;
         16'hca18, 16'hca19, 16'hca1a, 16'hca1b, 16'hca1c, 16'hca1d, 16'hca1e, 16'hca1f 	:	val_out <= 16'h03e8;
         16'hca20, 16'hca21, 16'hca22, 16'hca23, 16'hca24, 16'hca25, 16'hca26, 16'hca27 	:	val_out <= 16'h03ee;
         16'hca28, 16'hca29, 16'hca2a, 16'hca2b, 16'hca2c, 16'hca2d, 16'hca2e, 16'hca2f 	:	val_out <= 16'h03f4;
         16'hca30, 16'hca31, 16'hca32, 16'hca33, 16'hca34, 16'hca35, 16'hca36, 16'hca37 	:	val_out <= 16'h03fa;
         16'hca38, 16'hca39, 16'hca3a, 16'hca3b, 16'hca3c, 16'hca3d, 16'hca3e, 16'hca3f 	:	val_out <= 16'h0401;
         16'hca40, 16'hca41, 16'hca42, 16'hca43, 16'hca44, 16'hca45, 16'hca46, 16'hca47 	:	val_out <= 16'h0407;
         16'hca48, 16'hca49, 16'hca4a, 16'hca4b, 16'hca4c, 16'hca4d, 16'hca4e, 16'hca4f 	:	val_out <= 16'h040d;
         16'hca50, 16'hca51, 16'hca52, 16'hca53, 16'hca54, 16'hca55, 16'hca56, 16'hca57 	:	val_out <= 16'h0414;
         16'hca58, 16'hca59, 16'hca5a, 16'hca5b, 16'hca5c, 16'hca5d, 16'hca5e, 16'hca5f 	:	val_out <= 16'h041a;
         16'hca60, 16'hca61, 16'hca62, 16'hca63, 16'hca64, 16'hca65, 16'hca66, 16'hca67 	:	val_out <= 16'h0420;
         16'hca68, 16'hca69, 16'hca6a, 16'hca6b, 16'hca6c, 16'hca6d, 16'hca6e, 16'hca6f 	:	val_out <= 16'h0426;
         16'hca70, 16'hca71, 16'hca72, 16'hca73, 16'hca74, 16'hca75, 16'hca76, 16'hca77 	:	val_out <= 16'h042d;
         16'hca78, 16'hca79, 16'hca7a, 16'hca7b, 16'hca7c, 16'hca7d, 16'hca7e, 16'hca7f 	:	val_out <= 16'h0433;
         16'hca80, 16'hca81, 16'hca82, 16'hca83, 16'hca84, 16'hca85, 16'hca86, 16'hca87 	:	val_out <= 16'h043a;
         16'hca88, 16'hca89, 16'hca8a, 16'hca8b, 16'hca8c, 16'hca8d, 16'hca8e, 16'hca8f 	:	val_out <= 16'h0440;
         16'hca90, 16'hca91, 16'hca92, 16'hca93, 16'hca94, 16'hca95, 16'hca96, 16'hca97 	:	val_out <= 16'h0446;
         16'hca98, 16'hca99, 16'hca9a, 16'hca9b, 16'hca9c, 16'hca9d, 16'hca9e, 16'hca9f 	:	val_out <= 16'h044d;
         16'hcaa0, 16'hcaa1, 16'hcaa2, 16'hcaa3, 16'hcaa4, 16'hcaa5, 16'hcaa6, 16'hcaa7 	:	val_out <= 16'h0453;
         16'hcaa8, 16'hcaa9, 16'hcaaa, 16'hcaab, 16'hcaac, 16'hcaad, 16'hcaae, 16'hcaaf 	:	val_out <= 16'h045a;
         16'hcab0, 16'hcab1, 16'hcab2, 16'hcab3, 16'hcab4, 16'hcab5, 16'hcab6, 16'hcab7 	:	val_out <= 16'h0460;
         16'hcab8, 16'hcab9, 16'hcaba, 16'hcabb, 16'hcabc, 16'hcabd, 16'hcabe, 16'hcabf 	:	val_out <= 16'h0467;
         16'hcac0, 16'hcac1, 16'hcac2, 16'hcac3, 16'hcac4, 16'hcac5, 16'hcac6, 16'hcac7 	:	val_out <= 16'h046d;
         16'hcac8, 16'hcac9, 16'hcaca, 16'hcacb, 16'hcacc, 16'hcacd, 16'hcace, 16'hcacf 	:	val_out <= 16'h0474;
         16'hcad0, 16'hcad1, 16'hcad2, 16'hcad3, 16'hcad4, 16'hcad5, 16'hcad6, 16'hcad7 	:	val_out <= 16'h047b;
         16'hcad8, 16'hcad9, 16'hcada, 16'hcadb, 16'hcadc, 16'hcadd, 16'hcade, 16'hcadf 	:	val_out <= 16'h0481;
         16'hcae0, 16'hcae1, 16'hcae2, 16'hcae3, 16'hcae4, 16'hcae5, 16'hcae6, 16'hcae7 	:	val_out <= 16'h0488;
         16'hcae8, 16'hcae9, 16'hcaea, 16'hcaeb, 16'hcaec, 16'hcaed, 16'hcaee, 16'hcaef 	:	val_out <= 16'h048e;
         16'hcaf0, 16'hcaf1, 16'hcaf2, 16'hcaf3, 16'hcaf4, 16'hcaf5, 16'hcaf6, 16'hcaf7 	:	val_out <= 16'h0495;
         16'hcaf8, 16'hcaf9, 16'hcafa, 16'hcafb, 16'hcafc, 16'hcafd, 16'hcafe, 16'hcaff 	:	val_out <= 16'h049c;
         16'hcb00, 16'hcb01, 16'hcb02, 16'hcb03, 16'hcb04, 16'hcb05, 16'hcb06, 16'hcb07 	:	val_out <= 16'h04a2;
         16'hcb08, 16'hcb09, 16'hcb0a, 16'hcb0b, 16'hcb0c, 16'hcb0d, 16'hcb0e, 16'hcb0f 	:	val_out <= 16'h04a9;
         16'hcb10, 16'hcb11, 16'hcb12, 16'hcb13, 16'hcb14, 16'hcb15, 16'hcb16, 16'hcb17 	:	val_out <= 16'h04b0;
         16'hcb18, 16'hcb19, 16'hcb1a, 16'hcb1b, 16'hcb1c, 16'hcb1d, 16'hcb1e, 16'hcb1f 	:	val_out <= 16'h04b7;
         16'hcb20, 16'hcb21, 16'hcb22, 16'hcb23, 16'hcb24, 16'hcb25, 16'hcb26, 16'hcb27 	:	val_out <= 16'h04bd;
         16'hcb28, 16'hcb29, 16'hcb2a, 16'hcb2b, 16'hcb2c, 16'hcb2d, 16'hcb2e, 16'hcb2f 	:	val_out <= 16'h04c4;
         16'hcb30, 16'hcb31, 16'hcb32, 16'hcb33, 16'hcb34, 16'hcb35, 16'hcb36, 16'hcb37 	:	val_out <= 16'h04cb;
         16'hcb38, 16'hcb39, 16'hcb3a, 16'hcb3b, 16'hcb3c, 16'hcb3d, 16'hcb3e, 16'hcb3f 	:	val_out <= 16'h04d2;
         16'hcb40, 16'hcb41, 16'hcb42, 16'hcb43, 16'hcb44, 16'hcb45, 16'hcb46, 16'hcb47 	:	val_out <= 16'h04d9;
         16'hcb48, 16'hcb49, 16'hcb4a, 16'hcb4b, 16'hcb4c, 16'hcb4d, 16'hcb4e, 16'hcb4f 	:	val_out <= 16'h04e0;
         16'hcb50, 16'hcb51, 16'hcb52, 16'hcb53, 16'hcb54, 16'hcb55, 16'hcb56, 16'hcb57 	:	val_out <= 16'h04e6;
         16'hcb58, 16'hcb59, 16'hcb5a, 16'hcb5b, 16'hcb5c, 16'hcb5d, 16'hcb5e, 16'hcb5f 	:	val_out <= 16'h04ed;
         16'hcb60, 16'hcb61, 16'hcb62, 16'hcb63, 16'hcb64, 16'hcb65, 16'hcb66, 16'hcb67 	:	val_out <= 16'h04f4;
         16'hcb68, 16'hcb69, 16'hcb6a, 16'hcb6b, 16'hcb6c, 16'hcb6d, 16'hcb6e, 16'hcb6f 	:	val_out <= 16'h04fb;
         16'hcb70, 16'hcb71, 16'hcb72, 16'hcb73, 16'hcb74, 16'hcb75, 16'hcb76, 16'hcb77 	:	val_out <= 16'h0502;
         16'hcb78, 16'hcb79, 16'hcb7a, 16'hcb7b, 16'hcb7c, 16'hcb7d, 16'hcb7e, 16'hcb7f 	:	val_out <= 16'h0509;
         16'hcb80, 16'hcb81, 16'hcb82, 16'hcb83, 16'hcb84, 16'hcb85, 16'hcb86, 16'hcb87 	:	val_out <= 16'h0510;
         16'hcb88, 16'hcb89, 16'hcb8a, 16'hcb8b, 16'hcb8c, 16'hcb8d, 16'hcb8e, 16'hcb8f 	:	val_out <= 16'h0517;
         16'hcb90, 16'hcb91, 16'hcb92, 16'hcb93, 16'hcb94, 16'hcb95, 16'hcb96, 16'hcb97 	:	val_out <= 16'h051e;
         16'hcb98, 16'hcb99, 16'hcb9a, 16'hcb9b, 16'hcb9c, 16'hcb9d, 16'hcb9e, 16'hcb9f 	:	val_out <= 16'h0525;
         16'hcba0, 16'hcba1, 16'hcba2, 16'hcba3, 16'hcba4, 16'hcba5, 16'hcba6, 16'hcba7 	:	val_out <= 16'h052c;
         16'hcba8, 16'hcba9, 16'hcbaa, 16'hcbab, 16'hcbac, 16'hcbad, 16'hcbae, 16'hcbaf 	:	val_out <= 16'h0533;
         16'hcbb0, 16'hcbb1, 16'hcbb2, 16'hcbb3, 16'hcbb4, 16'hcbb5, 16'hcbb6, 16'hcbb7 	:	val_out <= 16'h053a;
         16'hcbb8, 16'hcbb9, 16'hcbba, 16'hcbbb, 16'hcbbc, 16'hcbbd, 16'hcbbe, 16'hcbbf 	:	val_out <= 16'h0542;
         16'hcbc0, 16'hcbc1, 16'hcbc2, 16'hcbc3, 16'hcbc4, 16'hcbc5, 16'hcbc6, 16'hcbc7 	:	val_out <= 16'h0549;
         16'hcbc8, 16'hcbc9, 16'hcbca, 16'hcbcb, 16'hcbcc, 16'hcbcd, 16'hcbce, 16'hcbcf 	:	val_out <= 16'h0550;
         16'hcbd0, 16'hcbd1, 16'hcbd2, 16'hcbd3, 16'hcbd4, 16'hcbd5, 16'hcbd6, 16'hcbd7 	:	val_out <= 16'h0557;
         16'hcbd8, 16'hcbd9, 16'hcbda, 16'hcbdb, 16'hcbdc, 16'hcbdd, 16'hcbde, 16'hcbdf 	:	val_out <= 16'h055e;
         16'hcbe0, 16'hcbe1, 16'hcbe2, 16'hcbe3, 16'hcbe4, 16'hcbe5, 16'hcbe6, 16'hcbe7 	:	val_out <= 16'h0565;
         16'hcbe8, 16'hcbe9, 16'hcbea, 16'hcbeb, 16'hcbec, 16'hcbed, 16'hcbee, 16'hcbef 	:	val_out <= 16'h056d;
         16'hcbf0, 16'hcbf1, 16'hcbf2, 16'hcbf3, 16'hcbf4, 16'hcbf5, 16'hcbf6, 16'hcbf7 	:	val_out <= 16'h0574;
         16'hcbf8, 16'hcbf9, 16'hcbfa, 16'hcbfb, 16'hcbfc, 16'hcbfd, 16'hcbfe, 16'hcbff 	:	val_out <= 16'h057b;
         16'hcc00, 16'hcc01, 16'hcc02, 16'hcc03, 16'hcc04, 16'hcc05, 16'hcc06, 16'hcc07 	:	val_out <= 16'h0582;
         16'hcc08, 16'hcc09, 16'hcc0a, 16'hcc0b, 16'hcc0c, 16'hcc0d, 16'hcc0e, 16'hcc0f 	:	val_out <= 16'h058a;
         16'hcc10, 16'hcc11, 16'hcc12, 16'hcc13, 16'hcc14, 16'hcc15, 16'hcc16, 16'hcc17 	:	val_out <= 16'h0591;
         16'hcc18, 16'hcc19, 16'hcc1a, 16'hcc1b, 16'hcc1c, 16'hcc1d, 16'hcc1e, 16'hcc1f 	:	val_out <= 16'h0598;
         16'hcc20, 16'hcc21, 16'hcc22, 16'hcc23, 16'hcc24, 16'hcc25, 16'hcc26, 16'hcc27 	:	val_out <= 16'h05a0;
         16'hcc28, 16'hcc29, 16'hcc2a, 16'hcc2b, 16'hcc2c, 16'hcc2d, 16'hcc2e, 16'hcc2f 	:	val_out <= 16'h05a7;
         16'hcc30, 16'hcc31, 16'hcc32, 16'hcc33, 16'hcc34, 16'hcc35, 16'hcc36, 16'hcc37 	:	val_out <= 16'h05af;
         16'hcc38, 16'hcc39, 16'hcc3a, 16'hcc3b, 16'hcc3c, 16'hcc3d, 16'hcc3e, 16'hcc3f 	:	val_out <= 16'h05b6;
         16'hcc40, 16'hcc41, 16'hcc42, 16'hcc43, 16'hcc44, 16'hcc45, 16'hcc46, 16'hcc47 	:	val_out <= 16'h05bd;
         16'hcc48, 16'hcc49, 16'hcc4a, 16'hcc4b, 16'hcc4c, 16'hcc4d, 16'hcc4e, 16'hcc4f 	:	val_out <= 16'h05c5;
         16'hcc50, 16'hcc51, 16'hcc52, 16'hcc53, 16'hcc54, 16'hcc55, 16'hcc56, 16'hcc57 	:	val_out <= 16'h05cc;
         16'hcc58, 16'hcc59, 16'hcc5a, 16'hcc5b, 16'hcc5c, 16'hcc5d, 16'hcc5e, 16'hcc5f 	:	val_out <= 16'h05d4;
         16'hcc60, 16'hcc61, 16'hcc62, 16'hcc63, 16'hcc64, 16'hcc65, 16'hcc66, 16'hcc67 	:	val_out <= 16'h05db;
         16'hcc68, 16'hcc69, 16'hcc6a, 16'hcc6b, 16'hcc6c, 16'hcc6d, 16'hcc6e, 16'hcc6f 	:	val_out <= 16'h05e3;
         16'hcc70, 16'hcc71, 16'hcc72, 16'hcc73, 16'hcc74, 16'hcc75, 16'hcc76, 16'hcc77 	:	val_out <= 16'h05ea;
         16'hcc78, 16'hcc79, 16'hcc7a, 16'hcc7b, 16'hcc7c, 16'hcc7d, 16'hcc7e, 16'hcc7f 	:	val_out <= 16'h05f2;
         16'hcc80, 16'hcc81, 16'hcc82, 16'hcc83, 16'hcc84, 16'hcc85, 16'hcc86, 16'hcc87 	:	val_out <= 16'h05fa;
         16'hcc88, 16'hcc89, 16'hcc8a, 16'hcc8b, 16'hcc8c, 16'hcc8d, 16'hcc8e, 16'hcc8f 	:	val_out <= 16'h0601;
         16'hcc90, 16'hcc91, 16'hcc92, 16'hcc93, 16'hcc94, 16'hcc95, 16'hcc96, 16'hcc97 	:	val_out <= 16'h0609;
         16'hcc98, 16'hcc99, 16'hcc9a, 16'hcc9b, 16'hcc9c, 16'hcc9d, 16'hcc9e, 16'hcc9f 	:	val_out <= 16'h0610;
         16'hcca0, 16'hcca1, 16'hcca2, 16'hcca3, 16'hcca4, 16'hcca5, 16'hcca6, 16'hcca7 	:	val_out <= 16'h0618;
         16'hcca8, 16'hcca9, 16'hccaa, 16'hccab, 16'hccac, 16'hccad, 16'hccae, 16'hccaf 	:	val_out <= 16'h0620;
         16'hccb0, 16'hccb1, 16'hccb2, 16'hccb3, 16'hccb4, 16'hccb5, 16'hccb6, 16'hccb7 	:	val_out <= 16'h0627;
         16'hccb8, 16'hccb9, 16'hccba, 16'hccbb, 16'hccbc, 16'hccbd, 16'hccbe, 16'hccbf 	:	val_out <= 16'h062f;
         16'hccc0, 16'hccc1, 16'hccc2, 16'hccc3, 16'hccc4, 16'hccc5, 16'hccc6, 16'hccc7 	:	val_out <= 16'h0637;
         16'hccc8, 16'hccc9, 16'hccca, 16'hcccb, 16'hcccc, 16'hcccd, 16'hccce, 16'hcccf 	:	val_out <= 16'h063f;
         16'hccd0, 16'hccd1, 16'hccd2, 16'hccd3, 16'hccd4, 16'hccd5, 16'hccd6, 16'hccd7 	:	val_out <= 16'h0646;
         16'hccd8, 16'hccd9, 16'hccda, 16'hccdb, 16'hccdc, 16'hccdd, 16'hccde, 16'hccdf 	:	val_out <= 16'h064e;
         16'hcce0, 16'hcce1, 16'hcce2, 16'hcce3, 16'hcce4, 16'hcce5, 16'hcce6, 16'hcce7 	:	val_out <= 16'h0656;
         16'hcce8, 16'hcce9, 16'hccea, 16'hcceb, 16'hccec, 16'hcced, 16'hccee, 16'hccef 	:	val_out <= 16'h065e;
         16'hccf0, 16'hccf1, 16'hccf2, 16'hccf3, 16'hccf4, 16'hccf5, 16'hccf6, 16'hccf7 	:	val_out <= 16'h0666;
         16'hccf8, 16'hccf9, 16'hccfa, 16'hccfb, 16'hccfc, 16'hccfd, 16'hccfe, 16'hccff 	:	val_out <= 16'h066d;
         16'hcd00, 16'hcd01, 16'hcd02, 16'hcd03, 16'hcd04, 16'hcd05, 16'hcd06, 16'hcd07 	:	val_out <= 16'h0675;
         16'hcd08, 16'hcd09, 16'hcd0a, 16'hcd0b, 16'hcd0c, 16'hcd0d, 16'hcd0e, 16'hcd0f 	:	val_out <= 16'h067d;
         16'hcd10, 16'hcd11, 16'hcd12, 16'hcd13, 16'hcd14, 16'hcd15, 16'hcd16, 16'hcd17 	:	val_out <= 16'h0685;
         16'hcd18, 16'hcd19, 16'hcd1a, 16'hcd1b, 16'hcd1c, 16'hcd1d, 16'hcd1e, 16'hcd1f 	:	val_out <= 16'h068d;
         16'hcd20, 16'hcd21, 16'hcd22, 16'hcd23, 16'hcd24, 16'hcd25, 16'hcd26, 16'hcd27 	:	val_out <= 16'h0695;
         16'hcd28, 16'hcd29, 16'hcd2a, 16'hcd2b, 16'hcd2c, 16'hcd2d, 16'hcd2e, 16'hcd2f 	:	val_out <= 16'h069d;
         16'hcd30, 16'hcd31, 16'hcd32, 16'hcd33, 16'hcd34, 16'hcd35, 16'hcd36, 16'hcd37 	:	val_out <= 16'h06a5;
         16'hcd38, 16'hcd39, 16'hcd3a, 16'hcd3b, 16'hcd3c, 16'hcd3d, 16'hcd3e, 16'hcd3f 	:	val_out <= 16'h06ad;
         16'hcd40, 16'hcd41, 16'hcd42, 16'hcd43, 16'hcd44, 16'hcd45, 16'hcd46, 16'hcd47 	:	val_out <= 16'h06b5;
         16'hcd48, 16'hcd49, 16'hcd4a, 16'hcd4b, 16'hcd4c, 16'hcd4d, 16'hcd4e, 16'hcd4f 	:	val_out <= 16'h06bd;
         16'hcd50, 16'hcd51, 16'hcd52, 16'hcd53, 16'hcd54, 16'hcd55, 16'hcd56, 16'hcd57 	:	val_out <= 16'h06c5;
         16'hcd58, 16'hcd59, 16'hcd5a, 16'hcd5b, 16'hcd5c, 16'hcd5d, 16'hcd5e, 16'hcd5f 	:	val_out <= 16'h06cd;
         16'hcd60, 16'hcd61, 16'hcd62, 16'hcd63, 16'hcd64, 16'hcd65, 16'hcd66, 16'hcd67 	:	val_out <= 16'h06d5;
         16'hcd68, 16'hcd69, 16'hcd6a, 16'hcd6b, 16'hcd6c, 16'hcd6d, 16'hcd6e, 16'hcd6f 	:	val_out <= 16'h06dd;
         16'hcd70, 16'hcd71, 16'hcd72, 16'hcd73, 16'hcd74, 16'hcd75, 16'hcd76, 16'hcd77 	:	val_out <= 16'h06e6;
         16'hcd78, 16'hcd79, 16'hcd7a, 16'hcd7b, 16'hcd7c, 16'hcd7d, 16'hcd7e, 16'hcd7f 	:	val_out <= 16'h06ee;
         16'hcd80, 16'hcd81, 16'hcd82, 16'hcd83, 16'hcd84, 16'hcd85, 16'hcd86, 16'hcd87 	:	val_out <= 16'h06f6;
         16'hcd88, 16'hcd89, 16'hcd8a, 16'hcd8b, 16'hcd8c, 16'hcd8d, 16'hcd8e, 16'hcd8f 	:	val_out <= 16'h06fe;
         16'hcd90, 16'hcd91, 16'hcd92, 16'hcd93, 16'hcd94, 16'hcd95, 16'hcd96, 16'hcd97 	:	val_out <= 16'h0706;
         16'hcd98, 16'hcd99, 16'hcd9a, 16'hcd9b, 16'hcd9c, 16'hcd9d, 16'hcd9e, 16'hcd9f 	:	val_out <= 16'h070e;
         16'hcda0, 16'hcda1, 16'hcda2, 16'hcda3, 16'hcda4, 16'hcda5, 16'hcda6, 16'hcda7 	:	val_out <= 16'h0717;
         16'hcda8, 16'hcda9, 16'hcdaa, 16'hcdab, 16'hcdac, 16'hcdad, 16'hcdae, 16'hcdaf 	:	val_out <= 16'h071f;
         16'hcdb0, 16'hcdb1, 16'hcdb2, 16'hcdb3, 16'hcdb4, 16'hcdb5, 16'hcdb6, 16'hcdb7 	:	val_out <= 16'h0727;
         16'hcdb8, 16'hcdb9, 16'hcdba, 16'hcdbb, 16'hcdbc, 16'hcdbd, 16'hcdbe, 16'hcdbf 	:	val_out <= 16'h0730;
         16'hcdc0, 16'hcdc1, 16'hcdc2, 16'hcdc3, 16'hcdc4, 16'hcdc5, 16'hcdc6, 16'hcdc7 	:	val_out <= 16'h0738;
         16'hcdc8, 16'hcdc9, 16'hcdca, 16'hcdcb, 16'hcdcc, 16'hcdcd, 16'hcdce, 16'hcdcf 	:	val_out <= 16'h0740;
         16'hcdd0, 16'hcdd1, 16'hcdd2, 16'hcdd3, 16'hcdd4, 16'hcdd5, 16'hcdd6, 16'hcdd7 	:	val_out <= 16'h0749;
         16'hcdd8, 16'hcdd9, 16'hcdda, 16'hcddb, 16'hcddc, 16'hcddd, 16'hcdde, 16'hcddf 	:	val_out <= 16'h0751;
         16'hcde0, 16'hcde1, 16'hcde2, 16'hcde3, 16'hcde4, 16'hcde5, 16'hcde6, 16'hcde7 	:	val_out <= 16'h0759;
         16'hcde8, 16'hcde9, 16'hcdea, 16'hcdeb, 16'hcdec, 16'hcded, 16'hcdee, 16'hcdef 	:	val_out <= 16'h0762;
         16'hcdf0, 16'hcdf1, 16'hcdf2, 16'hcdf3, 16'hcdf4, 16'hcdf5, 16'hcdf6, 16'hcdf7 	:	val_out <= 16'h076a;
         16'hcdf8, 16'hcdf9, 16'hcdfa, 16'hcdfb, 16'hcdfc, 16'hcdfd, 16'hcdfe, 16'hcdff 	:	val_out <= 16'h0773;
         16'hce00, 16'hce01, 16'hce02, 16'hce03, 16'hce04, 16'hce05, 16'hce06, 16'hce07 	:	val_out <= 16'h077b;
         16'hce08, 16'hce09, 16'hce0a, 16'hce0b, 16'hce0c, 16'hce0d, 16'hce0e, 16'hce0f 	:	val_out <= 16'h0783;
         16'hce10, 16'hce11, 16'hce12, 16'hce13, 16'hce14, 16'hce15, 16'hce16, 16'hce17 	:	val_out <= 16'h078c;
         16'hce18, 16'hce19, 16'hce1a, 16'hce1b, 16'hce1c, 16'hce1d, 16'hce1e, 16'hce1f 	:	val_out <= 16'h0794;
         16'hce20, 16'hce21, 16'hce22, 16'hce23, 16'hce24, 16'hce25, 16'hce26, 16'hce27 	:	val_out <= 16'h079d;
         16'hce28, 16'hce29, 16'hce2a, 16'hce2b, 16'hce2c, 16'hce2d, 16'hce2e, 16'hce2f 	:	val_out <= 16'h07a6;
         16'hce30, 16'hce31, 16'hce32, 16'hce33, 16'hce34, 16'hce35, 16'hce36, 16'hce37 	:	val_out <= 16'h07ae;
         16'hce38, 16'hce39, 16'hce3a, 16'hce3b, 16'hce3c, 16'hce3d, 16'hce3e, 16'hce3f 	:	val_out <= 16'h07b7;
         16'hce40, 16'hce41, 16'hce42, 16'hce43, 16'hce44, 16'hce45, 16'hce46, 16'hce47 	:	val_out <= 16'h07bf;
         16'hce48, 16'hce49, 16'hce4a, 16'hce4b, 16'hce4c, 16'hce4d, 16'hce4e, 16'hce4f 	:	val_out <= 16'h07c8;
         16'hce50, 16'hce51, 16'hce52, 16'hce53, 16'hce54, 16'hce55, 16'hce56, 16'hce57 	:	val_out <= 16'h07d1;
         16'hce58, 16'hce59, 16'hce5a, 16'hce5b, 16'hce5c, 16'hce5d, 16'hce5e, 16'hce5f 	:	val_out <= 16'h07d9;
         16'hce60, 16'hce61, 16'hce62, 16'hce63, 16'hce64, 16'hce65, 16'hce66, 16'hce67 	:	val_out <= 16'h07e2;
         16'hce68, 16'hce69, 16'hce6a, 16'hce6b, 16'hce6c, 16'hce6d, 16'hce6e, 16'hce6f 	:	val_out <= 16'h07eb;
         16'hce70, 16'hce71, 16'hce72, 16'hce73, 16'hce74, 16'hce75, 16'hce76, 16'hce77 	:	val_out <= 16'h07f3;
         16'hce78, 16'hce79, 16'hce7a, 16'hce7b, 16'hce7c, 16'hce7d, 16'hce7e, 16'hce7f 	:	val_out <= 16'h07fc;
         16'hce80, 16'hce81, 16'hce82, 16'hce83, 16'hce84, 16'hce85, 16'hce86, 16'hce87 	:	val_out <= 16'h0805;
         16'hce88, 16'hce89, 16'hce8a, 16'hce8b, 16'hce8c, 16'hce8d, 16'hce8e, 16'hce8f 	:	val_out <= 16'h080e;
         16'hce90, 16'hce91, 16'hce92, 16'hce93, 16'hce94, 16'hce95, 16'hce96, 16'hce97 	:	val_out <= 16'h0816;
         16'hce98, 16'hce99, 16'hce9a, 16'hce9b, 16'hce9c, 16'hce9d, 16'hce9e, 16'hce9f 	:	val_out <= 16'h081f;
         16'hcea0, 16'hcea1, 16'hcea2, 16'hcea3, 16'hcea4, 16'hcea5, 16'hcea6, 16'hcea7 	:	val_out <= 16'h0828;
         16'hcea8, 16'hcea9, 16'hceaa, 16'hceab, 16'hceac, 16'hcead, 16'hceae, 16'hceaf 	:	val_out <= 16'h0831;
         16'hceb0, 16'hceb1, 16'hceb2, 16'hceb3, 16'hceb4, 16'hceb5, 16'hceb6, 16'hceb7 	:	val_out <= 16'h083a;
         16'hceb8, 16'hceb9, 16'hceba, 16'hcebb, 16'hcebc, 16'hcebd, 16'hcebe, 16'hcebf 	:	val_out <= 16'h0843;
         16'hcec0, 16'hcec1, 16'hcec2, 16'hcec3, 16'hcec4, 16'hcec5, 16'hcec6, 16'hcec7 	:	val_out <= 16'h084b;
         16'hcec8, 16'hcec9, 16'hceca, 16'hcecb, 16'hcecc, 16'hcecd, 16'hcece, 16'hcecf 	:	val_out <= 16'h0854;
         16'hced0, 16'hced1, 16'hced2, 16'hced3, 16'hced4, 16'hced5, 16'hced6, 16'hced7 	:	val_out <= 16'h085d;
         16'hced8, 16'hced9, 16'hceda, 16'hcedb, 16'hcedc, 16'hcedd, 16'hcede, 16'hcedf 	:	val_out <= 16'h0866;
         16'hcee0, 16'hcee1, 16'hcee2, 16'hcee3, 16'hcee4, 16'hcee5, 16'hcee6, 16'hcee7 	:	val_out <= 16'h086f;
         16'hcee8, 16'hcee9, 16'hceea, 16'hceeb, 16'hceec, 16'hceed, 16'hceee, 16'hceef 	:	val_out <= 16'h0878;
         16'hcef0, 16'hcef1, 16'hcef2, 16'hcef3, 16'hcef4, 16'hcef5, 16'hcef6, 16'hcef7 	:	val_out <= 16'h0881;
         16'hcef8, 16'hcef9, 16'hcefa, 16'hcefb, 16'hcefc, 16'hcefd, 16'hcefe, 16'hceff 	:	val_out <= 16'h088a;
         16'hcf00, 16'hcf01, 16'hcf02, 16'hcf03, 16'hcf04, 16'hcf05, 16'hcf06, 16'hcf07 	:	val_out <= 16'h0893;
         16'hcf08, 16'hcf09, 16'hcf0a, 16'hcf0b, 16'hcf0c, 16'hcf0d, 16'hcf0e, 16'hcf0f 	:	val_out <= 16'h089c;
         16'hcf10, 16'hcf11, 16'hcf12, 16'hcf13, 16'hcf14, 16'hcf15, 16'hcf16, 16'hcf17 	:	val_out <= 16'h08a5;
         16'hcf18, 16'hcf19, 16'hcf1a, 16'hcf1b, 16'hcf1c, 16'hcf1d, 16'hcf1e, 16'hcf1f 	:	val_out <= 16'h08ae;
         16'hcf20, 16'hcf21, 16'hcf22, 16'hcf23, 16'hcf24, 16'hcf25, 16'hcf26, 16'hcf27 	:	val_out <= 16'h08b8;
         16'hcf28, 16'hcf29, 16'hcf2a, 16'hcf2b, 16'hcf2c, 16'hcf2d, 16'hcf2e, 16'hcf2f 	:	val_out <= 16'h08c1;
         16'hcf30, 16'hcf31, 16'hcf32, 16'hcf33, 16'hcf34, 16'hcf35, 16'hcf36, 16'hcf37 	:	val_out <= 16'h08ca;
         16'hcf38, 16'hcf39, 16'hcf3a, 16'hcf3b, 16'hcf3c, 16'hcf3d, 16'hcf3e, 16'hcf3f 	:	val_out <= 16'h08d3;
         16'hcf40, 16'hcf41, 16'hcf42, 16'hcf43, 16'hcf44, 16'hcf45, 16'hcf46, 16'hcf47 	:	val_out <= 16'h08dc;
         16'hcf48, 16'hcf49, 16'hcf4a, 16'hcf4b, 16'hcf4c, 16'hcf4d, 16'hcf4e, 16'hcf4f 	:	val_out <= 16'h08e5;
         16'hcf50, 16'hcf51, 16'hcf52, 16'hcf53, 16'hcf54, 16'hcf55, 16'hcf56, 16'hcf57 	:	val_out <= 16'h08ef;
         16'hcf58, 16'hcf59, 16'hcf5a, 16'hcf5b, 16'hcf5c, 16'hcf5d, 16'hcf5e, 16'hcf5f 	:	val_out <= 16'h08f8;
         16'hcf60, 16'hcf61, 16'hcf62, 16'hcf63, 16'hcf64, 16'hcf65, 16'hcf66, 16'hcf67 	:	val_out <= 16'h0901;
         16'hcf68, 16'hcf69, 16'hcf6a, 16'hcf6b, 16'hcf6c, 16'hcf6d, 16'hcf6e, 16'hcf6f 	:	val_out <= 16'h090a;
         16'hcf70, 16'hcf71, 16'hcf72, 16'hcf73, 16'hcf74, 16'hcf75, 16'hcf76, 16'hcf77 	:	val_out <= 16'h0914;
         16'hcf78, 16'hcf79, 16'hcf7a, 16'hcf7b, 16'hcf7c, 16'hcf7d, 16'hcf7e, 16'hcf7f 	:	val_out <= 16'h091d;
         16'hcf80, 16'hcf81, 16'hcf82, 16'hcf83, 16'hcf84, 16'hcf85, 16'hcf86, 16'hcf87 	:	val_out <= 16'h0926;
         16'hcf88, 16'hcf89, 16'hcf8a, 16'hcf8b, 16'hcf8c, 16'hcf8d, 16'hcf8e, 16'hcf8f 	:	val_out <= 16'h0930;
         16'hcf90, 16'hcf91, 16'hcf92, 16'hcf93, 16'hcf94, 16'hcf95, 16'hcf96, 16'hcf97 	:	val_out <= 16'h0939;
         16'hcf98, 16'hcf99, 16'hcf9a, 16'hcf9b, 16'hcf9c, 16'hcf9d, 16'hcf9e, 16'hcf9f 	:	val_out <= 16'h0942;
         16'hcfa0, 16'hcfa1, 16'hcfa2, 16'hcfa3, 16'hcfa4, 16'hcfa5, 16'hcfa6, 16'hcfa7 	:	val_out <= 16'h094c;
         16'hcfa8, 16'hcfa9, 16'hcfaa, 16'hcfab, 16'hcfac, 16'hcfad, 16'hcfae, 16'hcfaf 	:	val_out <= 16'h0955;
         16'hcfb0, 16'hcfb1, 16'hcfb2, 16'hcfb3, 16'hcfb4, 16'hcfb5, 16'hcfb6, 16'hcfb7 	:	val_out <= 16'h095f;
         16'hcfb8, 16'hcfb9, 16'hcfba, 16'hcfbb, 16'hcfbc, 16'hcfbd, 16'hcfbe, 16'hcfbf 	:	val_out <= 16'h0968;
         16'hcfc0, 16'hcfc1, 16'hcfc2, 16'hcfc3, 16'hcfc4, 16'hcfc5, 16'hcfc6, 16'hcfc7 	:	val_out <= 16'h0971;
         16'hcfc8, 16'hcfc9, 16'hcfca, 16'hcfcb, 16'hcfcc, 16'hcfcd, 16'hcfce, 16'hcfcf 	:	val_out <= 16'h097b;
         16'hcfd0, 16'hcfd1, 16'hcfd2, 16'hcfd3, 16'hcfd4, 16'hcfd5, 16'hcfd6, 16'hcfd7 	:	val_out <= 16'h0984;
         16'hcfd8, 16'hcfd9, 16'hcfda, 16'hcfdb, 16'hcfdc, 16'hcfdd, 16'hcfde, 16'hcfdf 	:	val_out <= 16'h098e;
         16'hcfe0, 16'hcfe1, 16'hcfe2, 16'hcfe3, 16'hcfe4, 16'hcfe5, 16'hcfe6, 16'hcfe7 	:	val_out <= 16'h0997;
         16'hcfe8, 16'hcfe9, 16'hcfea, 16'hcfeb, 16'hcfec, 16'hcfed, 16'hcfee, 16'hcfef 	:	val_out <= 16'h09a1;
         16'hcff0, 16'hcff1, 16'hcff2, 16'hcff3, 16'hcff4, 16'hcff5, 16'hcff6, 16'hcff7 	:	val_out <= 16'h09ab;
         16'hcff8, 16'hcff9, 16'hcffa, 16'hcffb, 16'hcffc, 16'hcffd, 16'hcffe, 16'hcfff 	:	val_out <= 16'h09b4;
         16'hd000, 16'hd001, 16'hd002, 16'hd003, 16'hd004, 16'hd005, 16'hd006, 16'hd007 	:	val_out <= 16'h09be;
         16'hd008, 16'hd009, 16'hd00a, 16'hd00b, 16'hd00c, 16'hd00d, 16'hd00e, 16'hd00f 	:	val_out <= 16'h09c7;
         16'hd010, 16'hd011, 16'hd012, 16'hd013, 16'hd014, 16'hd015, 16'hd016, 16'hd017 	:	val_out <= 16'h09d1;
         16'hd018, 16'hd019, 16'hd01a, 16'hd01b, 16'hd01c, 16'hd01d, 16'hd01e, 16'hd01f 	:	val_out <= 16'h09db;
         16'hd020, 16'hd021, 16'hd022, 16'hd023, 16'hd024, 16'hd025, 16'hd026, 16'hd027 	:	val_out <= 16'h09e4;
         16'hd028, 16'hd029, 16'hd02a, 16'hd02b, 16'hd02c, 16'hd02d, 16'hd02e, 16'hd02f 	:	val_out <= 16'h09ee;
         16'hd030, 16'hd031, 16'hd032, 16'hd033, 16'hd034, 16'hd035, 16'hd036, 16'hd037 	:	val_out <= 16'h09f8;
         16'hd038, 16'hd039, 16'hd03a, 16'hd03b, 16'hd03c, 16'hd03d, 16'hd03e, 16'hd03f 	:	val_out <= 16'h0a02;
         16'hd040, 16'hd041, 16'hd042, 16'hd043, 16'hd044, 16'hd045, 16'hd046, 16'hd047 	:	val_out <= 16'h0a0b;
         16'hd048, 16'hd049, 16'hd04a, 16'hd04b, 16'hd04c, 16'hd04d, 16'hd04e, 16'hd04f 	:	val_out <= 16'h0a15;
         16'hd050, 16'hd051, 16'hd052, 16'hd053, 16'hd054, 16'hd055, 16'hd056, 16'hd057 	:	val_out <= 16'h0a1f;
         16'hd058, 16'hd059, 16'hd05a, 16'hd05b, 16'hd05c, 16'hd05d, 16'hd05e, 16'hd05f 	:	val_out <= 16'h0a29;
         16'hd060, 16'hd061, 16'hd062, 16'hd063, 16'hd064, 16'hd065, 16'hd066, 16'hd067 	:	val_out <= 16'h0a33;
         16'hd068, 16'hd069, 16'hd06a, 16'hd06b, 16'hd06c, 16'hd06d, 16'hd06e, 16'hd06f 	:	val_out <= 16'h0a3c;
         16'hd070, 16'hd071, 16'hd072, 16'hd073, 16'hd074, 16'hd075, 16'hd076, 16'hd077 	:	val_out <= 16'h0a46;
         16'hd078, 16'hd079, 16'hd07a, 16'hd07b, 16'hd07c, 16'hd07d, 16'hd07e, 16'hd07f 	:	val_out <= 16'h0a50;
         16'hd080, 16'hd081, 16'hd082, 16'hd083, 16'hd084, 16'hd085, 16'hd086, 16'hd087 	:	val_out <= 16'h0a5a;
         16'hd088, 16'hd089, 16'hd08a, 16'hd08b, 16'hd08c, 16'hd08d, 16'hd08e, 16'hd08f 	:	val_out <= 16'h0a64;
         16'hd090, 16'hd091, 16'hd092, 16'hd093, 16'hd094, 16'hd095, 16'hd096, 16'hd097 	:	val_out <= 16'h0a6e;
         16'hd098, 16'hd099, 16'hd09a, 16'hd09b, 16'hd09c, 16'hd09d, 16'hd09e, 16'hd09f 	:	val_out <= 16'h0a78;
         16'hd0a0, 16'hd0a1, 16'hd0a2, 16'hd0a3, 16'hd0a4, 16'hd0a5, 16'hd0a6, 16'hd0a7 	:	val_out <= 16'h0a82;
         16'hd0a8, 16'hd0a9, 16'hd0aa, 16'hd0ab, 16'hd0ac, 16'hd0ad, 16'hd0ae, 16'hd0af 	:	val_out <= 16'h0a8c;
         16'hd0b0, 16'hd0b1, 16'hd0b2, 16'hd0b3, 16'hd0b4, 16'hd0b5, 16'hd0b6, 16'hd0b7 	:	val_out <= 16'h0a96;
         16'hd0b8, 16'hd0b9, 16'hd0ba, 16'hd0bb, 16'hd0bc, 16'hd0bd, 16'hd0be, 16'hd0bf 	:	val_out <= 16'h0aa0;
         16'hd0c0, 16'hd0c1, 16'hd0c2, 16'hd0c3, 16'hd0c4, 16'hd0c5, 16'hd0c6, 16'hd0c7 	:	val_out <= 16'h0aaa;
         16'hd0c8, 16'hd0c9, 16'hd0ca, 16'hd0cb, 16'hd0cc, 16'hd0cd, 16'hd0ce, 16'hd0cf 	:	val_out <= 16'h0ab4;
         16'hd0d0, 16'hd0d1, 16'hd0d2, 16'hd0d3, 16'hd0d4, 16'hd0d5, 16'hd0d6, 16'hd0d7 	:	val_out <= 16'h0abe;
         16'hd0d8, 16'hd0d9, 16'hd0da, 16'hd0db, 16'hd0dc, 16'hd0dd, 16'hd0de, 16'hd0df 	:	val_out <= 16'h0ac8;
         16'hd0e0, 16'hd0e1, 16'hd0e2, 16'hd0e3, 16'hd0e4, 16'hd0e5, 16'hd0e6, 16'hd0e7 	:	val_out <= 16'h0ad2;
         16'hd0e8, 16'hd0e9, 16'hd0ea, 16'hd0eb, 16'hd0ec, 16'hd0ed, 16'hd0ee, 16'hd0ef 	:	val_out <= 16'h0adc;
         16'hd0f0, 16'hd0f1, 16'hd0f2, 16'hd0f3, 16'hd0f4, 16'hd0f5, 16'hd0f6, 16'hd0f7 	:	val_out <= 16'h0ae6;
         16'hd0f8, 16'hd0f9, 16'hd0fa, 16'hd0fb, 16'hd0fc, 16'hd0fd, 16'hd0fe, 16'hd0ff 	:	val_out <= 16'h0af0;
         16'hd100, 16'hd101, 16'hd102, 16'hd103, 16'hd104, 16'hd105, 16'hd106, 16'hd107 	:	val_out <= 16'h0afb;
         16'hd108, 16'hd109, 16'hd10a, 16'hd10b, 16'hd10c, 16'hd10d, 16'hd10e, 16'hd10f 	:	val_out <= 16'h0b05;
         16'hd110, 16'hd111, 16'hd112, 16'hd113, 16'hd114, 16'hd115, 16'hd116, 16'hd117 	:	val_out <= 16'h0b0f;
         16'hd118, 16'hd119, 16'hd11a, 16'hd11b, 16'hd11c, 16'hd11d, 16'hd11e, 16'hd11f 	:	val_out <= 16'h0b19;
         16'hd120, 16'hd121, 16'hd122, 16'hd123, 16'hd124, 16'hd125, 16'hd126, 16'hd127 	:	val_out <= 16'h0b24;
         16'hd128, 16'hd129, 16'hd12a, 16'hd12b, 16'hd12c, 16'hd12d, 16'hd12e, 16'hd12f 	:	val_out <= 16'h0b2e;
         16'hd130, 16'hd131, 16'hd132, 16'hd133, 16'hd134, 16'hd135, 16'hd136, 16'hd137 	:	val_out <= 16'h0b38;
         16'hd138, 16'hd139, 16'hd13a, 16'hd13b, 16'hd13c, 16'hd13d, 16'hd13e, 16'hd13f 	:	val_out <= 16'h0b42;
         16'hd140, 16'hd141, 16'hd142, 16'hd143, 16'hd144, 16'hd145, 16'hd146, 16'hd147 	:	val_out <= 16'h0b4d;
         16'hd148, 16'hd149, 16'hd14a, 16'hd14b, 16'hd14c, 16'hd14d, 16'hd14e, 16'hd14f 	:	val_out <= 16'h0b57;
         16'hd150, 16'hd151, 16'hd152, 16'hd153, 16'hd154, 16'hd155, 16'hd156, 16'hd157 	:	val_out <= 16'h0b61;
         16'hd158, 16'hd159, 16'hd15a, 16'hd15b, 16'hd15c, 16'hd15d, 16'hd15e, 16'hd15f 	:	val_out <= 16'h0b6c;
         16'hd160, 16'hd161, 16'hd162, 16'hd163, 16'hd164, 16'hd165, 16'hd166, 16'hd167 	:	val_out <= 16'h0b76;
         16'hd168, 16'hd169, 16'hd16a, 16'hd16b, 16'hd16c, 16'hd16d, 16'hd16e, 16'hd16f 	:	val_out <= 16'h0b81;
         16'hd170, 16'hd171, 16'hd172, 16'hd173, 16'hd174, 16'hd175, 16'hd176, 16'hd177 	:	val_out <= 16'h0b8b;
         16'hd178, 16'hd179, 16'hd17a, 16'hd17b, 16'hd17c, 16'hd17d, 16'hd17e, 16'hd17f 	:	val_out <= 16'h0b95;
         16'hd180, 16'hd181, 16'hd182, 16'hd183, 16'hd184, 16'hd185, 16'hd186, 16'hd187 	:	val_out <= 16'h0ba0;
         16'hd188, 16'hd189, 16'hd18a, 16'hd18b, 16'hd18c, 16'hd18d, 16'hd18e, 16'hd18f 	:	val_out <= 16'h0baa;
         16'hd190, 16'hd191, 16'hd192, 16'hd193, 16'hd194, 16'hd195, 16'hd196, 16'hd197 	:	val_out <= 16'h0bb5;
         16'hd198, 16'hd199, 16'hd19a, 16'hd19b, 16'hd19c, 16'hd19d, 16'hd19e, 16'hd19f 	:	val_out <= 16'h0bbf;
         16'hd1a0, 16'hd1a1, 16'hd1a2, 16'hd1a3, 16'hd1a4, 16'hd1a5, 16'hd1a6, 16'hd1a7 	:	val_out <= 16'h0bca;
         16'hd1a8, 16'hd1a9, 16'hd1aa, 16'hd1ab, 16'hd1ac, 16'hd1ad, 16'hd1ae, 16'hd1af 	:	val_out <= 16'h0bd4;
         16'hd1b0, 16'hd1b1, 16'hd1b2, 16'hd1b3, 16'hd1b4, 16'hd1b5, 16'hd1b6, 16'hd1b7 	:	val_out <= 16'h0bdf;
         16'hd1b8, 16'hd1b9, 16'hd1ba, 16'hd1bb, 16'hd1bc, 16'hd1bd, 16'hd1be, 16'hd1bf 	:	val_out <= 16'h0bea;
         16'hd1c0, 16'hd1c1, 16'hd1c2, 16'hd1c3, 16'hd1c4, 16'hd1c5, 16'hd1c6, 16'hd1c7 	:	val_out <= 16'h0bf4;
         16'hd1c8, 16'hd1c9, 16'hd1ca, 16'hd1cb, 16'hd1cc, 16'hd1cd, 16'hd1ce, 16'hd1cf 	:	val_out <= 16'h0bff;
         16'hd1d0, 16'hd1d1, 16'hd1d2, 16'hd1d3, 16'hd1d4, 16'hd1d5, 16'hd1d6, 16'hd1d7 	:	val_out <= 16'h0c09;
         16'hd1d8, 16'hd1d9, 16'hd1da, 16'hd1db, 16'hd1dc, 16'hd1dd, 16'hd1de, 16'hd1df 	:	val_out <= 16'h0c14;
         16'hd1e0, 16'hd1e1, 16'hd1e2, 16'hd1e3, 16'hd1e4, 16'hd1e5, 16'hd1e6, 16'hd1e7 	:	val_out <= 16'h0c1f;
         16'hd1e8, 16'hd1e9, 16'hd1ea, 16'hd1eb, 16'hd1ec, 16'hd1ed, 16'hd1ee, 16'hd1ef 	:	val_out <= 16'h0c29;
         16'hd1f0, 16'hd1f1, 16'hd1f2, 16'hd1f3, 16'hd1f4, 16'hd1f5, 16'hd1f6, 16'hd1f7 	:	val_out <= 16'h0c34;
         16'hd1f8, 16'hd1f9, 16'hd1fa, 16'hd1fb, 16'hd1fc, 16'hd1fd, 16'hd1fe, 16'hd1ff 	:	val_out <= 16'h0c3f;
         16'hd200, 16'hd201, 16'hd202, 16'hd203, 16'hd204, 16'hd205, 16'hd206, 16'hd207 	:	val_out <= 16'h0c4a;
         16'hd208, 16'hd209, 16'hd20a, 16'hd20b, 16'hd20c, 16'hd20d, 16'hd20e, 16'hd20f 	:	val_out <= 16'h0c54;
         16'hd210, 16'hd211, 16'hd212, 16'hd213, 16'hd214, 16'hd215, 16'hd216, 16'hd217 	:	val_out <= 16'h0c5f;
         16'hd218, 16'hd219, 16'hd21a, 16'hd21b, 16'hd21c, 16'hd21d, 16'hd21e, 16'hd21f 	:	val_out <= 16'h0c6a;
         16'hd220, 16'hd221, 16'hd222, 16'hd223, 16'hd224, 16'hd225, 16'hd226, 16'hd227 	:	val_out <= 16'h0c75;
         16'hd228, 16'hd229, 16'hd22a, 16'hd22b, 16'hd22c, 16'hd22d, 16'hd22e, 16'hd22f 	:	val_out <= 16'h0c80;
         16'hd230, 16'hd231, 16'hd232, 16'hd233, 16'hd234, 16'hd235, 16'hd236, 16'hd237 	:	val_out <= 16'h0c8a;
         16'hd238, 16'hd239, 16'hd23a, 16'hd23b, 16'hd23c, 16'hd23d, 16'hd23e, 16'hd23f 	:	val_out <= 16'h0c95;
         16'hd240, 16'hd241, 16'hd242, 16'hd243, 16'hd244, 16'hd245, 16'hd246, 16'hd247 	:	val_out <= 16'h0ca0;
         16'hd248, 16'hd249, 16'hd24a, 16'hd24b, 16'hd24c, 16'hd24d, 16'hd24e, 16'hd24f 	:	val_out <= 16'h0cab;
         16'hd250, 16'hd251, 16'hd252, 16'hd253, 16'hd254, 16'hd255, 16'hd256, 16'hd257 	:	val_out <= 16'h0cb6;
         16'hd258, 16'hd259, 16'hd25a, 16'hd25b, 16'hd25c, 16'hd25d, 16'hd25e, 16'hd25f 	:	val_out <= 16'h0cc1;
         16'hd260, 16'hd261, 16'hd262, 16'hd263, 16'hd264, 16'hd265, 16'hd266, 16'hd267 	:	val_out <= 16'h0ccc;
         16'hd268, 16'hd269, 16'hd26a, 16'hd26b, 16'hd26c, 16'hd26d, 16'hd26e, 16'hd26f 	:	val_out <= 16'h0cd7;
         16'hd270, 16'hd271, 16'hd272, 16'hd273, 16'hd274, 16'hd275, 16'hd276, 16'hd277 	:	val_out <= 16'h0ce2;
         16'hd278, 16'hd279, 16'hd27a, 16'hd27b, 16'hd27c, 16'hd27d, 16'hd27e, 16'hd27f 	:	val_out <= 16'h0ced;
         16'hd280, 16'hd281, 16'hd282, 16'hd283, 16'hd284, 16'hd285, 16'hd286, 16'hd287 	:	val_out <= 16'h0cf8;
         16'hd288, 16'hd289, 16'hd28a, 16'hd28b, 16'hd28c, 16'hd28d, 16'hd28e, 16'hd28f 	:	val_out <= 16'h0d03;
         16'hd290, 16'hd291, 16'hd292, 16'hd293, 16'hd294, 16'hd295, 16'hd296, 16'hd297 	:	val_out <= 16'h0d0e;
         16'hd298, 16'hd299, 16'hd29a, 16'hd29b, 16'hd29c, 16'hd29d, 16'hd29e, 16'hd29f 	:	val_out <= 16'h0d19;
         16'hd2a0, 16'hd2a1, 16'hd2a2, 16'hd2a3, 16'hd2a4, 16'hd2a5, 16'hd2a6, 16'hd2a7 	:	val_out <= 16'h0d24;
         16'hd2a8, 16'hd2a9, 16'hd2aa, 16'hd2ab, 16'hd2ac, 16'hd2ad, 16'hd2ae, 16'hd2af 	:	val_out <= 16'h0d2f;
         16'hd2b0, 16'hd2b1, 16'hd2b2, 16'hd2b3, 16'hd2b4, 16'hd2b5, 16'hd2b6, 16'hd2b7 	:	val_out <= 16'h0d3a;
         16'hd2b8, 16'hd2b9, 16'hd2ba, 16'hd2bb, 16'hd2bc, 16'hd2bd, 16'hd2be, 16'hd2bf 	:	val_out <= 16'h0d45;
         16'hd2c0, 16'hd2c1, 16'hd2c2, 16'hd2c3, 16'hd2c4, 16'hd2c5, 16'hd2c6, 16'hd2c7 	:	val_out <= 16'h0d50;
         16'hd2c8, 16'hd2c9, 16'hd2ca, 16'hd2cb, 16'hd2cc, 16'hd2cd, 16'hd2ce, 16'hd2cf 	:	val_out <= 16'h0d5c;
         16'hd2d0, 16'hd2d1, 16'hd2d2, 16'hd2d3, 16'hd2d4, 16'hd2d5, 16'hd2d6, 16'hd2d7 	:	val_out <= 16'h0d67;
         16'hd2d8, 16'hd2d9, 16'hd2da, 16'hd2db, 16'hd2dc, 16'hd2dd, 16'hd2de, 16'hd2df 	:	val_out <= 16'h0d72;
         16'hd2e0, 16'hd2e1, 16'hd2e2, 16'hd2e3, 16'hd2e4, 16'hd2e5, 16'hd2e6, 16'hd2e7 	:	val_out <= 16'h0d7d;
         16'hd2e8, 16'hd2e9, 16'hd2ea, 16'hd2eb, 16'hd2ec, 16'hd2ed, 16'hd2ee, 16'hd2ef 	:	val_out <= 16'h0d89;
         16'hd2f0, 16'hd2f1, 16'hd2f2, 16'hd2f3, 16'hd2f4, 16'hd2f5, 16'hd2f6, 16'hd2f7 	:	val_out <= 16'h0d94;
         16'hd2f8, 16'hd2f9, 16'hd2fa, 16'hd2fb, 16'hd2fc, 16'hd2fd, 16'hd2fe, 16'hd2ff 	:	val_out <= 16'h0d9f;
         16'hd300, 16'hd301, 16'hd302, 16'hd303, 16'hd304, 16'hd305, 16'hd306, 16'hd307 	:	val_out <= 16'h0daa;
         16'hd308, 16'hd309, 16'hd30a, 16'hd30b, 16'hd30c, 16'hd30d, 16'hd30e, 16'hd30f 	:	val_out <= 16'h0db6;
         16'hd310, 16'hd311, 16'hd312, 16'hd313, 16'hd314, 16'hd315, 16'hd316, 16'hd317 	:	val_out <= 16'h0dc1;
         16'hd318, 16'hd319, 16'hd31a, 16'hd31b, 16'hd31c, 16'hd31d, 16'hd31e, 16'hd31f 	:	val_out <= 16'h0dcc;
         16'hd320, 16'hd321, 16'hd322, 16'hd323, 16'hd324, 16'hd325, 16'hd326, 16'hd327 	:	val_out <= 16'h0dd8;
         16'hd328, 16'hd329, 16'hd32a, 16'hd32b, 16'hd32c, 16'hd32d, 16'hd32e, 16'hd32f 	:	val_out <= 16'h0de3;
         16'hd330, 16'hd331, 16'hd332, 16'hd333, 16'hd334, 16'hd335, 16'hd336, 16'hd337 	:	val_out <= 16'h0dee;
         16'hd338, 16'hd339, 16'hd33a, 16'hd33b, 16'hd33c, 16'hd33d, 16'hd33e, 16'hd33f 	:	val_out <= 16'h0dfa;
         16'hd340, 16'hd341, 16'hd342, 16'hd343, 16'hd344, 16'hd345, 16'hd346, 16'hd347 	:	val_out <= 16'h0e05;
         16'hd348, 16'hd349, 16'hd34a, 16'hd34b, 16'hd34c, 16'hd34d, 16'hd34e, 16'hd34f 	:	val_out <= 16'h0e11;
         16'hd350, 16'hd351, 16'hd352, 16'hd353, 16'hd354, 16'hd355, 16'hd356, 16'hd357 	:	val_out <= 16'h0e1c;
         16'hd358, 16'hd359, 16'hd35a, 16'hd35b, 16'hd35c, 16'hd35d, 16'hd35e, 16'hd35f 	:	val_out <= 16'h0e28;
         16'hd360, 16'hd361, 16'hd362, 16'hd363, 16'hd364, 16'hd365, 16'hd366, 16'hd367 	:	val_out <= 16'h0e33;
         16'hd368, 16'hd369, 16'hd36a, 16'hd36b, 16'hd36c, 16'hd36d, 16'hd36e, 16'hd36f 	:	val_out <= 16'h0e3f;
         16'hd370, 16'hd371, 16'hd372, 16'hd373, 16'hd374, 16'hd375, 16'hd376, 16'hd377 	:	val_out <= 16'h0e4a;
         16'hd378, 16'hd379, 16'hd37a, 16'hd37b, 16'hd37c, 16'hd37d, 16'hd37e, 16'hd37f 	:	val_out <= 16'h0e56;
         16'hd380, 16'hd381, 16'hd382, 16'hd383, 16'hd384, 16'hd385, 16'hd386, 16'hd387 	:	val_out <= 16'h0e61;
         16'hd388, 16'hd389, 16'hd38a, 16'hd38b, 16'hd38c, 16'hd38d, 16'hd38e, 16'hd38f 	:	val_out <= 16'h0e6d;
         16'hd390, 16'hd391, 16'hd392, 16'hd393, 16'hd394, 16'hd395, 16'hd396, 16'hd397 	:	val_out <= 16'h0e79;
         16'hd398, 16'hd399, 16'hd39a, 16'hd39b, 16'hd39c, 16'hd39d, 16'hd39e, 16'hd39f 	:	val_out <= 16'h0e84;
         16'hd3a0, 16'hd3a1, 16'hd3a2, 16'hd3a3, 16'hd3a4, 16'hd3a5, 16'hd3a6, 16'hd3a7 	:	val_out <= 16'h0e90;
         16'hd3a8, 16'hd3a9, 16'hd3aa, 16'hd3ab, 16'hd3ac, 16'hd3ad, 16'hd3ae, 16'hd3af 	:	val_out <= 16'h0e9b;
         16'hd3b0, 16'hd3b1, 16'hd3b2, 16'hd3b3, 16'hd3b4, 16'hd3b5, 16'hd3b6, 16'hd3b7 	:	val_out <= 16'h0ea7;
         16'hd3b8, 16'hd3b9, 16'hd3ba, 16'hd3bb, 16'hd3bc, 16'hd3bd, 16'hd3be, 16'hd3bf 	:	val_out <= 16'h0eb3;
         16'hd3c0, 16'hd3c1, 16'hd3c2, 16'hd3c3, 16'hd3c4, 16'hd3c5, 16'hd3c6, 16'hd3c7 	:	val_out <= 16'h0ebe;
         16'hd3c8, 16'hd3c9, 16'hd3ca, 16'hd3cb, 16'hd3cc, 16'hd3cd, 16'hd3ce, 16'hd3cf 	:	val_out <= 16'h0eca;
         16'hd3d0, 16'hd3d1, 16'hd3d2, 16'hd3d3, 16'hd3d4, 16'hd3d5, 16'hd3d6, 16'hd3d7 	:	val_out <= 16'h0ed6;
         16'hd3d8, 16'hd3d9, 16'hd3da, 16'hd3db, 16'hd3dc, 16'hd3dd, 16'hd3de, 16'hd3df 	:	val_out <= 16'h0ee2;
         16'hd3e0, 16'hd3e1, 16'hd3e2, 16'hd3e3, 16'hd3e4, 16'hd3e5, 16'hd3e6, 16'hd3e7 	:	val_out <= 16'h0eed;
         16'hd3e8, 16'hd3e9, 16'hd3ea, 16'hd3eb, 16'hd3ec, 16'hd3ed, 16'hd3ee, 16'hd3ef 	:	val_out <= 16'h0ef9;
         16'hd3f0, 16'hd3f1, 16'hd3f2, 16'hd3f3, 16'hd3f4, 16'hd3f5, 16'hd3f6, 16'hd3f7 	:	val_out <= 16'h0f05;
         16'hd3f8, 16'hd3f9, 16'hd3fa, 16'hd3fb, 16'hd3fc, 16'hd3fd, 16'hd3fe, 16'hd3ff 	:	val_out <= 16'h0f11;
         16'hd400, 16'hd401, 16'hd402, 16'hd403, 16'hd404, 16'hd405, 16'hd406, 16'hd407 	:	val_out <= 16'h0f1d;
         16'hd408, 16'hd409, 16'hd40a, 16'hd40b, 16'hd40c, 16'hd40d, 16'hd40e, 16'hd40f 	:	val_out <= 16'h0f29;
         16'hd410, 16'hd411, 16'hd412, 16'hd413, 16'hd414, 16'hd415, 16'hd416, 16'hd417 	:	val_out <= 16'h0f34;
         16'hd418, 16'hd419, 16'hd41a, 16'hd41b, 16'hd41c, 16'hd41d, 16'hd41e, 16'hd41f 	:	val_out <= 16'h0f40;
         16'hd420, 16'hd421, 16'hd422, 16'hd423, 16'hd424, 16'hd425, 16'hd426, 16'hd427 	:	val_out <= 16'h0f4c;
         16'hd428, 16'hd429, 16'hd42a, 16'hd42b, 16'hd42c, 16'hd42d, 16'hd42e, 16'hd42f 	:	val_out <= 16'h0f58;
         16'hd430, 16'hd431, 16'hd432, 16'hd433, 16'hd434, 16'hd435, 16'hd436, 16'hd437 	:	val_out <= 16'h0f64;
         16'hd438, 16'hd439, 16'hd43a, 16'hd43b, 16'hd43c, 16'hd43d, 16'hd43e, 16'hd43f 	:	val_out <= 16'h0f70;
         16'hd440, 16'hd441, 16'hd442, 16'hd443, 16'hd444, 16'hd445, 16'hd446, 16'hd447 	:	val_out <= 16'h0f7c;
         16'hd448, 16'hd449, 16'hd44a, 16'hd44b, 16'hd44c, 16'hd44d, 16'hd44e, 16'hd44f 	:	val_out <= 16'h0f88;
         16'hd450, 16'hd451, 16'hd452, 16'hd453, 16'hd454, 16'hd455, 16'hd456, 16'hd457 	:	val_out <= 16'h0f94;
         16'hd458, 16'hd459, 16'hd45a, 16'hd45b, 16'hd45c, 16'hd45d, 16'hd45e, 16'hd45f 	:	val_out <= 16'h0fa0;
         16'hd460, 16'hd461, 16'hd462, 16'hd463, 16'hd464, 16'hd465, 16'hd466, 16'hd467 	:	val_out <= 16'h0fac;
         16'hd468, 16'hd469, 16'hd46a, 16'hd46b, 16'hd46c, 16'hd46d, 16'hd46e, 16'hd46f 	:	val_out <= 16'h0fb8;
         16'hd470, 16'hd471, 16'hd472, 16'hd473, 16'hd474, 16'hd475, 16'hd476, 16'hd477 	:	val_out <= 16'h0fc4;
         16'hd478, 16'hd479, 16'hd47a, 16'hd47b, 16'hd47c, 16'hd47d, 16'hd47e, 16'hd47f 	:	val_out <= 16'h0fd0;
         16'hd480, 16'hd481, 16'hd482, 16'hd483, 16'hd484, 16'hd485, 16'hd486, 16'hd487 	:	val_out <= 16'h0fdc;
         16'hd488, 16'hd489, 16'hd48a, 16'hd48b, 16'hd48c, 16'hd48d, 16'hd48e, 16'hd48f 	:	val_out <= 16'h0fe9;
         16'hd490, 16'hd491, 16'hd492, 16'hd493, 16'hd494, 16'hd495, 16'hd496, 16'hd497 	:	val_out <= 16'h0ff5;
         16'hd498, 16'hd499, 16'hd49a, 16'hd49b, 16'hd49c, 16'hd49d, 16'hd49e, 16'hd49f 	:	val_out <= 16'h1001;
         16'hd4a0, 16'hd4a1, 16'hd4a2, 16'hd4a3, 16'hd4a4, 16'hd4a5, 16'hd4a6, 16'hd4a7 	:	val_out <= 16'h100d;
         16'hd4a8, 16'hd4a9, 16'hd4aa, 16'hd4ab, 16'hd4ac, 16'hd4ad, 16'hd4ae, 16'hd4af 	:	val_out <= 16'h1019;
         16'hd4b0, 16'hd4b1, 16'hd4b2, 16'hd4b3, 16'hd4b4, 16'hd4b5, 16'hd4b6, 16'hd4b7 	:	val_out <= 16'h1025;
         16'hd4b8, 16'hd4b9, 16'hd4ba, 16'hd4bb, 16'hd4bc, 16'hd4bd, 16'hd4be, 16'hd4bf 	:	val_out <= 16'h1032;
         16'hd4c0, 16'hd4c1, 16'hd4c2, 16'hd4c3, 16'hd4c4, 16'hd4c5, 16'hd4c6, 16'hd4c7 	:	val_out <= 16'h103e;
         16'hd4c8, 16'hd4c9, 16'hd4ca, 16'hd4cb, 16'hd4cc, 16'hd4cd, 16'hd4ce, 16'hd4cf 	:	val_out <= 16'h104a;
         16'hd4d0, 16'hd4d1, 16'hd4d2, 16'hd4d3, 16'hd4d4, 16'hd4d5, 16'hd4d6, 16'hd4d7 	:	val_out <= 16'h1056;
         16'hd4d8, 16'hd4d9, 16'hd4da, 16'hd4db, 16'hd4dc, 16'hd4dd, 16'hd4de, 16'hd4df 	:	val_out <= 16'h1063;
         16'hd4e0, 16'hd4e1, 16'hd4e2, 16'hd4e3, 16'hd4e4, 16'hd4e5, 16'hd4e6, 16'hd4e7 	:	val_out <= 16'h106f;
         16'hd4e8, 16'hd4e9, 16'hd4ea, 16'hd4eb, 16'hd4ec, 16'hd4ed, 16'hd4ee, 16'hd4ef 	:	val_out <= 16'h107b;
         16'hd4f0, 16'hd4f1, 16'hd4f2, 16'hd4f3, 16'hd4f4, 16'hd4f5, 16'hd4f6, 16'hd4f7 	:	val_out <= 16'h1088;
         16'hd4f8, 16'hd4f9, 16'hd4fa, 16'hd4fb, 16'hd4fc, 16'hd4fd, 16'hd4fe, 16'hd4ff 	:	val_out <= 16'h1094;
         16'hd500, 16'hd501, 16'hd502, 16'hd503, 16'hd504, 16'hd505, 16'hd506, 16'hd507 	:	val_out <= 16'h10a0;
         16'hd508, 16'hd509, 16'hd50a, 16'hd50b, 16'hd50c, 16'hd50d, 16'hd50e, 16'hd50f 	:	val_out <= 16'h10ad;
         16'hd510, 16'hd511, 16'hd512, 16'hd513, 16'hd514, 16'hd515, 16'hd516, 16'hd517 	:	val_out <= 16'h10b9;
         16'hd518, 16'hd519, 16'hd51a, 16'hd51b, 16'hd51c, 16'hd51d, 16'hd51e, 16'hd51f 	:	val_out <= 16'h10c6;
         16'hd520, 16'hd521, 16'hd522, 16'hd523, 16'hd524, 16'hd525, 16'hd526, 16'hd527 	:	val_out <= 16'h10d2;
         16'hd528, 16'hd529, 16'hd52a, 16'hd52b, 16'hd52c, 16'hd52d, 16'hd52e, 16'hd52f 	:	val_out <= 16'h10df;
         16'hd530, 16'hd531, 16'hd532, 16'hd533, 16'hd534, 16'hd535, 16'hd536, 16'hd537 	:	val_out <= 16'h10eb;
         16'hd538, 16'hd539, 16'hd53a, 16'hd53b, 16'hd53c, 16'hd53d, 16'hd53e, 16'hd53f 	:	val_out <= 16'h10f8;
         16'hd540, 16'hd541, 16'hd542, 16'hd543, 16'hd544, 16'hd545, 16'hd546, 16'hd547 	:	val_out <= 16'h1104;
         16'hd548, 16'hd549, 16'hd54a, 16'hd54b, 16'hd54c, 16'hd54d, 16'hd54e, 16'hd54f 	:	val_out <= 16'h1111;
         16'hd550, 16'hd551, 16'hd552, 16'hd553, 16'hd554, 16'hd555, 16'hd556, 16'hd557 	:	val_out <= 16'h111d;
         16'hd558, 16'hd559, 16'hd55a, 16'hd55b, 16'hd55c, 16'hd55d, 16'hd55e, 16'hd55f 	:	val_out <= 16'h112a;
         16'hd560, 16'hd561, 16'hd562, 16'hd563, 16'hd564, 16'hd565, 16'hd566, 16'hd567 	:	val_out <= 16'h1136;
         16'hd568, 16'hd569, 16'hd56a, 16'hd56b, 16'hd56c, 16'hd56d, 16'hd56e, 16'hd56f 	:	val_out <= 16'h1143;
         16'hd570, 16'hd571, 16'hd572, 16'hd573, 16'hd574, 16'hd575, 16'hd576, 16'hd577 	:	val_out <= 16'h1150;
         16'hd578, 16'hd579, 16'hd57a, 16'hd57b, 16'hd57c, 16'hd57d, 16'hd57e, 16'hd57f 	:	val_out <= 16'h115c;
         16'hd580, 16'hd581, 16'hd582, 16'hd583, 16'hd584, 16'hd585, 16'hd586, 16'hd587 	:	val_out <= 16'h1169;
         16'hd588, 16'hd589, 16'hd58a, 16'hd58b, 16'hd58c, 16'hd58d, 16'hd58e, 16'hd58f 	:	val_out <= 16'h1176;
         16'hd590, 16'hd591, 16'hd592, 16'hd593, 16'hd594, 16'hd595, 16'hd596, 16'hd597 	:	val_out <= 16'h1182;
         16'hd598, 16'hd599, 16'hd59a, 16'hd59b, 16'hd59c, 16'hd59d, 16'hd59e, 16'hd59f 	:	val_out <= 16'h118f;
         16'hd5a0, 16'hd5a1, 16'hd5a2, 16'hd5a3, 16'hd5a4, 16'hd5a5, 16'hd5a6, 16'hd5a7 	:	val_out <= 16'h119c;
         16'hd5a8, 16'hd5a9, 16'hd5aa, 16'hd5ab, 16'hd5ac, 16'hd5ad, 16'hd5ae, 16'hd5af 	:	val_out <= 16'h11a8;
         16'hd5b0, 16'hd5b1, 16'hd5b2, 16'hd5b3, 16'hd5b4, 16'hd5b5, 16'hd5b6, 16'hd5b7 	:	val_out <= 16'h11b5;
         16'hd5b8, 16'hd5b9, 16'hd5ba, 16'hd5bb, 16'hd5bc, 16'hd5bd, 16'hd5be, 16'hd5bf 	:	val_out <= 16'h11c2;
         16'hd5c0, 16'hd5c1, 16'hd5c2, 16'hd5c3, 16'hd5c4, 16'hd5c5, 16'hd5c6, 16'hd5c7 	:	val_out <= 16'h11cf;
         16'hd5c8, 16'hd5c9, 16'hd5ca, 16'hd5cb, 16'hd5cc, 16'hd5cd, 16'hd5ce, 16'hd5cf 	:	val_out <= 16'h11db;
         16'hd5d0, 16'hd5d1, 16'hd5d2, 16'hd5d3, 16'hd5d4, 16'hd5d5, 16'hd5d6, 16'hd5d7 	:	val_out <= 16'h11e8;
         16'hd5d8, 16'hd5d9, 16'hd5da, 16'hd5db, 16'hd5dc, 16'hd5dd, 16'hd5de, 16'hd5df 	:	val_out <= 16'h11f5;
         16'hd5e0, 16'hd5e1, 16'hd5e2, 16'hd5e3, 16'hd5e4, 16'hd5e5, 16'hd5e6, 16'hd5e7 	:	val_out <= 16'h1202;
         16'hd5e8, 16'hd5e9, 16'hd5ea, 16'hd5eb, 16'hd5ec, 16'hd5ed, 16'hd5ee, 16'hd5ef 	:	val_out <= 16'h120f;
         16'hd5f0, 16'hd5f1, 16'hd5f2, 16'hd5f3, 16'hd5f4, 16'hd5f5, 16'hd5f6, 16'hd5f7 	:	val_out <= 16'h121c;
         16'hd5f8, 16'hd5f9, 16'hd5fa, 16'hd5fb, 16'hd5fc, 16'hd5fd, 16'hd5fe, 16'hd5ff 	:	val_out <= 16'h1229;
         16'hd600, 16'hd601, 16'hd602, 16'hd603, 16'hd604, 16'hd605, 16'hd606, 16'hd607 	:	val_out <= 16'h1235;
         16'hd608, 16'hd609, 16'hd60a, 16'hd60b, 16'hd60c, 16'hd60d, 16'hd60e, 16'hd60f 	:	val_out <= 16'h1242;
         16'hd610, 16'hd611, 16'hd612, 16'hd613, 16'hd614, 16'hd615, 16'hd616, 16'hd617 	:	val_out <= 16'h124f;
         16'hd618, 16'hd619, 16'hd61a, 16'hd61b, 16'hd61c, 16'hd61d, 16'hd61e, 16'hd61f 	:	val_out <= 16'h125c;
         16'hd620, 16'hd621, 16'hd622, 16'hd623, 16'hd624, 16'hd625, 16'hd626, 16'hd627 	:	val_out <= 16'h1269;
         16'hd628, 16'hd629, 16'hd62a, 16'hd62b, 16'hd62c, 16'hd62d, 16'hd62e, 16'hd62f 	:	val_out <= 16'h1276;
         16'hd630, 16'hd631, 16'hd632, 16'hd633, 16'hd634, 16'hd635, 16'hd636, 16'hd637 	:	val_out <= 16'h1283;
         16'hd638, 16'hd639, 16'hd63a, 16'hd63b, 16'hd63c, 16'hd63d, 16'hd63e, 16'hd63f 	:	val_out <= 16'h1290;
         16'hd640, 16'hd641, 16'hd642, 16'hd643, 16'hd644, 16'hd645, 16'hd646, 16'hd647 	:	val_out <= 16'h129d;
         16'hd648, 16'hd649, 16'hd64a, 16'hd64b, 16'hd64c, 16'hd64d, 16'hd64e, 16'hd64f 	:	val_out <= 16'h12aa;
         16'hd650, 16'hd651, 16'hd652, 16'hd653, 16'hd654, 16'hd655, 16'hd656, 16'hd657 	:	val_out <= 16'h12b7;
         16'hd658, 16'hd659, 16'hd65a, 16'hd65b, 16'hd65c, 16'hd65d, 16'hd65e, 16'hd65f 	:	val_out <= 16'h12c5;
         16'hd660, 16'hd661, 16'hd662, 16'hd663, 16'hd664, 16'hd665, 16'hd666, 16'hd667 	:	val_out <= 16'h12d2;
         16'hd668, 16'hd669, 16'hd66a, 16'hd66b, 16'hd66c, 16'hd66d, 16'hd66e, 16'hd66f 	:	val_out <= 16'h12df;
         16'hd670, 16'hd671, 16'hd672, 16'hd673, 16'hd674, 16'hd675, 16'hd676, 16'hd677 	:	val_out <= 16'h12ec;
         16'hd678, 16'hd679, 16'hd67a, 16'hd67b, 16'hd67c, 16'hd67d, 16'hd67e, 16'hd67f 	:	val_out <= 16'h12f9;
         16'hd680, 16'hd681, 16'hd682, 16'hd683, 16'hd684, 16'hd685, 16'hd686, 16'hd687 	:	val_out <= 16'h1306;
         16'hd688, 16'hd689, 16'hd68a, 16'hd68b, 16'hd68c, 16'hd68d, 16'hd68e, 16'hd68f 	:	val_out <= 16'h1313;
         16'hd690, 16'hd691, 16'hd692, 16'hd693, 16'hd694, 16'hd695, 16'hd696, 16'hd697 	:	val_out <= 16'h1321;
         16'hd698, 16'hd699, 16'hd69a, 16'hd69b, 16'hd69c, 16'hd69d, 16'hd69e, 16'hd69f 	:	val_out <= 16'h132e;
         16'hd6a0, 16'hd6a1, 16'hd6a2, 16'hd6a3, 16'hd6a4, 16'hd6a5, 16'hd6a6, 16'hd6a7 	:	val_out <= 16'h133b;
         16'hd6a8, 16'hd6a9, 16'hd6aa, 16'hd6ab, 16'hd6ac, 16'hd6ad, 16'hd6ae, 16'hd6af 	:	val_out <= 16'h1348;
         16'hd6b0, 16'hd6b1, 16'hd6b2, 16'hd6b3, 16'hd6b4, 16'hd6b5, 16'hd6b6, 16'hd6b7 	:	val_out <= 16'h1356;
         16'hd6b8, 16'hd6b9, 16'hd6ba, 16'hd6bb, 16'hd6bc, 16'hd6bd, 16'hd6be, 16'hd6bf 	:	val_out <= 16'h1363;
         16'hd6c0, 16'hd6c1, 16'hd6c2, 16'hd6c3, 16'hd6c4, 16'hd6c5, 16'hd6c6, 16'hd6c7 	:	val_out <= 16'h1370;
         16'hd6c8, 16'hd6c9, 16'hd6ca, 16'hd6cb, 16'hd6cc, 16'hd6cd, 16'hd6ce, 16'hd6cf 	:	val_out <= 16'h137e;
         16'hd6d0, 16'hd6d1, 16'hd6d2, 16'hd6d3, 16'hd6d4, 16'hd6d5, 16'hd6d6, 16'hd6d7 	:	val_out <= 16'h138b;
         16'hd6d8, 16'hd6d9, 16'hd6da, 16'hd6db, 16'hd6dc, 16'hd6dd, 16'hd6de, 16'hd6df 	:	val_out <= 16'h1398;
         16'hd6e0, 16'hd6e1, 16'hd6e2, 16'hd6e3, 16'hd6e4, 16'hd6e5, 16'hd6e6, 16'hd6e7 	:	val_out <= 16'h13a6;
         16'hd6e8, 16'hd6e9, 16'hd6ea, 16'hd6eb, 16'hd6ec, 16'hd6ed, 16'hd6ee, 16'hd6ef 	:	val_out <= 16'h13b3;
         16'hd6f0, 16'hd6f1, 16'hd6f2, 16'hd6f3, 16'hd6f4, 16'hd6f5, 16'hd6f6, 16'hd6f7 	:	val_out <= 16'h13c0;
         16'hd6f8, 16'hd6f9, 16'hd6fa, 16'hd6fb, 16'hd6fc, 16'hd6fd, 16'hd6fe, 16'hd6ff 	:	val_out <= 16'h13ce;
         16'hd700, 16'hd701, 16'hd702, 16'hd703, 16'hd704, 16'hd705, 16'hd706, 16'hd707 	:	val_out <= 16'h13db;
         16'hd708, 16'hd709, 16'hd70a, 16'hd70b, 16'hd70c, 16'hd70d, 16'hd70e, 16'hd70f 	:	val_out <= 16'h13e9;
         16'hd710, 16'hd711, 16'hd712, 16'hd713, 16'hd714, 16'hd715, 16'hd716, 16'hd717 	:	val_out <= 16'h13f6;
         16'hd718, 16'hd719, 16'hd71a, 16'hd71b, 16'hd71c, 16'hd71d, 16'hd71e, 16'hd71f 	:	val_out <= 16'h1404;
         16'hd720, 16'hd721, 16'hd722, 16'hd723, 16'hd724, 16'hd725, 16'hd726, 16'hd727 	:	val_out <= 16'h1411;
         16'hd728, 16'hd729, 16'hd72a, 16'hd72b, 16'hd72c, 16'hd72d, 16'hd72e, 16'hd72f 	:	val_out <= 16'h141f;
         16'hd730, 16'hd731, 16'hd732, 16'hd733, 16'hd734, 16'hd735, 16'hd736, 16'hd737 	:	val_out <= 16'h142c;
         16'hd738, 16'hd739, 16'hd73a, 16'hd73b, 16'hd73c, 16'hd73d, 16'hd73e, 16'hd73f 	:	val_out <= 16'h143a;
         16'hd740, 16'hd741, 16'hd742, 16'hd743, 16'hd744, 16'hd745, 16'hd746, 16'hd747 	:	val_out <= 16'h1447;
         16'hd748, 16'hd749, 16'hd74a, 16'hd74b, 16'hd74c, 16'hd74d, 16'hd74e, 16'hd74f 	:	val_out <= 16'h1455;
         16'hd750, 16'hd751, 16'hd752, 16'hd753, 16'hd754, 16'hd755, 16'hd756, 16'hd757 	:	val_out <= 16'h1463;
         16'hd758, 16'hd759, 16'hd75a, 16'hd75b, 16'hd75c, 16'hd75d, 16'hd75e, 16'hd75f 	:	val_out <= 16'h1470;
         16'hd760, 16'hd761, 16'hd762, 16'hd763, 16'hd764, 16'hd765, 16'hd766, 16'hd767 	:	val_out <= 16'h147e;
         16'hd768, 16'hd769, 16'hd76a, 16'hd76b, 16'hd76c, 16'hd76d, 16'hd76e, 16'hd76f 	:	val_out <= 16'h148c;
         16'hd770, 16'hd771, 16'hd772, 16'hd773, 16'hd774, 16'hd775, 16'hd776, 16'hd777 	:	val_out <= 16'h1499;
         16'hd778, 16'hd779, 16'hd77a, 16'hd77b, 16'hd77c, 16'hd77d, 16'hd77e, 16'hd77f 	:	val_out <= 16'h14a7;
         16'hd780, 16'hd781, 16'hd782, 16'hd783, 16'hd784, 16'hd785, 16'hd786, 16'hd787 	:	val_out <= 16'h14b5;
         16'hd788, 16'hd789, 16'hd78a, 16'hd78b, 16'hd78c, 16'hd78d, 16'hd78e, 16'hd78f 	:	val_out <= 16'h14c2;
         16'hd790, 16'hd791, 16'hd792, 16'hd793, 16'hd794, 16'hd795, 16'hd796, 16'hd797 	:	val_out <= 16'h14d0;
         16'hd798, 16'hd799, 16'hd79a, 16'hd79b, 16'hd79c, 16'hd79d, 16'hd79e, 16'hd79f 	:	val_out <= 16'h14de;
         16'hd7a0, 16'hd7a1, 16'hd7a2, 16'hd7a3, 16'hd7a4, 16'hd7a5, 16'hd7a6, 16'hd7a7 	:	val_out <= 16'h14ec;
         16'hd7a8, 16'hd7a9, 16'hd7aa, 16'hd7ab, 16'hd7ac, 16'hd7ad, 16'hd7ae, 16'hd7af 	:	val_out <= 16'h14f9;
         16'hd7b0, 16'hd7b1, 16'hd7b2, 16'hd7b3, 16'hd7b4, 16'hd7b5, 16'hd7b6, 16'hd7b7 	:	val_out <= 16'h1507;
         16'hd7b8, 16'hd7b9, 16'hd7ba, 16'hd7bb, 16'hd7bc, 16'hd7bd, 16'hd7be, 16'hd7bf 	:	val_out <= 16'h1515;
         16'hd7c0, 16'hd7c1, 16'hd7c2, 16'hd7c3, 16'hd7c4, 16'hd7c5, 16'hd7c6, 16'hd7c7 	:	val_out <= 16'h1523;
         16'hd7c8, 16'hd7c9, 16'hd7ca, 16'hd7cb, 16'hd7cc, 16'hd7cd, 16'hd7ce, 16'hd7cf 	:	val_out <= 16'h1531;
         16'hd7d0, 16'hd7d1, 16'hd7d2, 16'hd7d3, 16'hd7d4, 16'hd7d5, 16'hd7d6, 16'hd7d7 	:	val_out <= 16'h153e;
         16'hd7d8, 16'hd7d9, 16'hd7da, 16'hd7db, 16'hd7dc, 16'hd7dd, 16'hd7de, 16'hd7df 	:	val_out <= 16'h154c;
         16'hd7e0, 16'hd7e1, 16'hd7e2, 16'hd7e3, 16'hd7e4, 16'hd7e5, 16'hd7e6, 16'hd7e7 	:	val_out <= 16'h155a;
         16'hd7e8, 16'hd7e9, 16'hd7ea, 16'hd7eb, 16'hd7ec, 16'hd7ed, 16'hd7ee, 16'hd7ef 	:	val_out <= 16'h1568;
         16'hd7f0, 16'hd7f1, 16'hd7f2, 16'hd7f3, 16'hd7f4, 16'hd7f5, 16'hd7f6, 16'hd7f7 	:	val_out <= 16'h1576;
         16'hd7f8, 16'hd7f9, 16'hd7fa, 16'hd7fb, 16'hd7fc, 16'hd7fd, 16'hd7fe, 16'hd7ff 	:	val_out <= 16'h1584;
         16'hd800, 16'hd801, 16'hd802, 16'hd803, 16'hd804, 16'hd805, 16'hd806, 16'hd807 	:	val_out <= 16'h1592;
         16'hd808, 16'hd809, 16'hd80a, 16'hd80b, 16'hd80c, 16'hd80d, 16'hd80e, 16'hd80f 	:	val_out <= 16'h15a0;
         16'hd810, 16'hd811, 16'hd812, 16'hd813, 16'hd814, 16'hd815, 16'hd816, 16'hd817 	:	val_out <= 16'h15ae;
         16'hd818, 16'hd819, 16'hd81a, 16'hd81b, 16'hd81c, 16'hd81d, 16'hd81e, 16'hd81f 	:	val_out <= 16'h15bc;
         16'hd820, 16'hd821, 16'hd822, 16'hd823, 16'hd824, 16'hd825, 16'hd826, 16'hd827 	:	val_out <= 16'h15ca;
         16'hd828, 16'hd829, 16'hd82a, 16'hd82b, 16'hd82c, 16'hd82d, 16'hd82e, 16'hd82f 	:	val_out <= 16'h15d8;
         16'hd830, 16'hd831, 16'hd832, 16'hd833, 16'hd834, 16'hd835, 16'hd836, 16'hd837 	:	val_out <= 16'h15e6;
         16'hd838, 16'hd839, 16'hd83a, 16'hd83b, 16'hd83c, 16'hd83d, 16'hd83e, 16'hd83f 	:	val_out <= 16'h15f4;
         16'hd840, 16'hd841, 16'hd842, 16'hd843, 16'hd844, 16'hd845, 16'hd846, 16'hd847 	:	val_out <= 16'h1602;
         16'hd848, 16'hd849, 16'hd84a, 16'hd84b, 16'hd84c, 16'hd84d, 16'hd84e, 16'hd84f 	:	val_out <= 16'h1610;
         16'hd850, 16'hd851, 16'hd852, 16'hd853, 16'hd854, 16'hd855, 16'hd856, 16'hd857 	:	val_out <= 16'h161e;
         16'hd858, 16'hd859, 16'hd85a, 16'hd85b, 16'hd85c, 16'hd85d, 16'hd85e, 16'hd85f 	:	val_out <= 16'h162c;
         16'hd860, 16'hd861, 16'hd862, 16'hd863, 16'hd864, 16'hd865, 16'hd866, 16'hd867 	:	val_out <= 16'h163b;
         16'hd868, 16'hd869, 16'hd86a, 16'hd86b, 16'hd86c, 16'hd86d, 16'hd86e, 16'hd86f 	:	val_out <= 16'h1649;
         16'hd870, 16'hd871, 16'hd872, 16'hd873, 16'hd874, 16'hd875, 16'hd876, 16'hd877 	:	val_out <= 16'h1657;
         16'hd878, 16'hd879, 16'hd87a, 16'hd87b, 16'hd87c, 16'hd87d, 16'hd87e, 16'hd87f 	:	val_out <= 16'h1665;
         16'hd880, 16'hd881, 16'hd882, 16'hd883, 16'hd884, 16'hd885, 16'hd886, 16'hd887 	:	val_out <= 16'h1673;
         16'hd888, 16'hd889, 16'hd88a, 16'hd88b, 16'hd88c, 16'hd88d, 16'hd88e, 16'hd88f 	:	val_out <= 16'h1682;
         16'hd890, 16'hd891, 16'hd892, 16'hd893, 16'hd894, 16'hd895, 16'hd896, 16'hd897 	:	val_out <= 16'h1690;
         16'hd898, 16'hd899, 16'hd89a, 16'hd89b, 16'hd89c, 16'hd89d, 16'hd89e, 16'hd89f 	:	val_out <= 16'h169e;
         16'hd8a0, 16'hd8a1, 16'hd8a2, 16'hd8a3, 16'hd8a4, 16'hd8a5, 16'hd8a6, 16'hd8a7 	:	val_out <= 16'h16ac;
         16'hd8a8, 16'hd8a9, 16'hd8aa, 16'hd8ab, 16'hd8ac, 16'hd8ad, 16'hd8ae, 16'hd8af 	:	val_out <= 16'h16bb;
         16'hd8b0, 16'hd8b1, 16'hd8b2, 16'hd8b3, 16'hd8b4, 16'hd8b5, 16'hd8b6, 16'hd8b7 	:	val_out <= 16'h16c9;
         16'hd8b8, 16'hd8b9, 16'hd8ba, 16'hd8bb, 16'hd8bc, 16'hd8bd, 16'hd8be, 16'hd8bf 	:	val_out <= 16'h16d7;
         16'hd8c0, 16'hd8c1, 16'hd8c2, 16'hd8c3, 16'hd8c4, 16'hd8c5, 16'hd8c6, 16'hd8c7 	:	val_out <= 16'h16e6;
         16'hd8c8, 16'hd8c9, 16'hd8ca, 16'hd8cb, 16'hd8cc, 16'hd8cd, 16'hd8ce, 16'hd8cf 	:	val_out <= 16'h16f4;
         16'hd8d0, 16'hd8d1, 16'hd8d2, 16'hd8d3, 16'hd8d4, 16'hd8d5, 16'hd8d6, 16'hd8d7 	:	val_out <= 16'h1702;
         16'hd8d8, 16'hd8d9, 16'hd8da, 16'hd8db, 16'hd8dc, 16'hd8dd, 16'hd8de, 16'hd8df 	:	val_out <= 16'h1711;
         16'hd8e0, 16'hd8e1, 16'hd8e2, 16'hd8e3, 16'hd8e4, 16'hd8e5, 16'hd8e6, 16'hd8e7 	:	val_out <= 16'h171f;
         16'hd8e8, 16'hd8e9, 16'hd8ea, 16'hd8eb, 16'hd8ec, 16'hd8ed, 16'hd8ee, 16'hd8ef 	:	val_out <= 16'h172e;
         16'hd8f0, 16'hd8f1, 16'hd8f2, 16'hd8f3, 16'hd8f4, 16'hd8f5, 16'hd8f6, 16'hd8f7 	:	val_out <= 16'h173c;
         16'hd8f8, 16'hd8f9, 16'hd8fa, 16'hd8fb, 16'hd8fc, 16'hd8fd, 16'hd8fe, 16'hd8ff 	:	val_out <= 16'h174a;
         16'hd900, 16'hd901, 16'hd902, 16'hd903, 16'hd904, 16'hd905, 16'hd906, 16'hd907 	:	val_out <= 16'h1759;
         16'hd908, 16'hd909, 16'hd90a, 16'hd90b, 16'hd90c, 16'hd90d, 16'hd90e, 16'hd90f 	:	val_out <= 16'h1767;
         16'hd910, 16'hd911, 16'hd912, 16'hd913, 16'hd914, 16'hd915, 16'hd916, 16'hd917 	:	val_out <= 16'h1776;
         16'hd918, 16'hd919, 16'hd91a, 16'hd91b, 16'hd91c, 16'hd91d, 16'hd91e, 16'hd91f 	:	val_out <= 16'h1784;
         16'hd920, 16'hd921, 16'hd922, 16'hd923, 16'hd924, 16'hd925, 16'hd926, 16'hd927 	:	val_out <= 16'h1793;
         16'hd928, 16'hd929, 16'hd92a, 16'hd92b, 16'hd92c, 16'hd92d, 16'hd92e, 16'hd92f 	:	val_out <= 16'h17a1;
         16'hd930, 16'hd931, 16'hd932, 16'hd933, 16'hd934, 16'hd935, 16'hd936, 16'hd937 	:	val_out <= 16'h17b0;
         16'hd938, 16'hd939, 16'hd93a, 16'hd93b, 16'hd93c, 16'hd93d, 16'hd93e, 16'hd93f 	:	val_out <= 16'h17bf;
         16'hd940, 16'hd941, 16'hd942, 16'hd943, 16'hd944, 16'hd945, 16'hd946, 16'hd947 	:	val_out <= 16'h17cd;
         16'hd948, 16'hd949, 16'hd94a, 16'hd94b, 16'hd94c, 16'hd94d, 16'hd94e, 16'hd94f 	:	val_out <= 16'h17dc;
         16'hd950, 16'hd951, 16'hd952, 16'hd953, 16'hd954, 16'hd955, 16'hd956, 16'hd957 	:	val_out <= 16'h17ea;
         16'hd958, 16'hd959, 16'hd95a, 16'hd95b, 16'hd95c, 16'hd95d, 16'hd95e, 16'hd95f 	:	val_out <= 16'h17f9;
         16'hd960, 16'hd961, 16'hd962, 16'hd963, 16'hd964, 16'hd965, 16'hd966, 16'hd967 	:	val_out <= 16'h1808;
         16'hd968, 16'hd969, 16'hd96a, 16'hd96b, 16'hd96c, 16'hd96d, 16'hd96e, 16'hd96f 	:	val_out <= 16'h1816;
         16'hd970, 16'hd971, 16'hd972, 16'hd973, 16'hd974, 16'hd975, 16'hd976, 16'hd977 	:	val_out <= 16'h1825;
         16'hd978, 16'hd979, 16'hd97a, 16'hd97b, 16'hd97c, 16'hd97d, 16'hd97e, 16'hd97f 	:	val_out <= 16'h1834;
         16'hd980, 16'hd981, 16'hd982, 16'hd983, 16'hd984, 16'hd985, 16'hd986, 16'hd987 	:	val_out <= 16'h1842;
         16'hd988, 16'hd989, 16'hd98a, 16'hd98b, 16'hd98c, 16'hd98d, 16'hd98e, 16'hd98f 	:	val_out <= 16'h1851;
         16'hd990, 16'hd991, 16'hd992, 16'hd993, 16'hd994, 16'hd995, 16'hd996, 16'hd997 	:	val_out <= 16'h1860;
         16'hd998, 16'hd999, 16'hd99a, 16'hd99b, 16'hd99c, 16'hd99d, 16'hd99e, 16'hd99f 	:	val_out <= 16'h186f;
         16'hd9a0, 16'hd9a1, 16'hd9a2, 16'hd9a3, 16'hd9a4, 16'hd9a5, 16'hd9a6, 16'hd9a7 	:	val_out <= 16'h187d;
         16'hd9a8, 16'hd9a9, 16'hd9aa, 16'hd9ab, 16'hd9ac, 16'hd9ad, 16'hd9ae, 16'hd9af 	:	val_out <= 16'h188c;
         16'hd9b0, 16'hd9b1, 16'hd9b2, 16'hd9b3, 16'hd9b4, 16'hd9b5, 16'hd9b6, 16'hd9b7 	:	val_out <= 16'h189b;
         16'hd9b8, 16'hd9b9, 16'hd9ba, 16'hd9bb, 16'hd9bc, 16'hd9bd, 16'hd9be, 16'hd9bf 	:	val_out <= 16'h18aa;
         16'hd9c0, 16'hd9c1, 16'hd9c2, 16'hd9c3, 16'hd9c4, 16'hd9c5, 16'hd9c6, 16'hd9c7 	:	val_out <= 16'h18b9;
         16'hd9c8, 16'hd9c9, 16'hd9ca, 16'hd9cb, 16'hd9cc, 16'hd9cd, 16'hd9ce, 16'hd9cf 	:	val_out <= 16'h18c8;
         16'hd9d0, 16'hd9d1, 16'hd9d2, 16'hd9d3, 16'hd9d4, 16'hd9d5, 16'hd9d6, 16'hd9d7 	:	val_out <= 16'h18d6;
         16'hd9d8, 16'hd9d9, 16'hd9da, 16'hd9db, 16'hd9dc, 16'hd9dd, 16'hd9de, 16'hd9df 	:	val_out <= 16'h18e5;
         16'hd9e0, 16'hd9e1, 16'hd9e2, 16'hd9e3, 16'hd9e4, 16'hd9e5, 16'hd9e6, 16'hd9e7 	:	val_out <= 16'h18f4;
         16'hd9e8, 16'hd9e9, 16'hd9ea, 16'hd9eb, 16'hd9ec, 16'hd9ed, 16'hd9ee, 16'hd9ef 	:	val_out <= 16'h1903;
         16'hd9f0, 16'hd9f1, 16'hd9f2, 16'hd9f3, 16'hd9f4, 16'hd9f5, 16'hd9f6, 16'hd9f7 	:	val_out <= 16'h1912;
         16'hd9f8, 16'hd9f9, 16'hd9fa, 16'hd9fb, 16'hd9fc, 16'hd9fd, 16'hd9fe, 16'hd9ff 	:	val_out <= 16'h1921;
         16'hda00, 16'hda01, 16'hda02, 16'hda03, 16'hda04, 16'hda05, 16'hda06, 16'hda07 	:	val_out <= 16'h1930;
         16'hda08, 16'hda09, 16'hda0a, 16'hda0b, 16'hda0c, 16'hda0d, 16'hda0e, 16'hda0f 	:	val_out <= 16'h193f;
         16'hda10, 16'hda11, 16'hda12, 16'hda13, 16'hda14, 16'hda15, 16'hda16, 16'hda17 	:	val_out <= 16'h194e;
         16'hda18, 16'hda19, 16'hda1a, 16'hda1b, 16'hda1c, 16'hda1d, 16'hda1e, 16'hda1f 	:	val_out <= 16'h195d;
         16'hda20, 16'hda21, 16'hda22, 16'hda23, 16'hda24, 16'hda25, 16'hda26, 16'hda27 	:	val_out <= 16'h196c;
         16'hda28, 16'hda29, 16'hda2a, 16'hda2b, 16'hda2c, 16'hda2d, 16'hda2e, 16'hda2f 	:	val_out <= 16'h197b;
         16'hda30, 16'hda31, 16'hda32, 16'hda33, 16'hda34, 16'hda35, 16'hda36, 16'hda37 	:	val_out <= 16'h198a;
         16'hda38, 16'hda39, 16'hda3a, 16'hda3b, 16'hda3c, 16'hda3d, 16'hda3e, 16'hda3f 	:	val_out <= 16'h1999;
         16'hda40, 16'hda41, 16'hda42, 16'hda43, 16'hda44, 16'hda45, 16'hda46, 16'hda47 	:	val_out <= 16'h19a8;
         16'hda48, 16'hda49, 16'hda4a, 16'hda4b, 16'hda4c, 16'hda4d, 16'hda4e, 16'hda4f 	:	val_out <= 16'h19b7;
         16'hda50, 16'hda51, 16'hda52, 16'hda53, 16'hda54, 16'hda55, 16'hda56, 16'hda57 	:	val_out <= 16'h19c6;
         16'hda58, 16'hda59, 16'hda5a, 16'hda5b, 16'hda5c, 16'hda5d, 16'hda5e, 16'hda5f 	:	val_out <= 16'h19d6;
         16'hda60, 16'hda61, 16'hda62, 16'hda63, 16'hda64, 16'hda65, 16'hda66, 16'hda67 	:	val_out <= 16'h19e5;
         16'hda68, 16'hda69, 16'hda6a, 16'hda6b, 16'hda6c, 16'hda6d, 16'hda6e, 16'hda6f 	:	val_out <= 16'h19f4;
         16'hda70, 16'hda71, 16'hda72, 16'hda73, 16'hda74, 16'hda75, 16'hda76, 16'hda77 	:	val_out <= 16'h1a03;
         16'hda78, 16'hda79, 16'hda7a, 16'hda7b, 16'hda7c, 16'hda7d, 16'hda7e, 16'hda7f 	:	val_out <= 16'h1a12;
         16'hda80, 16'hda81, 16'hda82, 16'hda83, 16'hda84, 16'hda85, 16'hda86, 16'hda87 	:	val_out <= 16'h1a22;
         16'hda88, 16'hda89, 16'hda8a, 16'hda8b, 16'hda8c, 16'hda8d, 16'hda8e, 16'hda8f 	:	val_out <= 16'h1a31;
         16'hda90, 16'hda91, 16'hda92, 16'hda93, 16'hda94, 16'hda95, 16'hda96, 16'hda97 	:	val_out <= 16'h1a40;
         16'hda98, 16'hda99, 16'hda9a, 16'hda9b, 16'hda9c, 16'hda9d, 16'hda9e, 16'hda9f 	:	val_out <= 16'h1a4f;
         16'hdaa0, 16'hdaa1, 16'hdaa2, 16'hdaa3, 16'hdaa4, 16'hdaa5, 16'hdaa6, 16'hdaa7 	:	val_out <= 16'h1a5f;
         16'hdaa8, 16'hdaa9, 16'hdaaa, 16'hdaab, 16'hdaac, 16'hdaad, 16'hdaae, 16'hdaaf 	:	val_out <= 16'h1a6e;
         16'hdab0, 16'hdab1, 16'hdab2, 16'hdab3, 16'hdab4, 16'hdab5, 16'hdab6, 16'hdab7 	:	val_out <= 16'h1a7d;
         16'hdab8, 16'hdab9, 16'hdaba, 16'hdabb, 16'hdabc, 16'hdabd, 16'hdabe, 16'hdabf 	:	val_out <= 16'h1a8c;
         16'hdac0, 16'hdac1, 16'hdac2, 16'hdac3, 16'hdac4, 16'hdac5, 16'hdac6, 16'hdac7 	:	val_out <= 16'h1a9c;
         16'hdac8, 16'hdac9, 16'hdaca, 16'hdacb, 16'hdacc, 16'hdacd, 16'hdace, 16'hdacf 	:	val_out <= 16'h1aab;
         16'hdad0, 16'hdad1, 16'hdad2, 16'hdad3, 16'hdad4, 16'hdad5, 16'hdad6, 16'hdad7 	:	val_out <= 16'h1aba;
         16'hdad8, 16'hdad9, 16'hdada, 16'hdadb, 16'hdadc, 16'hdadd, 16'hdade, 16'hdadf 	:	val_out <= 16'h1aca;
         16'hdae0, 16'hdae1, 16'hdae2, 16'hdae3, 16'hdae4, 16'hdae5, 16'hdae6, 16'hdae7 	:	val_out <= 16'h1ad9;
         16'hdae8, 16'hdae9, 16'hdaea, 16'hdaeb, 16'hdaec, 16'hdaed, 16'hdaee, 16'hdaef 	:	val_out <= 16'h1ae9;
         16'hdaf0, 16'hdaf1, 16'hdaf2, 16'hdaf3, 16'hdaf4, 16'hdaf5, 16'hdaf6, 16'hdaf7 	:	val_out <= 16'h1af8;
         16'hdaf8, 16'hdaf9, 16'hdafa, 16'hdafb, 16'hdafc, 16'hdafd, 16'hdafe, 16'hdaff 	:	val_out <= 16'h1b08;
         16'hdb00, 16'hdb01, 16'hdb02, 16'hdb03, 16'hdb04, 16'hdb05, 16'hdb06, 16'hdb07 	:	val_out <= 16'h1b17;
         16'hdb08, 16'hdb09, 16'hdb0a, 16'hdb0b, 16'hdb0c, 16'hdb0d, 16'hdb0e, 16'hdb0f 	:	val_out <= 16'h1b26;
         16'hdb10, 16'hdb11, 16'hdb12, 16'hdb13, 16'hdb14, 16'hdb15, 16'hdb16, 16'hdb17 	:	val_out <= 16'h1b36;
         16'hdb18, 16'hdb19, 16'hdb1a, 16'hdb1b, 16'hdb1c, 16'hdb1d, 16'hdb1e, 16'hdb1f 	:	val_out <= 16'h1b45;
         16'hdb20, 16'hdb21, 16'hdb22, 16'hdb23, 16'hdb24, 16'hdb25, 16'hdb26, 16'hdb27 	:	val_out <= 16'h1b55;
         16'hdb28, 16'hdb29, 16'hdb2a, 16'hdb2b, 16'hdb2c, 16'hdb2d, 16'hdb2e, 16'hdb2f 	:	val_out <= 16'h1b64;
         16'hdb30, 16'hdb31, 16'hdb32, 16'hdb33, 16'hdb34, 16'hdb35, 16'hdb36, 16'hdb37 	:	val_out <= 16'h1b74;
         16'hdb38, 16'hdb39, 16'hdb3a, 16'hdb3b, 16'hdb3c, 16'hdb3d, 16'hdb3e, 16'hdb3f 	:	val_out <= 16'h1b84;
         16'hdb40, 16'hdb41, 16'hdb42, 16'hdb43, 16'hdb44, 16'hdb45, 16'hdb46, 16'hdb47 	:	val_out <= 16'h1b93;
         16'hdb48, 16'hdb49, 16'hdb4a, 16'hdb4b, 16'hdb4c, 16'hdb4d, 16'hdb4e, 16'hdb4f 	:	val_out <= 16'h1ba3;
         16'hdb50, 16'hdb51, 16'hdb52, 16'hdb53, 16'hdb54, 16'hdb55, 16'hdb56, 16'hdb57 	:	val_out <= 16'h1bb2;
         16'hdb58, 16'hdb59, 16'hdb5a, 16'hdb5b, 16'hdb5c, 16'hdb5d, 16'hdb5e, 16'hdb5f 	:	val_out <= 16'h1bc2;
         16'hdb60, 16'hdb61, 16'hdb62, 16'hdb63, 16'hdb64, 16'hdb65, 16'hdb66, 16'hdb67 	:	val_out <= 16'h1bd2;
         16'hdb68, 16'hdb69, 16'hdb6a, 16'hdb6b, 16'hdb6c, 16'hdb6d, 16'hdb6e, 16'hdb6f 	:	val_out <= 16'h1be1;
         16'hdb70, 16'hdb71, 16'hdb72, 16'hdb73, 16'hdb74, 16'hdb75, 16'hdb76, 16'hdb77 	:	val_out <= 16'h1bf1;
         16'hdb78, 16'hdb79, 16'hdb7a, 16'hdb7b, 16'hdb7c, 16'hdb7d, 16'hdb7e, 16'hdb7f 	:	val_out <= 16'h1c01;
         16'hdb80, 16'hdb81, 16'hdb82, 16'hdb83, 16'hdb84, 16'hdb85, 16'hdb86, 16'hdb87 	:	val_out <= 16'h1c10;
         16'hdb88, 16'hdb89, 16'hdb8a, 16'hdb8b, 16'hdb8c, 16'hdb8d, 16'hdb8e, 16'hdb8f 	:	val_out <= 16'h1c20;
         16'hdb90, 16'hdb91, 16'hdb92, 16'hdb93, 16'hdb94, 16'hdb95, 16'hdb96, 16'hdb97 	:	val_out <= 16'h1c30;
         16'hdb98, 16'hdb99, 16'hdb9a, 16'hdb9b, 16'hdb9c, 16'hdb9d, 16'hdb9e, 16'hdb9f 	:	val_out <= 16'h1c3f;
         16'hdba0, 16'hdba1, 16'hdba2, 16'hdba3, 16'hdba4, 16'hdba5, 16'hdba6, 16'hdba7 	:	val_out <= 16'h1c4f;
         16'hdba8, 16'hdba9, 16'hdbaa, 16'hdbab, 16'hdbac, 16'hdbad, 16'hdbae, 16'hdbaf 	:	val_out <= 16'h1c5f;
         16'hdbb0, 16'hdbb1, 16'hdbb2, 16'hdbb3, 16'hdbb4, 16'hdbb5, 16'hdbb6, 16'hdbb7 	:	val_out <= 16'h1c6f;
         16'hdbb8, 16'hdbb9, 16'hdbba, 16'hdbbb, 16'hdbbc, 16'hdbbd, 16'hdbbe, 16'hdbbf 	:	val_out <= 16'h1c7f;
         16'hdbc0, 16'hdbc1, 16'hdbc2, 16'hdbc3, 16'hdbc4, 16'hdbc5, 16'hdbc6, 16'hdbc7 	:	val_out <= 16'h1c8e;
         16'hdbc8, 16'hdbc9, 16'hdbca, 16'hdbcb, 16'hdbcc, 16'hdbcd, 16'hdbce, 16'hdbcf 	:	val_out <= 16'h1c9e;
         16'hdbd0, 16'hdbd1, 16'hdbd2, 16'hdbd3, 16'hdbd4, 16'hdbd5, 16'hdbd6, 16'hdbd7 	:	val_out <= 16'h1cae;
         16'hdbd8, 16'hdbd9, 16'hdbda, 16'hdbdb, 16'hdbdc, 16'hdbdd, 16'hdbde, 16'hdbdf 	:	val_out <= 16'h1cbe;
         16'hdbe0, 16'hdbe1, 16'hdbe2, 16'hdbe3, 16'hdbe4, 16'hdbe5, 16'hdbe6, 16'hdbe7 	:	val_out <= 16'h1cce;
         16'hdbe8, 16'hdbe9, 16'hdbea, 16'hdbeb, 16'hdbec, 16'hdbed, 16'hdbee, 16'hdbef 	:	val_out <= 16'h1cde;
         16'hdbf0, 16'hdbf1, 16'hdbf2, 16'hdbf3, 16'hdbf4, 16'hdbf5, 16'hdbf6, 16'hdbf7 	:	val_out <= 16'h1cee;
         16'hdbf8, 16'hdbf9, 16'hdbfa, 16'hdbfb, 16'hdbfc, 16'hdbfd, 16'hdbfe, 16'hdbff 	:	val_out <= 16'h1cfe;
         16'hdc00, 16'hdc01, 16'hdc02, 16'hdc03, 16'hdc04, 16'hdc05, 16'hdc06, 16'hdc07 	:	val_out <= 16'h1d0d;
         16'hdc08, 16'hdc09, 16'hdc0a, 16'hdc0b, 16'hdc0c, 16'hdc0d, 16'hdc0e, 16'hdc0f 	:	val_out <= 16'h1d1d;
         16'hdc10, 16'hdc11, 16'hdc12, 16'hdc13, 16'hdc14, 16'hdc15, 16'hdc16, 16'hdc17 	:	val_out <= 16'h1d2d;
         16'hdc18, 16'hdc19, 16'hdc1a, 16'hdc1b, 16'hdc1c, 16'hdc1d, 16'hdc1e, 16'hdc1f 	:	val_out <= 16'h1d3d;
         16'hdc20, 16'hdc21, 16'hdc22, 16'hdc23, 16'hdc24, 16'hdc25, 16'hdc26, 16'hdc27 	:	val_out <= 16'h1d4d;
         16'hdc28, 16'hdc29, 16'hdc2a, 16'hdc2b, 16'hdc2c, 16'hdc2d, 16'hdc2e, 16'hdc2f 	:	val_out <= 16'h1d5d;
         16'hdc30, 16'hdc31, 16'hdc32, 16'hdc33, 16'hdc34, 16'hdc35, 16'hdc36, 16'hdc37 	:	val_out <= 16'h1d6d;
         16'hdc38, 16'hdc39, 16'hdc3a, 16'hdc3b, 16'hdc3c, 16'hdc3d, 16'hdc3e, 16'hdc3f 	:	val_out <= 16'h1d7d;
         16'hdc40, 16'hdc41, 16'hdc42, 16'hdc43, 16'hdc44, 16'hdc45, 16'hdc46, 16'hdc47 	:	val_out <= 16'h1d8e;
         16'hdc48, 16'hdc49, 16'hdc4a, 16'hdc4b, 16'hdc4c, 16'hdc4d, 16'hdc4e, 16'hdc4f 	:	val_out <= 16'h1d9e;
         16'hdc50, 16'hdc51, 16'hdc52, 16'hdc53, 16'hdc54, 16'hdc55, 16'hdc56, 16'hdc57 	:	val_out <= 16'h1dae;
         16'hdc58, 16'hdc59, 16'hdc5a, 16'hdc5b, 16'hdc5c, 16'hdc5d, 16'hdc5e, 16'hdc5f 	:	val_out <= 16'h1dbe;
         16'hdc60, 16'hdc61, 16'hdc62, 16'hdc63, 16'hdc64, 16'hdc65, 16'hdc66, 16'hdc67 	:	val_out <= 16'h1dce;
         16'hdc68, 16'hdc69, 16'hdc6a, 16'hdc6b, 16'hdc6c, 16'hdc6d, 16'hdc6e, 16'hdc6f 	:	val_out <= 16'h1dde;
         16'hdc70, 16'hdc71, 16'hdc72, 16'hdc73, 16'hdc74, 16'hdc75, 16'hdc76, 16'hdc77 	:	val_out <= 16'h1dee;
         16'hdc78, 16'hdc79, 16'hdc7a, 16'hdc7b, 16'hdc7c, 16'hdc7d, 16'hdc7e, 16'hdc7f 	:	val_out <= 16'h1dfe;
         16'hdc80, 16'hdc81, 16'hdc82, 16'hdc83, 16'hdc84, 16'hdc85, 16'hdc86, 16'hdc87 	:	val_out <= 16'h1e0e;
         16'hdc88, 16'hdc89, 16'hdc8a, 16'hdc8b, 16'hdc8c, 16'hdc8d, 16'hdc8e, 16'hdc8f 	:	val_out <= 16'h1e1f;
         16'hdc90, 16'hdc91, 16'hdc92, 16'hdc93, 16'hdc94, 16'hdc95, 16'hdc96, 16'hdc97 	:	val_out <= 16'h1e2f;
         16'hdc98, 16'hdc99, 16'hdc9a, 16'hdc9b, 16'hdc9c, 16'hdc9d, 16'hdc9e, 16'hdc9f 	:	val_out <= 16'h1e3f;
         16'hdca0, 16'hdca1, 16'hdca2, 16'hdca3, 16'hdca4, 16'hdca5, 16'hdca6, 16'hdca7 	:	val_out <= 16'h1e4f;
         16'hdca8, 16'hdca9, 16'hdcaa, 16'hdcab, 16'hdcac, 16'hdcad, 16'hdcae, 16'hdcaf 	:	val_out <= 16'h1e60;
         16'hdcb0, 16'hdcb1, 16'hdcb2, 16'hdcb3, 16'hdcb4, 16'hdcb5, 16'hdcb6, 16'hdcb7 	:	val_out <= 16'h1e70;
         16'hdcb8, 16'hdcb9, 16'hdcba, 16'hdcbb, 16'hdcbc, 16'hdcbd, 16'hdcbe, 16'hdcbf 	:	val_out <= 16'h1e80;
         16'hdcc0, 16'hdcc1, 16'hdcc2, 16'hdcc3, 16'hdcc4, 16'hdcc5, 16'hdcc6, 16'hdcc7 	:	val_out <= 16'h1e90;
         16'hdcc8, 16'hdcc9, 16'hdcca, 16'hdccb, 16'hdccc, 16'hdccd, 16'hdcce, 16'hdccf 	:	val_out <= 16'h1ea1;
         16'hdcd0, 16'hdcd1, 16'hdcd2, 16'hdcd3, 16'hdcd4, 16'hdcd5, 16'hdcd6, 16'hdcd7 	:	val_out <= 16'h1eb1;
         16'hdcd8, 16'hdcd9, 16'hdcda, 16'hdcdb, 16'hdcdc, 16'hdcdd, 16'hdcde, 16'hdcdf 	:	val_out <= 16'h1ec1;
         16'hdce0, 16'hdce1, 16'hdce2, 16'hdce3, 16'hdce4, 16'hdce5, 16'hdce6, 16'hdce7 	:	val_out <= 16'h1ed2;
         16'hdce8, 16'hdce9, 16'hdcea, 16'hdceb, 16'hdcec, 16'hdced, 16'hdcee, 16'hdcef 	:	val_out <= 16'h1ee2;
         16'hdcf0, 16'hdcf1, 16'hdcf2, 16'hdcf3, 16'hdcf4, 16'hdcf5, 16'hdcf6, 16'hdcf7 	:	val_out <= 16'h1ef2;
         16'hdcf8, 16'hdcf9, 16'hdcfa, 16'hdcfb, 16'hdcfc, 16'hdcfd, 16'hdcfe, 16'hdcff 	:	val_out <= 16'h1f03;
         16'hdd00, 16'hdd01, 16'hdd02, 16'hdd03, 16'hdd04, 16'hdd05, 16'hdd06, 16'hdd07 	:	val_out <= 16'h1f13;
         16'hdd08, 16'hdd09, 16'hdd0a, 16'hdd0b, 16'hdd0c, 16'hdd0d, 16'hdd0e, 16'hdd0f 	:	val_out <= 16'h1f24;
         16'hdd10, 16'hdd11, 16'hdd12, 16'hdd13, 16'hdd14, 16'hdd15, 16'hdd16, 16'hdd17 	:	val_out <= 16'h1f34;
         16'hdd18, 16'hdd19, 16'hdd1a, 16'hdd1b, 16'hdd1c, 16'hdd1d, 16'hdd1e, 16'hdd1f 	:	val_out <= 16'h1f45;
         16'hdd20, 16'hdd21, 16'hdd22, 16'hdd23, 16'hdd24, 16'hdd25, 16'hdd26, 16'hdd27 	:	val_out <= 16'h1f55;
         16'hdd28, 16'hdd29, 16'hdd2a, 16'hdd2b, 16'hdd2c, 16'hdd2d, 16'hdd2e, 16'hdd2f 	:	val_out <= 16'h1f66;
         16'hdd30, 16'hdd31, 16'hdd32, 16'hdd33, 16'hdd34, 16'hdd35, 16'hdd36, 16'hdd37 	:	val_out <= 16'h1f76;
         16'hdd38, 16'hdd39, 16'hdd3a, 16'hdd3b, 16'hdd3c, 16'hdd3d, 16'hdd3e, 16'hdd3f 	:	val_out <= 16'h1f87;
         16'hdd40, 16'hdd41, 16'hdd42, 16'hdd43, 16'hdd44, 16'hdd45, 16'hdd46, 16'hdd47 	:	val_out <= 16'h1f97;
         16'hdd48, 16'hdd49, 16'hdd4a, 16'hdd4b, 16'hdd4c, 16'hdd4d, 16'hdd4e, 16'hdd4f 	:	val_out <= 16'h1fa8;
         16'hdd50, 16'hdd51, 16'hdd52, 16'hdd53, 16'hdd54, 16'hdd55, 16'hdd56, 16'hdd57 	:	val_out <= 16'h1fb8;
         16'hdd58, 16'hdd59, 16'hdd5a, 16'hdd5b, 16'hdd5c, 16'hdd5d, 16'hdd5e, 16'hdd5f 	:	val_out <= 16'h1fc9;
         16'hdd60, 16'hdd61, 16'hdd62, 16'hdd63, 16'hdd64, 16'hdd65, 16'hdd66, 16'hdd67 	:	val_out <= 16'h1fd9;
         16'hdd68, 16'hdd69, 16'hdd6a, 16'hdd6b, 16'hdd6c, 16'hdd6d, 16'hdd6e, 16'hdd6f 	:	val_out <= 16'h1fea;
         16'hdd70, 16'hdd71, 16'hdd72, 16'hdd73, 16'hdd74, 16'hdd75, 16'hdd76, 16'hdd77 	:	val_out <= 16'h1ffb;
         16'hdd78, 16'hdd79, 16'hdd7a, 16'hdd7b, 16'hdd7c, 16'hdd7d, 16'hdd7e, 16'hdd7f 	:	val_out <= 16'h200b;
         16'hdd80, 16'hdd81, 16'hdd82, 16'hdd83, 16'hdd84, 16'hdd85, 16'hdd86, 16'hdd87 	:	val_out <= 16'h201c;
         16'hdd88, 16'hdd89, 16'hdd8a, 16'hdd8b, 16'hdd8c, 16'hdd8d, 16'hdd8e, 16'hdd8f 	:	val_out <= 16'h202c;
         16'hdd90, 16'hdd91, 16'hdd92, 16'hdd93, 16'hdd94, 16'hdd95, 16'hdd96, 16'hdd97 	:	val_out <= 16'h203d;
         16'hdd98, 16'hdd99, 16'hdd9a, 16'hdd9b, 16'hdd9c, 16'hdd9d, 16'hdd9e, 16'hdd9f 	:	val_out <= 16'h204e;
         16'hdda0, 16'hdda1, 16'hdda2, 16'hdda3, 16'hdda4, 16'hdda5, 16'hdda6, 16'hdda7 	:	val_out <= 16'h205f;
         16'hdda8, 16'hdda9, 16'hddaa, 16'hddab, 16'hddac, 16'hddad, 16'hddae, 16'hddaf 	:	val_out <= 16'h206f;
         16'hddb0, 16'hddb1, 16'hddb2, 16'hddb3, 16'hddb4, 16'hddb5, 16'hddb6, 16'hddb7 	:	val_out <= 16'h2080;
         16'hddb8, 16'hddb9, 16'hddba, 16'hddbb, 16'hddbc, 16'hddbd, 16'hddbe, 16'hddbf 	:	val_out <= 16'h2091;
         16'hddc0, 16'hddc1, 16'hddc2, 16'hddc3, 16'hddc4, 16'hddc5, 16'hddc6, 16'hddc7 	:	val_out <= 16'h20a1;
         16'hddc8, 16'hddc9, 16'hddca, 16'hddcb, 16'hddcc, 16'hddcd, 16'hddce, 16'hddcf 	:	val_out <= 16'h20b2;
         16'hddd0, 16'hddd1, 16'hddd2, 16'hddd3, 16'hddd4, 16'hddd5, 16'hddd6, 16'hddd7 	:	val_out <= 16'h20c3;
         16'hddd8, 16'hddd9, 16'hddda, 16'hdddb, 16'hdddc, 16'hdddd, 16'hddde, 16'hdddf 	:	val_out <= 16'h20d4;
         16'hdde0, 16'hdde1, 16'hdde2, 16'hdde3, 16'hdde4, 16'hdde5, 16'hdde6, 16'hdde7 	:	val_out <= 16'h20e5;
         16'hdde8, 16'hdde9, 16'hddea, 16'hddeb, 16'hddec, 16'hdded, 16'hddee, 16'hddef 	:	val_out <= 16'h20f5;
         16'hddf0, 16'hddf1, 16'hddf2, 16'hddf3, 16'hddf4, 16'hddf5, 16'hddf6, 16'hddf7 	:	val_out <= 16'h2106;
         16'hddf8, 16'hddf9, 16'hddfa, 16'hddfb, 16'hddfc, 16'hddfd, 16'hddfe, 16'hddff 	:	val_out <= 16'h2117;
         16'hde00, 16'hde01, 16'hde02, 16'hde03, 16'hde04, 16'hde05, 16'hde06, 16'hde07 	:	val_out <= 16'h2128;
         16'hde08, 16'hde09, 16'hde0a, 16'hde0b, 16'hde0c, 16'hde0d, 16'hde0e, 16'hde0f 	:	val_out <= 16'h2139;
         16'hde10, 16'hde11, 16'hde12, 16'hde13, 16'hde14, 16'hde15, 16'hde16, 16'hde17 	:	val_out <= 16'h214a;
         16'hde18, 16'hde19, 16'hde1a, 16'hde1b, 16'hde1c, 16'hde1d, 16'hde1e, 16'hde1f 	:	val_out <= 16'h215b;
         16'hde20, 16'hde21, 16'hde22, 16'hde23, 16'hde24, 16'hde25, 16'hde26, 16'hde27 	:	val_out <= 16'h216c;
         16'hde28, 16'hde29, 16'hde2a, 16'hde2b, 16'hde2c, 16'hde2d, 16'hde2e, 16'hde2f 	:	val_out <= 16'h217d;
         16'hde30, 16'hde31, 16'hde32, 16'hde33, 16'hde34, 16'hde35, 16'hde36, 16'hde37 	:	val_out <= 16'h218e;
         16'hde38, 16'hde39, 16'hde3a, 16'hde3b, 16'hde3c, 16'hde3d, 16'hde3e, 16'hde3f 	:	val_out <= 16'h219f;
         16'hde40, 16'hde41, 16'hde42, 16'hde43, 16'hde44, 16'hde45, 16'hde46, 16'hde47 	:	val_out <= 16'h21af;
         16'hde48, 16'hde49, 16'hde4a, 16'hde4b, 16'hde4c, 16'hde4d, 16'hde4e, 16'hde4f 	:	val_out <= 16'h21c0;
         16'hde50, 16'hde51, 16'hde52, 16'hde53, 16'hde54, 16'hde55, 16'hde56, 16'hde57 	:	val_out <= 16'h21d2;
         16'hde58, 16'hde59, 16'hde5a, 16'hde5b, 16'hde5c, 16'hde5d, 16'hde5e, 16'hde5f 	:	val_out <= 16'h21e3;
         16'hde60, 16'hde61, 16'hde62, 16'hde63, 16'hde64, 16'hde65, 16'hde66, 16'hde67 	:	val_out <= 16'h21f4;
         16'hde68, 16'hde69, 16'hde6a, 16'hde6b, 16'hde6c, 16'hde6d, 16'hde6e, 16'hde6f 	:	val_out <= 16'h2205;
         16'hde70, 16'hde71, 16'hde72, 16'hde73, 16'hde74, 16'hde75, 16'hde76, 16'hde77 	:	val_out <= 16'h2216;
         16'hde78, 16'hde79, 16'hde7a, 16'hde7b, 16'hde7c, 16'hde7d, 16'hde7e, 16'hde7f 	:	val_out <= 16'h2227;
         16'hde80, 16'hde81, 16'hde82, 16'hde83, 16'hde84, 16'hde85, 16'hde86, 16'hde87 	:	val_out <= 16'h2238;
         16'hde88, 16'hde89, 16'hde8a, 16'hde8b, 16'hde8c, 16'hde8d, 16'hde8e, 16'hde8f 	:	val_out <= 16'h2249;
         16'hde90, 16'hde91, 16'hde92, 16'hde93, 16'hde94, 16'hde95, 16'hde96, 16'hde97 	:	val_out <= 16'h225a;
         16'hde98, 16'hde99, 16'hde9a, 16'hde9b, 16'hde9c, 16'hde9d, 16'hde9e, 16'hde9f 	:	val_out <= 16'h226b;
         16'hdea0, 16'hdea1, 16'hdea2, 16'hdea3, 16'hdea4, 16'hdea5, 16'hdea6, 16'hdea7 	:	val_out <= 16'h227c;
         16'hdea8, 16'hdea9, 16'hdeaa, 16'hdeab, 16'hdeac, 16'hdead, 16'hdeae, 16'hdeaf 	:	val_out <= 16'h228e;
         16'hdeb0, 16'hdeb1, 16'hdeb2, 16'hdeb3, 16'hdeb4, 16'hdeb5, 16'hdeb6, 16'hdeb7 	:	val_out <= 16'h229f;
         16'hdeb8, 16'hdeb9, 16'hdeba, 16'hdebb, 16'hdebc, 16'hdebd, 16'hdebe, 16'hdebf 	:	val_out <= 16'h22b0;
         16'hdec0, 16'hdec1, 16'hdec2, 16'hdec3, 16'hdec4, 16'hdec5, 16'hdec6, 16'hdec7 	:	val_out <= 16'h22c1;
         16'hdec8, 16'hdec9, 16'hdeca, 16'hdecb, 16'hdecc, 16'hdecd, 16'hdece, 16'hdecf 	:	val_out <= 16'h22d2;
         16'hded0, 16'hded1, 16'hded2, 16'hded3, 16'hded4, 16'hded5, 16'hded6, 16'hded7 	:	val_out <= 16'h22e4;
         16'hded8, 16'hded9, 16'hdeda, 16'hdedb, 16'hdedc, 16'hdedd, 16'hdede, 16'hdedf 	:	val_out <= 16'h22f5;
         16'hdee0, 16'hdee1, 16'hdee2, 16'hdee3, 16'hdee4, 16'hdee5, 16'hdee6, 16'hdee7 	:	val_out <= 16'h2306;
         16'hdee8, 16'hdee9, 16'hdeea, 16'hdeeb, 16'hdeec, 16'hdeed, 16'hdeee, 16'hdeef 	:	val_out <= 16'h2317;
         16'hdef0, 16'hdef1, 16'hdef2, 16'hdef3, 16'hdef4, 16'hdef5, 16'hdef6, 16'hdef7 	:	val_out <= 16'h2329;
         16'hdef8, 16'hdef9, 16'hdefa, 16'hdefb, 16'hdefc, 16'hdefd, 16'hdefe, 16'hdeff 	:	val_out <= 16'h233a;
         16'hdf00, 16'hdf01, 16'hdf02, 16'hdf03, 16'hdf04, 16'hdf05, 16'hdf06, 16'hdf07 	:	val_out <= 16'h234b;
         16'hdf08, 16'hdf09, 16'hdf0a, 16'hdf0b, 16'hdf0c, 16'hdf0d, 16'hdf0e, 16'hdf0f 	:	val_out <= 16'h235d;
         16'hdf10, 16'hdf11, 16'hdf12, 16'hdf13, 16'hdf14, 16'hdf15, 16'hdf16, 16'hdf17 	:	val_out <= 16'h236e;
         16'hdf18, 16'hdf19, 16'hdf1a, 16'hdf1b, 16'hdf1c, 16'hdf1d, 16'hdf1e, 16'hdf1f 	:	val_out <= 16'h237f;
         16'hdf20, 16'hdf21, 16'hdf22, 16'hdf23, 16'hdf24, 16'hdf25, 16'hdf26, 16'hdf27 	:	val_out <= 16'h2391;
         16'hdf28, 16'hdf29, 16'hdf2a, 16'hdf2b, 16'hdf2c, 16'hdf2d, 16'hdf2e, 16'hdf2f 	:	val_out <= 16'h23a2;
         16'hdf30, 16'hdf31, 16'hdf32, 16'hdf33, 16'hdf34, 16'hdf35, 16'hdf36, 16'hdf37 	:	val_out <= 16'h23b4;
         16'hdf38, 16'hdf39, 16'hdf3a, 16'hdf3b, 16'hdf3c, 16'hdf3d, 16'hdf3e, 16'hdf3f 	:	val_out <= 16'h23c5;
         16'hdf40, 16'hdf41, 16'hdf42, 16'hdf43, 16'hdf44, 16'hdf45, 16'hdf46, 16'hdf47 	:	val_out <= 16'h23d6;
         16'hdf48, 16'hdf49, 16'hdf4a, 16'hdf4b, 16'hdf4c, 16'hdf4d, 16'hdf4e, 16'hdf4f 	:	val_out <= 16'h23e8;
         16'hdf50, 16'hdf51, 16'hdf52, 16'hdf53, 16'hdf54, 16'hdf55, 16'hdf56, 16'hdf57 	:	val_out <= 16'h23f9;
         16'hdf58, 16'hdf59, 16'hdf5a, 16'hdf5b, 16'hdf5c, 16'hdf5d, 16'hdf5e, 16'hdf5f 	:	val_out <= 16'h240b;
         16'hdf60, 16'hdf61, 16'hdf62, 16'hdf63, 16'hdf64, 16'hdf65, 16'hdf66, 16'hdf67 	:	val_out <= 16'h241c;
         16'hdf68, 16'hdf69, 16'hdf6a, 16'hdf6b, 16'hdf6c, 16'hdf6d, 16'hdf6e, 16'hdf6f 	:	val_out <= 16'h242e;
         16'hdf70, 16'hdf71, 16'hdf72, 16'hdf73, 16'hdf74, 16'hdf75, 16'hdf76, 16'hdf77 	:	val_out <= 16'h243f;
         16'hdf78, 16'hdf79, 16'hdf7a, 16'hdf7b, 16'hdf7c, 16'hdf7d, 16'hdf7e, 16'hdf7f 	:	val_out <= 16'h2451;
         16'hdf80, 16'hdf81, 16'hdf82, 16'hdf83, 16'hdf84, 16'hdf85, 16'hdf86, 16'hdf87 	:	val_out <= 16'h2462;
         16'hdf88, 16'hdf89, 16'hdf8a, 16'hdf8b, 16'hdf8c, 16'hdf8d, 16'hdf8e, 16'hdf8f 	:	val_out <= 16'h2474;
         16'hdf90, 16'hdf91, 16'hdf92, 16'hdf93, 16'hdf94, 16'hdf95, 16'hdf96, 16'hdf97 	:	val_out <= 16'h2486;
         16'hdf98, 16'hdf99, 16'hdf9a, 16'hdf9b, 16'hdf9c, 16'hdf9d, 16'hdf9e, 16'hdf9f 	:	val_out <= 16'h2497;
         16'hdfa0, 16'hdfa1, 16'hdfa2, 16'hdfa3, 16'hdfa4, 16'hdfa5, 16'hdfa6, 16'hdfa7 	:	val_out <= 16'h24a9;
         16'hdfa8, 16'hdfa9, 16'hdfaa, 16'hdfab, 16'hdfac, 16'hdfad, 16'hdfae, 16'hdfaf 	:	val_out <= 16'h24ba;
         16'hdfb0, 16'hdfb1, 16'hdfb2, 16'hdfb3, 16'hdfb4, 16'hdfb5, 16'hdfb6, 16'hdfb7 	:	val_out <= 16'h24cc;
         16'hdfb8, 16'hdfb9, 16'hdfba, 16'hdfbb, 16'hdfbc, 16'hdfbd, 16'hdfbe, 16'hdfbf 	:	val_out <= 16'h24de;
         16'hdfc0, 16'hdfc1, 16'hdfc2, 16'hdfc3, 16'hdfc4, 16'hdfc5, 16'hdfc6, 16'hdfc7 	:	val_out <= 16'h24ef;
         16'hdfc8, 16'hdfc9, 16'hdfca, 16'hdfcb, 16'hdfcc, 16'hdfcd, 16'hdfce, 16'hdfcf 	:	val_out <= 16'h2501;
         16'hdfd0, 16'hdfd1, 16'hdfd2, 16'hdfd3, 16'hdfd4, 16'hdfd5, 16'hdfd6, 16'hdfd7 	:	val_out <= 16'h2513;
         16'hdfd8, 16'hdfd9, 16'hdfda, 16'hdfdb, 16'hdfdc, 16'hdfdd, 16'hdfde, 16'hdfdf 	:	val_out <= 16'h2524;
         16'hdfe0, 16'hdfe1, 16'hdfe2, 16'hdfe3, 16'hdfe4, 16'hdfe5, 16'hdfe6, 16'hdfe7 	:	val_out <= 16'h2536;
         16'hdfe8, 16'hdfe9, 16'hdfea, 16'hdfeb, 16'hdfec, 16'hdfed, 16'hdfee, 16'hdfef 	:	val_out <= 16'h2548;
         16'hdff0, 16'hdff1, 16'hdff2, 16'hdff3, 16'hdff4, 16'hdff5, 16'hdff6, 16'hdff7 	:	val_out <= 16'h255a;
         16'hdff8, 16'hdff9, 16'hdffa, 16'hdffb, 16'hdffc, 16'hdffd, 16'hdffe, 16'hdfff 	:	val_out <= 16'h256b;
         16'he000, 16'he001, 16'he002, 16'he003, 16'he004, 16'he005, 16'he006, 16'he007 	:	val_out <= 16'h257d;
         16'he008, 16'he009, 16'he00a, 16'he00b, 16'he00c, 16'he00d, 16'he00e, 16'he00f 	:	val_out <= 16'h258f;
         16'he010, 16'he011, 16'he012, 16'he013, 16'he014, 16'he015, 16'he016, 16'he017 	:	val_out <= 16'h25a1;
         16'he018, 16'he019, 16'he01a, 16'he01b, 16'he01c, 16'he01d, 16'he01e, 16'he01f 	:	val_out <= 16'h25b2;
         16'he020, 16'he021, 16'he022, 16'he023, 16'he024, 16'he025, 16'he026, 16'he027 	:	val_out <= 16'h25c4;
         16'he028, 16'he029, 16'he02a, 16'he02b, 16'he02c, 16'he02d, 16'he02e, 16'he02f 	:	val_out <= 16'h25d6;
         16'he030, 16'he031, 16'he032, 16'he033, 16'he034, 16'he035, 16'he036, 16'he037 	:	val_out <= 16'h25e8;
         16'he038, 16'he039, 16'he03a, 16'he03b, 16'he03c, 16'he03d, 16'he03e, 16'he03f 	:	val_out <= 16'h25fa;
         16'he040, 16'he041, 16'he042, 16'he043, 16'he044, 16'he045, 16'he046, 16'he047 	:	val_out <= 16'h260c;
         16'he048, 16'he049, 16'he04a, 16'he04b, 16'he04c, 16'he04d, 16'he04e, 16'he04f 	:	val_out <= 16'h261e;
         16'he050, 16'he051, 16'he052, 16'he053, 16'he054, 16'he055, 16'he056, 16'he057 	:	val_out <= 16'h262f;
         16'he058, 16'he059, 16'he05a, 16'he05b, 16'he05c, 16'he05d, 16'he05e, 16'he05f 	:	val_out <= 16'h2641;
         16'he060, 16'he061, 16'he062, 16'he063, 16'he064, 16'he065, 16'he066, 16'he067 	:	val_out <= 16'h2653;
         16'he068, 16'he069, 16'he06a, 16'he06b, 16'he06c, 16'he06d, 16'he06e, 16'he06f 	:	val_out <= 16'h2665;
         16'he070, 16'he071, 16'he072, 16'he073, 16'he074, 16'he075, 16'he076, 16'he077 	:	val_out <= 16'h2677;
         16'he078, 16'he079, 16'he07a, 16'he07b, 16'he07c, 16'he07d, 16'he07e, 16'he07f 	:	val_out <= 16'h2689;
         16'he080, 16'he081, 16'he082, 16'he083, 16'he084, 16'he085, 16'he086, 16'he087 	:	val_out <= 16'h269b;
         16'he088, 16'he089, 16'he08a, 16'he08b, 16'he08c, 16'he08d, 16'he08e, 16'he08f 	:	val_out <= 16'h26ad;
         16'he090, 16'he091, 16'he092, 16'he093, 16'he094, 16'he095, 16'he096, 16'he097 	:	val_out <= 16'h26bf;
         16'he098, 16'he099, 16'he09a, 16'he09b, 16'he09c, 16'he09d, 16'he09e, 16'he09f 	:	val_out <= 16'h26d1;
         16'he0a0, 16'he0a1, 16'he0a2, 16'he0a3, 16'he0a4, 16'he0a5, 16'he0a6, 16'he0a7 	:	val_out <= 16'h26e3;
         16'he0a8, 16'he0a9, 16'he0aa, 16'he0ab, 16'he0ac, 16'he0ad, 16'he0ae, 16'he0af 	:	val_out <= 16'h26f5;
         16'he0b0, 16'he0b1, 16'he0b2, 16'he0b3, 16'he0b4, 16'he0b5, 16'he0b6, 16'he0b7 	:	val_out <= 16'h2707;
         16'he0b8, 16'he0b9, 16'he0ba, 16'he0bb, 16'he0bc, 16'he0bd, 16'he0be, 16'he0bf 	:	val_out <= 16'h2719;
         16'he0c0, 16'he0c1, 16'he0c2, 16'he0c3, 16'he0c4, 16'he0c5, 16'he0c6, 16'he0c7 	:	val_out <= 16'h272b;
         16'he0c8, 16'he0c9, 16'he0ca, 16'he0cb, 16'he0cc, 16'he0cd, 16'he0ce, 16'he0cf 	:	val_out <= 16'h273e;
         16'he0d0, 16'he0d1, 16'he0d2, 16'he0d3, 16'he0d4, 16'he0d5, 16'he0d6, 16'he0d7 	:	val_out <= 16'h2750;
         16'he0d8, 16'he0d9, 16'he0da, 16'he0db, 16'he0dc, 16'he0dd, 16'he0de, 16'he0df 	:	val_out <= 16'h2762;
         16'he0e0, 16'he0e1, 16'he0e2, 16'he0e3, 16'he0e4, 16'he0e5, 16'he0e6, 16'he0e7 	:	val_out <= 16'h2774;
         16'he0e8, 16'he0e9, 16'he0ea, 16'he0eb, 16'he0ec, 16'he0ed, 16'he0ee, 16'he0ef 	:	val_out <= 16'h2786;
         16'he0f0, 16'he0f1, 16'he0f2, 16'he0f3, 16'he0f4, 16'he0f5, 16'he0f6, 16'he0f7 	:	val_out <= 16'h2798;
         16'he0f8, 16'he0f9, 16'he0fa, 16'he0fb, 16'he0fc, 16'he0fd, 16'he0fe, 16'he0ff 	:	val_out <= 16'h27aa;
         16'he100, 16'he101, 16'he102, 16'he103, 16'he104, 16'he105, 16'he106, 16'he107 	:	val_out <= 16'h27bd;
         16'he108, 16'he109, 16'he10a, 16'he10b, 16'he10c, 16'he10d, 16'he10e, 16'he10f 	:	val_out <= 16'h27cf;
         16'he110, 16'he111, 16'he112, 16'he113, 16'he114, 16'he115, 16'he116, 16'he117 	:	val_out <= 16'h27e1;
         16'he118, 16'he119, 16'he11a, 16'he11b, 16'he11c, 16'he11d, 16'he11e, 16'he11f 	:	val_out <= 16'h27f3;
         16'he120, 16'he121, 16'he122, 16'he123, 16'he124, 16'he125, 16'he126, 16'he127 	:	val_out <= 16'h2806;
         16'he128, 16'he129, 16'he12a, 16'he12b, 16'he12c, 16'he12d, 16'he12e, 16'he12f 	:	val_out <= 16'h2818;
         16'he130, 16'he131, 16'he132, 16'he133, 16'he134, 16'he135, 16'he136, 16'he137 	:	val_out <= 16'h282a;
         16'he138, 16'he139, 16'he13a, 16'he13b, 16'he13c, 16'he13d, 16'he13e, 16'he13f 	:	val_out <= 16'h283c;
         16'he140, 16'he141, 16'he142, 16'he143, 16'he144, 16'he145, 16'he146, 16'he147 	:	val_out <= 16'h284f;
         16'he148, 16'he149, 16'he14a, 16'he14b, 16'he14c, 16'he14d, 16'he14e, 16'he14f 	:	val_out <= 16'h2861;
         16'he150, 16'he151, 16'he152, 16'he153, 16'he154, 16'he155, 16'he156, 16'he157 	:	val_out <= 16'h2873;
         16'he158, 16'he159, 16'he15a, 16'he15b, 16'he15c, 16'he15d, 16'he15e, 16'he15f 	:	val_out <= 16'h2886;
         16'he160, 16'he161, 16'he162, 16'he163, 16'he164, 16'he165, 16'he166, 16'he167 	:	val_out <= 16'h2898;
         16'he168, 16'he169, 16'he16a, 16'he16b, 16'he16c, 16'he16d, 16'he16e, 16'he16f 	:	val_out <= 16'h28aa;
         16'he170, 16'he171, 16'he172, 16'he173, 16'he174, 16'he175, 16'he176, 16'he177 	:	val_out <= 16'h28bd;
         16'he178, 16'he179, 16'he17a, 16'he17b, 16'he17c, 16'he17d, 16'he17e, 16'he17f 	:	val_out <= 16'h28cf;
         16'he180, 16'he181, 16'he182, 16'he183, 16'he184, 16'he185, 16'he186, 16'he187 	:	val_out <= 16'h28e2;
         16'he188, 16'he189, 16'he18a, 16'he18b, 16'he18c, 16'he18d, 16'he18e, 16'he18f 	:	val_out <= 16'h28f4;
         16'he190, 16'he191, 16'he192, 16'he193, 16'he194, 16'he195, 16'he196, 16'he197 	:	val_out <= 16'h2906;
         16'he198, 16'he199, 16'he19a, 16'he19b, 16'he19c, 16'he19d, 16'he19e, 16'he19f 	:	val_out <= 16'h2919;
         16'he1a0, 16'he1a1, 16'he1a2, 16'he1a3, 16'he1a4, 16'he1a5, 16'he1a6, 16'he1a7 	:	val_out <= 16'h292b;
         16'he1a8, 16'he1a9, 16'he1aa, 16'he1ab, 16'he1ac, 16'he1ad, 16'he1ae, 16'he1af 	:	val_out <= 16'h293e;
         16'he1b0, 16'he1b1, 16'he1b2, 16'he1b3, 16'he1b4, 16'he1b5, 16'he1b6, 16'he1b7 	:	val_out <= 16'h2950;
         16'he1b8, 16'he1b9, 16'he1ba, 16'he1bb, 16'he1bc, 16'he1bd, 16'he1be, 16'he1bf 	:	val_out <= 16'h2963;
         16'he1c0, 16'he1c1, 16'he1c2, 16'he1c3, 16'he1c4, 16'he1c5, 16'he1c6, 16'he1c7 	:	val_out <= 16'h2975;
         16'he1c8, 16'he1c9, 16'he1ca, 16'he1cb, 16'he1cc, 16'he1cd, 16'he1ce, 16'he1cf 	:	val_out <= 16'h2988;
         16'he1d0, 16'he1d1, 16'he1d2, 16'he1d3, 16'he1d4, 16'he1d5, 16'he1d6, 16'he1d7 	:	val_out <= 16'h299a;
         16'he1d8, 16'he1d9, 16'he1da, 16'he1db, 16'he1dc, 16'he1dd, 16'he1de, 16'he1df 	:	val_out <= 16'h29ad;
         16'he1e0, 16'he1e1, 16'he1e2, 16'he1e3, 16'he1e4, 16'he1e5, 16'he1e6, 16'he1e7 	:	val_out <= 16'h29bf;
         16'he1e8, 16'he1e9, 16'he1ea, 16'he1eb, 16'he1ec, 16'he1ed, 16'he1ee, 16'he1ef 	:	val_out <= 16'h29d2;
         16'he1f0, 16'he1f1, 16'he1f2, 16'he1f3, 16'he1f4, 16'he1f5, 16'he1f6, 16'he1f7 	:	val_out <= 16'h29e5;
         16'he1f8, 16'he1f9, 16'he1fa, 16'he1fb, 16'he1fc, 16'he1fd, 16'he1fe, 16'he1ff 	:	val_out <= 16'h29f7;
         16'he200, 16'he201, 16'he202, 16'he203, 16'he204, 16'he205, 16'he206, 16'he207 	:	val_out <= 16'h2a0a;
         16'he208, 16'he209, 16'he20a, 16'he20b, 16'he20c, 16'he20d, 16'he20e, 16'he20f 	:	val_out <= 16'h2a1c;
         16'he210, 16'he211, 16'he212, 16'he213, 16'he214, 16'he215, 16'he216, 16'he217 	:	val_out <= 16'h2a2f;
         16'he218, 16'he219, 16'he21a, 16'he21b, 16'he21c, 16'he21d, 16'he21e, 16'he21f 	:	val_out <= 16'h2a42;
         16'he220, 16'he221, 16'he222, 16'he223, 16'he224, 16'he225, 16'he226, 16'he227 	:	val_out <= 16'h2a54;
         16'he228, 16'he229, 16'he22a, 16'he22b, 16'he22c, 16'he22d, 16'he22e, 16'he22f 	:	val_out <= 16'h2a67;
         16'he230, 16'he231, 16'he232, 16'he233, 16'he234, 16'he235, 16'he236, 16'he237 	:	val_out <= 16'h2a7a;
         16'he238, 16'he239, 16'he23a, 16'he23b, 16'he23c, 16'he23d, 16'he23e, 16'he23f 	:	val_out <= 16'h2a8d;
         16'he240, 16'he241, 16'he242, 16'he243, 16'he244, 16'he245, 16'he246, 16'he247 	:	val_out <= 16'h2a9f;
         16'he248, 16'he249, 16'he24a, 16'he24b, 16'he24c, 16'he24d, 16'he24e, 16'he24f 	:	val_out <= 16'h2ab2;
         16'he250, 16'he251, 16'he252, 16'he253, 16'he254, 16'he255, 16'he256, 16'he257 	:	val_out <= 16'h2ac5;
         16'he258, 16'he259, 16'he25a, 16'he25b, 16'he25c, 16'he25d, 16'he25e, 16'he25f 	:	val_out <= 16'h2ad7;
         16'he260, 16'he261, 16'he262, 16'he263, 16'he264, 16'he265, 16'he266, 16'he267 	:	val_out <= 16'h2aea;
         16'he268, 16'he269, 16'he26a, 16'he26b, 16'he26c, 16'he26d, 16'he26e, 16'he26f 	:	val_out <= 16'h2afd;
         16'he270, 16'he271, 16'he272, 16'he273, 16'he274, 16'he275, 16'he276, 16'he277 	:	val_out <= 16'h2b10;
         16'he278, 16'he279, 16'he27a, 16'he27b, 16'he27c, 16'he27d, 16'he27e, 16'he27f 	:	val_out <= 16'h2b23;
         16'he280, 16'he281, 16'he282, 16'he283, 16'he284, 16'he285, 16'he286, 16'he287 	:	val_out <= 16'h2b35;
         16'he288, 16'he289, 16'he28a, 16'he28b, 16'he28c, 16'he28d, 16'he28e, 16'he28f 	:	val_out <= 16'h2b48;
         16'he290, 16'he291, 16'he292, 16'he293, 16'he294, 16'he295, 16'he296, 16'he297 	:	val_out <= 16'h2b5b;
         16'he298, 16'he299, 16'he29a, 16'he29b, 16'he29c, 16'he29d, 16'he29e, 16'he29f 	:	val_out <= 16'h2b6e;
         16'he2a0, 16'he2a1, 16'he2a2, 16'he2a3, 16'he2a4, 16'he2a5, 16'he2a6, 16'he2a7 	:	val_out <= 16'h2b81;
         16'he2a8, 16'he2a9, 16'he2aa, 16'he2ab, 16'he2ac, 16'he2ad, 16'he2ae, 16'he2af 	:	val_out <= 16'h2b94;
         16'he2b0, 16'he2b1, 16'he2b2, 16'he2b3, 16'he2b4, 16'he2b5, 16'he2b6, 16'he2b7 	:	val_out <= 16'h2ba7;
         16'he2b8, 16'he2b9, 16'he2ba, 16'he2bb, 16'he2bc, 16'he2bd, 16'he2be, 16'he2bf 	:	val_out <= 16'h2bba;
         16'he2c0, 16'he2c1, 16'he2c2, 16'he2c3, 16'he2c4, 16'he2c5, 16'he2c6, 16'he2c7 	:	val_out <= 16'h2bcc;
         16'he2c8, 16'he2c9, 16'he2ca, 16'he2cb, 16'he2cc, 16'he2cd, 16'he2ce, 16'he2cf 	:	val_out <= 16'h2bdf;
         16'he2d0, 16'he2d1, 16'he2d2, 16'he2d3, 16'he2d4, 16'he2d5, 16'he2d6, 16'he2d7 	:	val_out <= 16'h2bf2;
         16'he2d8, 16'he2d9, 16'he2da, 16'he2db, 16'he2dc, 16'he2dd, 16'he2de, 16'he2df 	:	val_out <= 16'h2c05;
         16'he2e0, 16'he2e1, 16'he2e2, 16'he2e3, 16'he2e4, 16'he2e5, 16'he2e6, 16'he2e7 	:	val_out <= 16'h2c18;
         16'he2e8, 16'he2e9, 16'he2ea, 16'he2eb, 16'he2ec, 16'he2ed, 16'he2ee, 16'he2ef 	:	val_out <= 16'h2c2b;
         16'he2f0, 16'he2f1, 16'he2f2, 16'he2f3, 16'he2f4, 16'he2f5, 16'he2f6, 16'he2f7 	:	val_out <= 16'h2c3e;
         16'he2f8, 16'he2f9, 16'he2fa, 16'he2fb, 16'he2fc, 16'he2fd, 16'he2fe, 16'he2ff 	:	val_out <= 16'h2c51;
         16'he300, 16'he301, 16'he302, 16'he303, 16'he304, 16'he305, 16'he306, 16'he307 	:	val_out <= 16'h2c64;
         16'he308, 16'he309, 16'he30a, 16'he30b, 16'he30c, 16'he30d, 16'he30e, 16'he30f 	:	val_out <= 16'h2c77;
         16'he310, 16'he311, 16'he312, 16'he313, 16'he314, 16'he315, 16'he316, 16'he317 	:	val_out <= 16'h2c8a;
         16'he318, 16'he319, 16'he31a, 16'he31b, 16'he31c, 16'he31d, 16'he31e, 16'he31f 	:	val_out <= 16'h2c9d;
         16'he320, 16'he321, 16'he322, 16'he323, 16'he324, 16'he325, 16'he326, 16'he327 	:	val_out <= 16'h2cb1;
         16'he328, 16'he329, 16'he32a, 16'he32b, 16'he32c, 16'he32d, 16'he32e, 16'he32f 	:	val_out <= 16'h2cc4;
         16'he330, 16'he331, 16'he332, 16'he333, 16'he334, 16'he335, 16'he336, 16'he337 	:	val_out <= 16'h2cd7;
         16'he338, 16'he339, 16'he33a, 16'he33b, 16'he33c, 16'he33d, 16'he33e, 16'he33f 	:	val_out <= 16'h2cea;
         16'he340, 16'he341, 16'he342, 16'he343, 16'he344, 16'he345, 16'he346, 16'he347 	:	val_out <= 16'h2cfd;
         16'he348, 16'he349, 16'he34a, 16'he34b, 16'he34c, 16'he34d, 16'he34e, 16'he34f 	:	val_out <= 16'h2d10;
         16'he350, 16'he351, 16'he352, 16'he353, 16'he354, 16'he355, 16'he356, 16'he357 	:	val_out <= 16'h2d23;
         16'he358, 16'he359, 16'he35a, 16'he35b, 16'he35c, 16'he35d, 16'he35e, 16'he35f 	:	val_out <= 16'h2d36;
         16'he360, 16'he361, 16'he362, 16'he363, 16'he364, 16'he365, 16'he366, 16'he367 	:	val_out <= 16'h2d4a;
         16'he368, 16'he369, 16'he36a, 16'he36b, 16'he36c, 16'he36d, 16'he36e, 16'he36f 	:	val_out <= 16'h2d5d;
         16'he370, 16'he371, 16'he372, 16'he373, 16'he374, 16'he375, 16'he376, 16'he377 	:	val_out <= 16'h2d70;
         16'he378, 16'he379, 16'he37a, 16'he37b, 16'he37c, 16'he37d, 16'he37e, 16'he37f 	:	val_out <= 16'h2d83;
         16'he380, 16'he381, 16'he382, 16'he383, 16'he384, 16'he385, 16'he386, 16'he387 	:	val_out <= 16'h2d96;
         16'he388, 16'he389, 16'he38a, 16'he38b, 16'he38c, 16'he38d, 16'he38e, 16'he38f 	:	val_out <= 16'h2daa;
         16'he390, 16'he391, 16'he392, 16'he393, 16'he394, 16'he395, 16'he396, 16'he397 	:	val_out <= 16'h2dbd;
         16'he398, 16'he399, 16'he39a, 16'he39b, 16'he39c, 16'he39d, 16'he39e, 16'he39f 	:	val_out <= 16'h2dd0;
         16'he3a0, 16'he3a1, 16'he3a2, 16'he3a3, 16'he3a4, 16'he3a5, 16'he3a6, 16'he3a7 	:	val_out <= 16'h2de3;
         16'he3a8, 16'he3a9, 16'he3aa, 16'he3ab, 16'he3ac, 16'he3ad, 16'he3ae, 16'he3af 	:	val_out <= 16'h2df7;
         16'he3b0, 16'he3b1, 16'he3b2, 16'he3b3, 16'he3b4, 16'he3b5, 16'he3b6, 16'he3b7 	:	val_out <= 16'h2e0a;
         16'he3b8, 16'he3b9, 16'he3ba, 16'he3bb, 16'he3bc, 16'he3bd, 16'he3be, 16'he3bf 	:	val_out <= 16'h2e1d;
         16'he3c0, 16'he3c1, 16'he3c2, 16'he3c3, 16'he3c4, 16'he3c5, 16'he3c6, 16'he3c7 	:	val_out <= 16'h2e31;
         16'he3c8, 16'he3c9, 16'he3ca, 16'he3cb, 16'he3cc, 16'he3cd, 16'he3ce, 16'he3cf 	:	val_out <= 16'h2e44;
         16'he3d0, 16'he3d1, 16'he3d2, 16'he3d3, 16'he3d4, 16'he3d5, 16'he3d6, 16'he3d7 	:	val_out <= 16'h2e57;
         16'he3d8, 16'he3d9, 16'he3da, 16'he3db, 16'he3dc, 16'he3dd, 16'he3de, 16'he3df 	:	val_out <= 16'h2e6b;
         16'he3e0, 16'he3e1, 16'he3e2, 16'he3e3, 16'he3e4, 16'he3e5, 16'he3e6, 16'he3e7 	:	val_out <= 16'h2e7e;
         16'he3e8, 16'he3e9, 16'he3ea, 16'he3eb, 16'he3ec, 16'he3ed, 16'he3ee, 16'he3ef 	:	val_out <= 16'h2e91;
         16'he3f0, 16'he3f1, 16'he3f2, 16'he3f3, 16'he3f4, 16'he3f5, 16'he3f6, 16'he3f7 	:	val_out <= 16'h2ea5;
         16'he3f8, 16'he3f9, 16'he3fa, 16'he3fb, 16'he3fc, 16'he3fd, 16'he3fe, 16'he3ff 	:	val_out <= 16'h2eb8;
         16'he400, 16'he401, 16'he402, 16'he403, 16'he404, 16'he405, 16'he406, 16'he407 	:	val_out <= 16'h2ecc;
         16'he408, 16'he409, 16'he40a, 16'he40b, 16'he40c, 16'he40d, 16'he40e, 16'he40f 	:	val_out <= 16'h2edf;
         16'he410, 16'he411, 16'he412, 16'he413, 16'he414, 16'he415, 16'he416, 16'he417 	:	val_out <= 16'h2ef3;
         16'he418, 16'he419, 16'he41a, 16'he41b, 16'he41c, 16'he41d, 16'he41e, 16'he41f 	:	val_out <= 16'h2f06;
         16'he420, 16'he421, 16'he422, 16'he423, 16'he424, 16'he425, 16'he426, 16'he427 	:	val_out <= 16'h2f1a;
         16'he428, 16'he429, 16'he42a, 16'he42b, 16'he42c, 16'he42d, 16'he42e, 16'he42f 	:	val_out <= 16'h2f2d;
         16'he430, 16'he431, 16'he432, 16'he433, 16'he434, 16'he435, 16'he436, 16'he437 	:	val_out <= 16'h2f40;
         16'he438, 16'he439, 16'he43a, 16'he43b, 16'he43c, 16'he43d, 16'he43e, 16'he43f 	:	val_out <= 16'h2f54;
         16'he440, 16'he441, 16'he442, 16'he443, 16'he444, 16'he445, 16'he446, 16'he447 	:	val_out <= 16'h2f68;
         16'he448, 16'he449, 16'he44a, 16'he44b, 16'he44c, 16'he44d, 16'he44e, 16'he44f 	:	val_out <= 16'h2f7b;
         16'he450, 16'he451, 16'he452, 16'he453, 16'he454, 16'he455, 16'he456, 16'he457 	:	val_out <= 16'h2f8f;
         16'he458, 16'he459, 16'he45a, 16'he45b, 16'he45c, 16'he45d, 16'he45e, 16'he45f 	:	val_out <= 16'h2fa2;
         16'he460, 16'he461, 16'he462, 16'he463, 16'he464, 16'he465, 16'he466, 16'he467 	:	val_out <= 16'h2fb6;
         16'he468, 16'he469, 16'he46a, 16'he46b, 16'he46c, 16'he46d, 16'he46e, 16'he46f 	:	val_out <= 16'h2fc9;
         16'he470, 16'he471, 16'he472, 16'he473, 16'he474, 16'he475, 16'he476, 16'he477 	:	val_out <= 16'h2fdd;
         16'he478, 16'he479, 16'he47a, 16'he47b, 16'he47c, 16'he47d, 16'he47e, 16'he47f 	:	val_out <= 16'h2ff0;
         16'he480, 16'he481, 16'he482, 16'he483, 16'he484, 16'he485, 16'he486, 16'he487 	:	val_out <= 16'h3004;
         16'he488, 16'he489, 16'he48a, 16'he48b, 16'he48c, 16'he48d, 16'he48e, 16'he48f 	:	val_out <= 16'h3018;
         16'he490, 16'he491, 16'he492, 16'he493, 16'he494, 16'he495, 16'he496, 16'he497 	:	val_out <= 16'h302b;
         16'he498, 16'he499, 16'he49a, 16'he49b, 16'he49c, 16'he49d, 16'he49e, 16'he49f 	:	val_out <= 16'h303f;
         16'he4a0, 16'he4a1, 16'he4a2, 16'he4a3, 16'he4a4, 16'he4a5, 16'he4a6, 16'he4a7 	:	val_out <= 16'h3053;
         16'he4a8, 16'he4a9, 16'he4aa, 16'he4ab, 16'he4ac, 16'he4ad, 16'he4ae, 16'he4af 	:	val_out <= 16'h3066;
         16'he4b0, 16'he4b1, 16'he4b2, 16'he4b3, 16'he4b4, 16'he4b5, 16'he4b6, 16'he4b7 	:	val_out <= 16'h307a;
         16'he4b8, 16'he4b9, 16'he4ba, 16'he4bb, 16'he4bc, 16'he4bd, 16'he4be, 16'he4bf 	:	val_out <= 16'h308e;
         16'he4c0, 16'he4c1, 16'he4c2, 16'he4c3, 16'he4c4, 16'he4c5, 16'he4c6, 16'he4c7 	:	val_out <= 16'h30a1;
         16'he4c8, 16'he4c9, 16'he4ca, 16'he4cb, 16'he4cc, 16'he4cd, 16'he4ce, 16'he4cf 	:	val_out <= 16'h30b5;
         16'he4d0, 16'he4d1, 16'he4d2, 16'he4d3, 16'he4d4, 16'he4d5, 16'he4d6, 16'he4d7 	:	val_out <= 16'h30c9;
         16'he4d8, 16'he4d9, 16'he4da, 16'he4db, 16'he4dc, 16'he4dd, 16'he4de, 16'he4df 	:	val_out <= 16'h30dd;
         16'he4e0, 16'he4e1, 16'he4e2, 16'he4e3, 16'he4e4, 16'he4e5, 16'he4e6, 16'he4e7 	:	val_out <= 16'h30f0;
         16'he4e8, 16'he4e9, 16'he4ea, 16'he4eb, 16'he4ec, 16'he4ed, 16'he4ee, 16'he4ef 	:	val_out <= 16'h3104;
         16'he4f0, 16'he4f1, 16'he4f2, 16'he4f3, 16'he4f4, 16'he4f5, 16'he4f6, 16'he4f7 	:	val_out <= 16'h3118;
         16'he4f8, 16'he4f9, 16'he4fa, 16'he4fb, 16'he4fc, 16'he4fd, 16'he4fe, 16'he4ff 	:	val_out <= 16'h312c;
         16'he500, 16'he501, 16'he502, 16'he503, 16'he504, 16'he505, 16'he506, 16'he507 	:	val_out <= 16'h3140;
         16'he508, 16'he509, 16'he50a, 16'he50b, 16'he50c, 16'he50d, 16'he50e, 16'he50f 	:	val_out <= 16'h3153;
         16'he510, 16'he511, 16'he512, 16'he513, 16'he514, 16'he515, 16'he516, 16'he517 	:	val_out <= 16'h3167;
         16'he518, 16'he519, 16'he51a, 16'he51b, 16'he51c, 16'he51d, 16'he51e, 16'he51f 	:	val_out <= 16'h317b;
         16'he520, 16'he521, 16'he522, 16'he523, 16'he524, 16'he525, 16'he526, 16'he527 	:	val_out <= 16'h318f;
         16'he528, 16'he529, 16'he52a, 16'he52b, 16'he52c, 16'he52d, 16'he52e, 16'he52f 	:	val_out <= 16'h31a3;
         16'he530, 16'he531, 16'he532, 16'he533, 16'he534, 16'he535, 16'he536, 16'he537 	:	val_out <= 16'h31b7;
         16'he538, 16'he539, 16'he53a, 16'he53b, 16'he53c, 16'he53d, 16'he53e, 16'he53f 	:	val_out <= 16'h31cb;
         16'he540, 16'he541, 16'he542, 16'he543, 16'he544, 16'he545, 16'he546, 16'he547 	:	val_out <= 16'h31de;
         16'he548, 16'he549, 16'he54a, 16'he54b, 16'he54c, 16'he54d, 16'he54e, 16'he54f 	:	val_out <= 16'h31f2;
         16'he550, 16'he551, 16'he552, 16'he553, 16'he554, 16'he555, 16'he556, 16'he557 	:	val_out <= 16'h3206;
         16'he558, 16'he559, 16'he55a, 16'he55b, 16'he55c, 16'he55d, 16'he55e, 16'he55f 	:	val_out <= 16'h321a;
         16'he560, 16'he561, 16'he562, 16'he563, 16'he564, 16'he565, 16'he566, 16'he567 	:	val_out <= 16'h322e;
         16'he568, 16'he569, 16'he56a, 16'he56b, 16'he56c, 16'he56d, 16'he56e, 16'he56f 	:	val_out <= 16'h3242;
         16'he570, 16'he571, 16'he572, 16'he573, 16'he574, 16'he575, 16'he576, 16'he577 	:	val_out <= 16'h3256;
         16'he578, 16'he579, 16'he57a, 16'he57b, 16'he57c, 16'he57d, 16'he57e, 16'he57f 	:	val_out <= 16'h326a;
         16'he580, 16'he581, 16'he582, 16'he583, 16'he584, 16'he585, 16'he586, 16'he587 	:	val_out <= 16'h327e;
         16'he588, 16'he589, 16'he58a, 16'he58b, 16'he58c, 16'he58d, 16'he58e, 16'he58f 	:	val_out <= 16'h3292;
         16'he590, 16'he591, 16'he592, 16'he593, 16'he594, 16'he595, 16'he596, 16'he597 	:	val_out <= 16'h32a6;
         16'he598, 16'he599, 16'he59a, 16'he59b, 16'he59c, 16'he59d, 16'he59e, 16'he59f 	:	val_out <= 16'h32ba;
         16'he5a0, 16'he5a1, 16'he5a2, 16'he5a3, 16'he5a4, 16'he5a5, 16'he5a6, 16'he5a7 	:	val_out <= 16'h32ce;
         16'he5a8, 16'he5a9, 16'he5aa, 16'he5ab, 16'he5ac, 16'he5ad, 16'he5ae, 16'he5af 	:	val_out <= 16'h32e2;
         16'he5b0, 16'he5b1, 16'he5b2, 16'he5b3, 16'he5b4, 16'he5b5, 16'he5b6, 16'he5b7 	:	val_out <= 16'h32f6;
         16'he5b8, 16'he5b9, 16'he5ba, 16'he5bb, 16'he5bc, 16'he5bd, 16'he5be, 16'he5bf 	:	val_out <= 16'h330a;
         16'he5c0, 16'he5c1, 16'he5c2, 16'he5c3, 16'he5c4, 16'he5c5, 16'he5c6, 16'he5c7 	:	val_out <= 16'h331e;
         16'he5c8, 16'he5c9, 16'he5ca, 16'he5cb, 16'he5cc, 16'he5cd, 16'he5ce, 16'he5cf 	:	val_out <= 16'h3333;
         16'he5d0, 16'he5d1, 16'he5d2, 16'he5d3, 16'he5d4, 16'he5d5, 16'he5d6, 16'he5d7 	:	val_out <= 16'h3347;
         16'he5d8, 16'he5d9, 16'he5da, 16'he5db, 16'he5dc, 16'he5dd, 16'he5de, 16'he5df 	:	val_out <= 16'h335b;
         16'he5e0, 16'he5e1, 16'he5e2, 16'he5e3, 16'he5e4, 16'he5e5, 16'he5e6, 16'he5e7 	:	val_out <= 16'h336f;
         16'he5e8, 16'he5e9, 16'he5ea, 16'he5eb, 16'he5ec, 16'he5ed, 16'he5ee, 16'he5ef 	:	val_out <= 16'h3383;
         16'he5f0, 16'he5f1, 16'he5f2, 16'he5f3, 16'he5f4, 16'he5f5, 16'he5f6, 16'he5f7 	:	val_out <= 16'h3397;
         16'he5f8, 16'he5f9, 16'he5fa, 16'he5fb, 16'he5fc, 16'he5fd, 16'he5fe, 16'he5ff 	:	val_out <= 16'h33ab;
         16'he600, 16'he601, 16'he602, 16'he603, 16'he604, 16'he605, 16'he606, 16'he607 	:	val_out <= 16'h33c0;
         16'he608, 16'he609, 16'he60a, 16'he60b, 16'he60c, 16'he60d, 16'he60e, 16'he60f 	:	val_out <= 16'h33d4;
         16'he610, 16'he611, 16'he612, 16'he613, 16'he614, 16'he615, 16'he616, 16'he617 	:	val_out <= 16'h33e8;
         16'he618, 16'he619, 16'he61a, 16'he61b, 16'he61c, 16'he61d, 16'he61e, 16'he61f 	:	val_out <= 16'h33fc;
         16'he620, 16'he621, 16'he622, 16'he623, 16'he624, 16'he625, 16'he626, 16'he627 	:	val_out <= 16'h3410;
         16'he628, 16'he629, 16'he62a, 16'he62b, 16'he62c, 16'he62d, 16'he62e, 16'he62f 	:	val_out <= 16'h3425;
         16'he630, 16'he631, 16'he632, 16'he633, 16'he634, 16'he635, 16'he636, 16'he637 	:	val_out <= 16'h3439;
         16'he638, 16'he639, 16'he63a, 16'he63b, 16'he63c, 16'he63d, 16'he63e, 16'he63f 	:	val_out <= 16'h344d;
         16'he640, 16'he641, 16'he642, 16'he643, 16'he644, 16'he645, 16'he646, 16'he647 	:	val_out <= 16'h3461;
         16'he648, 16'he649, 16'he64a, 16'he64b, 16'he64c, 16'he64d, 16'he64e, 16'he64f 	:	val_out <= 16'h3476;
         16'he650, 16'he651, 16'he652, 16'he653, 16'he654, 16'he655, 16'he656, 16'he657 	:	val_out <= 16'h348a;
         16'he658, 16'he659, 16'he65a, 16'he65b, 16'he65c, 16'he65d, 16'he65e, 16'he65f 	:	val_out <= 16'h349e;
         16'he660, 16'he661, 16'he662, 16'he663, 16'he664, 16'he665, 16'he666, 16'he667 	:	val_out <= 16'h34b3;
         16'he668, 16'he669, 16'he66a, 16'he66b, 16'he66c, 16'he66d, 16'he66e, 16'he66f 	:	val_out <= 16'h34c7;
         16'he670, 16'he671, 16'he672, 16'he673, 16'he674, 16'he675, 16'he676, 16'he677 	:	val_out <= 16'h34db;
         16'he678, 16'he679, 16'he67a, 16'he67b, 16'he67c, 16'he67d, 16'he67e, 16'he67f 	:	val_out <= 16'h34f0;
         16'he680, 16'he681, 16'he682, 16'he683, 16'he684, 16'he685, 16'he686, 16'he687 	:	val_out <= 16'h3504;
         16'he688, 16'he689, 16'he68a, 16'he68b, 16'he68c, 16'he68d, 16'he68e, 16'he68f 	:	val_out <= 16'h3518;
         16'he690, 16'he691, 16'he692, 16'he693, 16'he694, 16'he695, 16'he696, 16'he697 	:	val_out <= 16'h352d;
         16'he698, 16'he699, 16'he69a, 16'he69b, 16'he69c, 16'he69d, 16'he69e, 16'he69f 	:	val_out <= 16'h3541;
         16'he6a0, 16'he6a1, 16'he6a2, 16'he6a3, 16'he6a4, 16'he6a5, 16'he6a6, 16'he6a7 	:	val_out <= 16'h3556;
         16'he6a8, 16'he6a9, 16'he6aa, 16'he6ab, 16'he6ac, 16'he6ad, 16'he6ae, 16'he6af 	:	val_out <= 16'h356a;
         16'he6b0, 16'he6b1, 16'he6b2, 16'he6b3, 16'he6b4, 16'he6b5, 16'he6b6, 16'he6b7 	:	val_out <= 16'h357e;
         16'he6b8, 16'he6b9, 16'he6ba, 16'he6bb, 16'he6bc, 16'he6bd, 16'he6be, 16'he6bf 	:	val_out <= 16'h3593;
         16'he6c0, 16'he6c1, 16'he6c2, 16'he6c3, 16'he6c4, 16'he6c5, 16'he6c6, 16'he6c7 	:	val_out <= 16'h35a7;
         16'he6c8, 16'he6c9, 16'he6ca, 16'he6cb, 16'he6cc, 16'he6cd, 16'he6ce, 16'he6cf 	:	val_out <= 16'h35bc;
         16'he6d0, 16'he6d1, 16'he6d2, 16'he6d3, 16'he6d4, 16'he6d5, 16'he6d6, 16'he6d7 	:	val_out <= 16'h35d0;
         16'he6d8, 16'he6d9, 16'he6da, 16'he6db, 16'he6dc, 16'he6dd, 16'he6de, 16'he6df 	:	val_out <= 16'h35e5;
         16'he6e0, 16'he6e1, 16'he6e2, 16'he6e3, 16'he6e4, 16'he6e5, 16'he6e6, 16'he6e7 	:	val_out <= 16'h35f9;
         16'he6e8, 16'he6e9, 16'he6ea, 16'he6eb, 16'he6ec, 16'he6ed, 16'he6ee, 16'he6ef 	:	val_out <= 16'h360e;
         16'he6f0, 16'he6f1, 16'he6f2, 16'he6f3, 16'he6f4, 16'he6f5, 16'he6f6, 16'he6f7 	:	val_out <= 16'h3622;
         16'he6f8, 16'he6f9, 16'he6fa, 16'he6fb, 16'he6fc, 16'he6fd, 16'he6fe, 16'he6ff 	:	val_out <= 16'h3637;
         16'he700, 16'he701, 16'he702, 16'he703, 16'he704, 16'he705, 16'he706, 16'he707 	:	val_out <= 16'h364b;
         16'he708, 16'he709, 16'he70a, 16'he70b, 16'he70c, 16'he70d, 16'he70e, 16'he70f 	:	val_out <= 16'h3660;
         16'he710, 16'he711, 16'he712, 16'he713, 16'he714, 16'he715, 16'he716, 16'he717 	:	val_out <= 16'h3675;
         16'he718, 16'he719, 16'he71a, 16'he71b, 16'he71c, 16'he71d, 16'he71e, 16'he71f 	:	val_out <= 16'h3689;
         16'he720, 16'he721, 16'he722, 16'he723, 16'he724, 16'he725, 16'he726, 16'he727 	:	val_out <= 16'h369e;
         16'he728, 16'he729, 16'he72a, 16'he72b, 16'he72c, 16'he72d, 16'he72e, 16'he72f 	:	val_out <= 16'h36b2;
         16'he730, 16'he731, 16'he732, 16'he733, 16'he734, 16'he735, 16'he736, 16'he737 	:	val_out <= 16'h36c7;
         16'he738, 16'he739, 16'he73a, 16'he73b, 16'he73c, 16'he73d, 16'he73e, 16'he73f 	:	val_out <= 16'h36dc;
         16'he740, 16'he741, 16'he742, 16'he743, 16'he744, 16'he745, 16'he746, 16'he747 	:	val_out <= 16'h36f0;
         16'he748, 16'he749, 16'he74a, 16'he74b, 16'he74c, 16'he74d, 16'he74e, 16'he74f 	:	val_out <= 16'h3705;
         16'he750, 16'he751, 16'he752, 16'he753, 16'he754, 16'he755, 16'he756, 16'he757 	:	val_out <= 16'h3719;
         16'he758, 16'he759, 16'he75a, 16'he75b, 16'he75c, 16'he75d, 16'he75e, 16'he75f 	:	val_out <= 16'h372e;
         16'he760, 16'he761, 16'he762, 16'he763, 16'he764, 16'he765, 16'he766, 16'he767 	:	val_out <= 16'h3743;
         16'he768, 16'he769, 16'he76a, 16'he76b, 16'he76c, 16'he76d, 16'he76e, 16'he76f 	:	val_out <= 16'h3757;
         16'he770, 16'he771, 16'he772, 16'he773, 16'he774, 16'he775, 16'he776, 16'he777 	:	val_out <= 16'h376c;
         16'he778, 16'he779, 16'he77a, 16'he77b, 16'he77c, 16'he77d, 16'he77e, 16'he77f 	:	val_out <= 16'h3781;
         16'he780, 16'he781, 16'he782, 16'he783, 16'he784, 16'he785, 16'he786, 16'he787 	:	val_out <= 16'h3796;
         16'he788, 16'he789, 16'he78a, 16'he78b, 16'he78c, 16'he78d, 16'he78e, 16'he78f 	:	val_out <= 16'h37aa;
         16'he790, 16'he791, 16'he792, 16'he793, 16'he794, 16'he795, 16'he796, 16'he797 	:	val_out <= 16'h37bf;
         16'he798, 16'he799, 16'he79a, 16'he79b, 16'he79c, 16'he79d, 16'he79e, 16'he79f 	:	val_out <= 16'h37d4;
         16'he7a0, 16'he7a1, 16'he7a2, 16'he7a3, 16'he7a4, 16'he7a5, 16'he7a6, 16'he7a7 	:	val_out <= 16'h37e9;
         16'he7a8, 16'he7a9, 16'he7aa, 16'he7ab, 16'he7ac, 16'he7ad, 16'he7ae, 16'he7af 	:	val_out <= 16'h37fd;
         16'he7b0, 16'he7b1, 16'he7b2, 16'he7b3, 16'he7b4, 16'he7b5, 16'he7b6, 16'he7b7 	:	val_out <= 16'h3812;
         16'he7b8, 16'he7b9, 16'he7ba, 16'he7bb, 16'he7bc, 16'he7bd, 16'he7be, 16'he7bf 	:	val_out <= 16'h3827;
         16'he7c0, 16'he7c1, 16'he7c2, 16'he7c3, 16'he7c4, 16'he7c5, 16'he7c6, 16'he7c7 	:	val_out <= 16'h383c;
         16'he7c8, 16'he7c9, 16'he7ca, 16'he7cb, 16'he7cc, 16'he7cd, 16'he7ce, 16'he7cf 	:	val_out <= 16'h3851;
         16'he7d0, 16'he7d1, 16'he7d2, 16'he7d3, 16'he7d4, 16'he7d5, 16'he7d6, 16'he7d7 	:	val_out <= 16'h3865;
         16'he7d8, 16'he7d9, 16'he7da, 16'he7db, 16'he7dc, 16'he7dd, 16'he7de, 16'he7df 	:	val_out <= 16'h387a;
         16'he7e0, 16'he7e1, 16'he7e2, 16'he7e3, 16'he7e4, 16'he7e5, 16'he7e6, 16'he7e7 	:	val_out <= 16'h388f;
         16'he7e8, 16'he7e9, 16'he7ea, 16'he7eb, 16'he7ec, 16'he7ed, 16'he7ee, 16'he7ef 	:	val_out <= 16'h38a4;
         16'he7f0, 16'he7f1, 16'he7f2, 16'he7f3, 16'he7f4, 16'he7f5, 16'he7f6, 16'he7f7 	:	val_out <= 16'h38b9;
         16'he7f8, 16'he7f9, 16'he7fa, 16'he7fb, 16'he7fc, 16'he7fd, 16'he7fe, 16'he7ff 	:	val_out <= 16'h38ce;
         16'he800, 16'he801, 16'he802, 16'he803, 16'he804, 16'he805, 16'he806, 16'he807 	:	val_out <= 16'h38e3;
         16'he808, 16'he809, 16'he80a, 16'he80b, 16'he80c, 16'he80d, 16'he80e, 16'he80f 	:	val_out <= 16'h38f7;
         16'he810, 16'he811, 16'he812, 16'he813, 16'he814, 16'he815, 16'he816, 16'he817 	:	val_out <= 16'h390c;
         16'he818, 16'he819, 16'he81a, 16'he81b, 16'he81c, 16'he81d, 16'he81e, 16'he81f 	:	val_out <= 16'h3921;
         16'he820, 16'he821, 16'he822, 16'he823, 16'he824, 16'he825, 16'he826, 16'he827 	:	val_out <= 16'h3936;
         16'he828, 16'he829, 16'he82a, 16'he82b, 16'he82c, 16'he82d, 16'he82e, 16'he82f 	:	val_out <= 16'h394b;
         16'he830, 16'he831, 16'he832, 16'he833, 16'he834, 16'he835, 16'he836, 16'he837 	:	val_out <= 16'h3960;
         16'he838, 16'he839, 16'he83a, 16'he83b, 16'he83c, 16'he83d, 16'he83e, 16'he83f 	:	val_out <= 16'h3975;
         16'he840, 16'he841, 16'he842, 16'he843, 16'he844, 16'he845, 16'he846, 16'he847 	:	val_out <= 16'h398a;
         16'he848, 16'he849, 16'he84a, 16'he84b, 16'he84c, 16'he84d, 16'he84e, 16'he84f 	:	val_out <= 16'h399f;
         16'he850, 16'he851, 16'he852, 16'he853, 16'he854, 16'he855, 16'he856, 16'he857 	:	val_out <= 16'h39b4;
         16'he858, 16'he859, 16'he85a, 16'he85b, 16'he85c, 16'he85d, 16'he85e, 16'he85f 	:	val_out <= 16'h39c9;
         16'he860, 16'he861, 16'he862, 16'he863, 16'he864, 16'he865, 16'he866, 16'he867 	:	val_out <= 16'h39de;
         16'he868, 16'he869, 16'he86a, 16'he86b, 16'he86c, 16'he86d, 16'he86e, 16'he86f 	:	val_out <= 16'h39f3;
         16'he870, 16'he871, 16'he872, 16'he873, 16'he874, 16'he875, 16'he876, 16'he877 	:	val_out <= 16'h3a08;
         16'he878, 16'he879, 16'he87a, 16'he87b, 16'he87c, 16'he87d, 16'he87e, 16'he87f 	:	val_out <= 16'h3a1d;
         16'he880, 16'he881, 16'he882, 16'he883, 16'he884, 16'he885, 16'he886, 16'he887 	:	val_out <= 16'h3a32;
         16'he888, 16'he889, 16'he88a, 16'he88b, 16'he88c, 16'he88d, 16'he88e, 16'he88f 	:	val_out <= 16'h3a47;
         16'he890, 16'he891, 16'he892, 16'he893, 16'he894, 16'he895, 16'he896, 16'he897 	:	val_out <= 16'h3a5c;
         16'he898, 16'he899, 16'he89a, 16'he89b, 16'he89c, 16'he89d, 16'he89e, 16'he89f 	:	val_out <= 16'h3a72;
         16'he8a0, 16'he8a1, 16'he8a2, 16'he8a3, 16'he8a4, 16'he8a5, 16'he8a6, 16'he8a7 	:	val_out <= 16'h3a87;
         16'he8a8, 16'he8a9, 16'he8aa, 16'he8ab, 16'he8ac, 16'he8ad, 16'he8ae, 16'he8af 	:	val_out <= 16'h3a9c;
         16'he8b0, 16'he8b1, 16'he8b2, 16'he8b3, 16'he8b4, 16'he8b5, 16'he8b6, 16'he8b7 	:	val_out <= 16'h3ab1;
         16'he8b8, 16'he8b9, 16'he8ba, 16'he8bb, 16'he8bc, 16'he8bd, 16'he8be, 16'he8bf 	:	val_out <= 16'h3ac6;
         16'he8c0, 16'he8c1, 16'he8c2, 16'he8c3, 16'he8c4, 16'he8c5, 16'he8c6, 16'he8c7 	:	val_out <= 16'h3adb;
         16'he8c8, 16'he8c9, 16'he8ca, 16'he8cb, 16'he8cc, 16'he8cd, 16'he8ce, 16'he8cf 	:	val_out <= 16'h3af0;
         16'he8d0, 16'he8d1, 16'he8d2, 16'he8d3, 16'he8d4, 16'he8d5, 16'he8d6, 16'he8d7 	:	val_out <= 16'h3b05;
         16'he8d8, 16'he8d9, 16'he8da, 16'he8db, 16'he8dc, 16'he8dd, 16'he8de, 16'he8df 	:	val_out <= 16'h3b1b;
         16'he8e0, 16'he8e1, 16'he8e2, 16'he8e3, 16'he8e4, 16'he8e5, 16'he8e6, 16'he8e7 	:	val_out <= 16'h3b30;
         16'he8e8, 16'he8e9, 16'he8ea, 16'he8eb, 16'he8ec, 16'he8ed, 16'he8ee, 16'he8ef 	:	val_out <= 16'h3b45;
         16'he8f0, 16'he8f1, 16'he8f2, 16'he8f3, 16'he8f4, 16'he8f5, 16'he8f6, 16'he8f7 	:	val_out <= 16'h3b5a;
         16'he8f8, 16'he8f9, 16'he8fa, 16'he8fb, 16'he8fc, 16'he8fd, 16'he8fe, 16'he8ff 	:	val_out <= 16'h3b6f;
         16'he900, 16'he901, 16'he902, 16'he903, 16'he904, 16'he905, 16'he906, 16'he907 	:	val_out <= 16'h3b85;
         16'he908, 16'he909, 16'he90a, 16'he90b, 16'he90c, 16'he90d, 16'he90e, 16'he90f 	:	val_out <= 16'h3b9a;
         16'he910, 16'he911, 16'he912, 16'he913, 16'he914, 16'he915, 16'he916, 16'he917 	:	val_out <= 16'h3baf;
         16'he918, 16'he919, 16'he91a, 16'he91b, 16'he91c, 16'he91d, 16'he91e, 16'he91f 	:	val_out <= 16'h3bc4;
         16'he920, 16'he921, 16'he922, 16'he923, 16'he924, 16'he925, 16'he926, 16'he927 	:	val_out <= 16'h3bda;
         16'he928, 16'he929, 16'he92a, 16'he92b, 16'he92c, 16'he92d, 16'he92e, 16'he92f 	:	val_out <= 16'h3bef;
         16'he930, 16'he931, 16'he932, 16'he933, 16'he934, 16'he935, 16'he936, 16'he937 	:	val_out <= 16'h3c04;
         16'he938, 16'he939, 16'he93a, 16'he93b, 16'he93c, 16'he93d, 16'he93e, 16'he93f 	:	val_out <= 16'h3c1a;
         16'he940, 16'he941, 16'he942, 16'he943, 16'he944, 16'he945, 16'he946, 16'he947 	:	val_out <= 16'h3c2f;
         16'he948, 16'he949, 16'he94a, 16'he94b, 16'he94c, 16'he94d, 16'he94e, 16'he94f 	:	val_out <= 16'h3c44;
         16'he950, 16'he951, 16'he952, 16'he953, 16'he954, 16'he955, 16'he956, 16'he957 	:	val_out <= 16'h3c5a;
         16'he958, 16'he959, 16'he95a, 16'he95b, 16'he95c, 16'he95d, 16'he95e, 16'he95f 	:	val_out <= 16'h3c6f;
         16'he960, 16'he961, 16'he962, 16'he963, 16'he964, 16'he965, 16'he966, 16'he967 	:	val_out <= 16'h3c84;
         16'he968, 16'he969, 16'he96a, 16'he96b, 16'he96c, 16'he96d, 16'he96e, 16'he96f 	:	val_out <= 16'h3c9a;
         16'he970, 16'he971, 16'he972, 16'he973, 16'he974, 16'he975, 16'he976, 16'he977 	:	val_out <= 16'h3caf;
         16'he978, 16'he979, 16'he97a, 16'he97b, 16'he97c, 16'he97d, 16'he97e, 16'he97f 	:	val_out <= 16'h3cc4;
         16'he980, 16'he981, 16'he982, 16'he983, 16'he984, 16'he985, 16'he986, 16'he987 	:	val_out <= 16'h3cda;
         16'he988, 16'he989, 16'he98a, 16'he98b, 16'he98c, 16'he98d, 16'he98e, 16'he98f 	:	val_out <= 16'h3cef;
         16'he990, 16'he991, 16'he992, 16'he993, 16'he994, 16'he995, 16'he996, 16'he997 	:	val_out <= 16'h3d05;
         16'he998, 16'he999, 16'he99a, 16'he99b, 16'he99c, 16'he99d, 16'he99e, 16'he99f 	:	val_out <= 16'h3d1a;
         16'he9a0, 16'he9a1, 16'he9a2, 16'he9a3, 16'he9a4, 16'he9a5, 16'he9a6, 16'he9a7 	:	val_out <= 16'h3d2f;
         16'he9a8, 16'he9a9, 16'he9aa, 16'he9ab, 16'he9ac, 16'he9ad, 16'he9ae, 16'he9af 	:	val_out <= 16'h3d45;
         16'he9b0, 16'he9b1, 16'he9b2, 16'he9b3, 16'he9b4, 16'he9b5, 16'he9b6, 16'he9b7 	:	val_out <= 16'h3d5a;
         16'he9b8, 16'he9b9, 16'he9ba, 16'he9bb, 16'he9bc, 16'he9bd, 16'he9be, 16'he9bf 	:	val_out <= 16'h3d70;
         16'he9c0, 16'he9c1, 16'he9c2, 16'he9c3, 16'he9c4, 16'he9c5, 16'he9c6, 16'he9c7 	:	val_out <= 16'h3d85;
         16'he9c8, 16'he9c9, 16'he9ca, 16'he9cb, 16'he9cc, 16'he9cd, 16'he9ce, 16'he9cf 	:	val_out <= 16'h3d9b;
         16'he9d0, 16'he9d1, 16'he9d2, 16'he9d3, 16'he9d4, 16'he9d5, 16'he9d6, 16'he9d7 	:	val_out <= 16'h3db0;
         16'he9d8, 16'he9d9, 16'he9da, 16'he9db, 16'he9dc, 16'he9dd, 16'he9de, 16'he9df 	:	val_out <= 16'h3dc6;
         16'he9e0, 16'he9e1, 16'he9e2, 16'he9e3, 16'he9e4, 16'he9e5, 16'he9e6, 16'he9e7 	:	val_out <= 16'h3ddb;
         16'he9e8, 16'he9e9, 16'he9ea, 16'he9eb, 16'he9ec, 16'he9ed, 16'he9ee, 16'he9ef 	:	val_out <= 16'h3df1;
         16'he9f0, 16'he9f1, 16'he9f2, 16'he9f3, 16'he9f4, 16'he9f5, 16'he9f6, 16'he9f7 	:	val_out <= 16'h3e06;
         16'he9f8, 16'he9f9, 16'he9fa, 16'he9fb, 16'he9fc, 16'he9fd, 16'he9fe, 16'he9ff 	:	val_out <= 16'h3e1c;
         16'hea00, 16'hea01, 16'hea02, 16'hea03, 16'hea04, 16'hea05, 16'hea06, 16'hea07 	:	val_out <= 16'h3e31;
         16'hea08, 16'hea09, 16'hea0a, 16'hea0b, 16'hea0c, 16'hea0d, 16'hea0e, 16'hea0f 	:	val_out <= 16'h3e47;
         16'hea10, 16'hea11, 16'hea12, 16'hea13, 16'hea14, 16'hea15, 16'hea16, 16'hea17 	:	val_out <= 16'h3e5d;
         16'hea18, 16'hea19, 16'hea1a, 16'hea1b, 16'hea1c, 16'hea1d, 16'hea1e, 16'hea1f 	:	val_out <= 16'h3e72;
         16'hea20, 16'hea21, 16'hea22, 16'hea23, 16'hea24, 16'hea25, 16'hea26, 16'hea27 	:	val_out <= 16'h3e88;
         16'hea28, 16'hea29, 16'hea2a, 16'hea2b, 16'hea2c, 16'hea2d, 16'hea2e, 16'hea2f 	:	val_out <= 16'h3e9d;
         16'hea30, 16'hea31, 16'hea32, 16'hea33, 16'hea34, 16'hea35, 16'hea36, 16'hea37 	:	val_out <= 16'h3eb3;
         16'hea38, 16'hea39, 16'hea3a, 16'hea3b, 16'hea3c, 16'hea3d, 16'hea3e, 16'hea3f 	:	val_out <= 16'h3ec9;
         16'hea40, 16'hea41, 16'hea42, 16'hea43, 16'hea44, 16'hea45, 16'hea46, 16'hea47 	:	val_out <= 16'h3ede;
         16'hea48, 16'hea49, 16'hea4a, 16'hea4b, 16'hea4c, 16'hea4d, 16'hea4e, 16'hea4f 	:	val_out <= 16'h3ef4;
         16'hea50, 16'hea51, 16'hea52, 16'hea53, 16'hea54, 16'hea55, 16'hea56, 16'hea57 	:	val_out <= 16'h3f09;
         16'hea58, 16'hea59, 16'hea5a, 16'hea5b, 16'hea5c, 16'hea5d, 16'hea5e, 16'hea5f 	:	val_out <= 16'h3f1f;
         16'hea60, 16'hea61, 16'hea62, 16'hea63, 16'hea64, 16'hea65, 16'hea66, 16'hea67 	:	val_out <= 16'h3f35;
         16'hea68, 16'hea69, 16'hea6a, 16'hea6b, 16'hea6c, 16'hea6d, 16'hea6e, 16'hea6f 	:	val_out <= 16'h3f4a;
         16'hea70, 16'hea71, 16'hea72, 16'hea73, 16'hea74, 16'hea75, 16'hea76, 16'hea77 	:	val_out <= 16'h3f60;
         16'hea78, 16'hea79, 16'hea7a, 16'hea7b, 16'hea7c, 16'hea7d, 16'hea7e, 16'hea7f 	:	val_out <= 16'h3f76;
         16'hea80, 16'hea81, 16'hea82, 16'hea83, 16'hea84, 16'hea85, 16'hea86, 16'hea87 	:	val_out <= 16'h3f8c;
         16'hea88, 16'hea89, 16'hea8a, 16'hea8b, 16'hea8c, 16'hea8d, 16'hea8e, 16'hea8f 	:	val_out <= 16'h3fa1;
         16'hea90, 16'hea91, 16'hea92, 16'hea93, 16'hea94, 16'hea95, 16'hea96, 16'hea97 	:	val_out <= 16'h3fb7;
         16'hea98, 16'hea99, 16'hea9a, 16'hea9b, 16'hea9c, 16'hea9d, 16'hea9e, 16'hea9f 	:	val_out <= 16'h3fcd;
         16'heaa0, 16'heaa1, 16'heaa2, 16'heaa3, 16'heaa4, 16'heaa5, 16'heaa6, 16'heaa7 	:	val_out <= 16'h3fe2;
         16'heaa8, 16'heaa9, 16'heaaa, 16'heaab, 16'heaac, 16'heaad, 16'heaae, 16'heaaf 	:	val_out <= 16'h3ff8;
         16'heab0, 16'heab1, 16'heab2, 16'heab3, 16'heab4, 16'heab5, 16'heab6, 16'heab7 	:	val_out <= 16'h400e;
         16'heab8, 16'heab9, 16'heaba, 16'heabb, 16'heabc, 16'heabd, 16'heabe, 16'heabf 	:	val_out <= 16'h4024;
         16'heac0, 16'heac1, 16'heac2, 16'heac3, 16'heac4, 16'heac5, 16'heac6, 16'heac7 	:	val_out <= 16'h403a;
         16'heac8, 16'heac9, 16'heaca, 16'heacb, 16'heacc, 16'heacd, 16'heace, 16'heacf 	:	val_out <= 16'h404f;
         16'head0, 16'head1, 16'head2, 16'head3, 16'head4, 16'head5, 16'head6, 16'head7 	:	val_out <= 16'h4065;
         16'head8, 16'head9, 16'heada, 16'headb, 16'headc, 16'headd, 16'heade, 16'headf 	:	val_out <= 16'h407b;
         16'heae0, 16'heae1, 16'heae2, 16'heae3, 16'heae4, 16'heae5, 16'heae6, 16'heae7 	:	val_out <= 16'h4091;
         16'heae8, 16'heae9, 16'heaea, 16'heaeb, 16'heaec, 16'heaed, 16'heaee, 16'heaef 	:	val_out <= 16'h40a7;
         16'heaf0, 16'heaf1, 16'heaf2, 16'heaf3, 16'heaf4, 16'heaf5, 16'heaf6, 16'heaf7 	:	val_out <= 16'h40bc;
         16'heaf8, 16'heaf9, 16'heafa, 16'heafb, 16'heafc, 16'heafd, 16'heafe, 16'heaff 	:	val_out <= 16'h40d2;
         16'heb00, 16'heb01, 16'heb02, 16'heb03, 16'heb04, 16'heb05, 16'heb06, 16'heb07 	:	val_out <= 16'h40e8;
         16'heb08, 16'heb09, 16'heb0a, 16'heb0b, 16'heb0c, 16'heb0d, 16'heb0e, 16'heb0f 	:	val_out <= 16'h40fe;
         16'heb10, 16'heb11, 16'heb12, 16'heb13, 16'heb14, 16'heb15, 16'heb16, 16'heb17 	:	val_out <= 16'h4114;
         16'heb18, 16'heb19, 16'heb1a, 16'heb1b, 16'heb1c, 16'heb1d, 16'heb1e, 16'heb1f 	:	val_out <= 16'h412a;
         16'heb20, 16'heb21, 16'heb22, 16'heb23, 16'heb24, 16'heb25, 16'heb26, 16'heb27 	:	val_out <= 16'h4140;
         16'heb28, 16'heb29, 16'heb2a, 16'heb2b, 16'heb2c, 16'heb2d, 16'heb2e, 16'heb2f 	:	val_out <= 16'h4156;
         16'heb30, 16'heb31, 16'heb32, 16'heb33, 16'heb34, 16'heb35, 16'heb36, 16'heb37 	:	val_out <= 16'h416c;
         16'heb38, 16'heb39, 16'heb3a, 16'heb3b, 16'heb3c, 16'heb3d, 16'heb3e, 16'heb3f 	:	val_out <= 16'h4182;
         16'heb40, 16'heb41, 16'heb42, 16'heb43, 16'heb44, 16'heb45, 16'heb46, 16'heb47 	:	val_out <= 16'h4197;
         16'heb48, 16'heb49, 16'heb4a, 16'heb4b, 16'heb4c, 16'heb4d, 16'heb4e, 16'heb4f 	:	val_out <= 16'h41ad;
         16'heb50, 16'heb51, 16'heb52, 16'heb53, 16'heb54, 16'heb55, 16'heb56, 16'heb57 	:	val_out <= 16'h41c3;
         16'heb58, 16'heb59, 16'heb5a, 16'heb5b, 16'heb5c, 16'heb5d, 16'heb5e, 16'heb5f 	:	val_out <= 16'h41d9;
         16'heb60, 16'heb61, 16'heb62, 16'heb63, 16'heb64, 16'heb65, 16'heb66, 16'heb67 	:	val_out <= 16'h41ef;
         16'heb68, 16'heb69, 16'heb6a, 16'heb6b, 16'heb6c, 16'heb6d, 16'heb6e, 16'heb6f 	:	val_out <= 16'h4205;
         16'heb70, 16'heb71, 16'heb72, 16'heb73, 16'heb74, 16'heb75, 16'heb76, 16'heb77 	:	val_out <= 16'h421b;
         16'heb78, 16'heb79, 16'heb7a, 16'heb7b, 16'heb7c, 16'heb7d, 16'heb7e, 16'heb7f 	:	val_out <= 16'h4231;
         16'heb80, 16'heb81, 16'heb82, 16'heb83, 16'heb84, 16'heb85, 16'heb86, 16'heb87 	:	val_out <= 16'h4247;
         16'heb88, 16'heb89, 16'heb8a, 16'heb8b, 16'heb8c, 16'heb8d, 16'heb8e, 16'heb8f 	:	val_out <= 16'h425d;
         16'heb90, 16'heb91, 16'heb92, 16'heb93, 16'heb94, 16'heb95, 16'heb96, 16'heb97 	:	val_out <= 16'h4273;
         16'heb98, 16'heb99, 16'heb9a, 16'heb9b, 16'heb9c, 16'heb9d, 16'heb9e, 16'heb9f 	:	val_out <= 16'h4289;
         16'heba0, 16'heba1, 16'heba2, 16'heba3, 16'heba4, 16'heba5, 16'heba6, 16'heba7 	:	val_out <= 16'h429f;
         16'heba8, 16'heba9, 16'hebaa, 16'hebab, 16'hebac, 16'hebad, 16'hebae, 16'hebaf 	:	val_out <= 16'h42b6;
         16'hebb0, 16'hebb1, 16'hebb2, 16'hebb3, 16'hebb4, 16'hebb5, 16'hebb6, 16'hebb7 	:	val_out <= 16'h42cc;
         16'hebb8, 16'hebb9, 16'hebba, 16'hebbb, 16'hebbc, 16'hebbd, 16'hebbe, 16'hebbf 	:	val_out <= 16'h42e2;
         16'hebc0, 16'hebc1, 16'hebc2, 16'hebc3, 16'hebc4, 16'hebc5, 16'hebc6, 16'hebc7 	:	val_out <= 16'h42f8;
         16'hebc8, 16'hebc9, 16'hebca, 16'hebcb, 16'hebcc, 16'hebcd, 16'hebce, 16'hebcf 	:	val_out <= 16'h430e;
         16'hebd0, 16'hebd1, 16'hebd2, 16'hebd3, 16'hebd4, 16'hebd5, 16'hebd6, 16'hebd7 	:	val_out <= 16'h4324;
         16'hebd8, 16'hebd9, 16'hebda, 16'hebdb, 16'hebdc, 16'hebdd, 16'hebde, 16'hebdf 	:	val_out <= 16'h433a;
         16'hebe0, 16'hebe1, 16'hebe2, 16'hebe3, 16'hebe4, 16'hebe5, 16'hebe6, 16'hebe7 	:	val_out <= 16'h4350;
         16'hebe8, 16'hebe9, 16'hebea, 16'hebeb, 16'hebec, 16'hebed, 16'hebee, 16'hebef 	:	val_out <= 16'h4366;
         16'hebf0, 16'hebf1, 16'hebf2, 16'hebf3, 16'hebf4, 16'hebf5, 16'hebf6, 16'hebf7 	:	val_out <= 16'h437c;
         16'hebf8, 16'hebf9, 16'hebfa, 16'hebfb, 16'hebfc, 16'hebfd, 16'hebfe, 16'hebff 	:	val_out <= 16'h4393;
         16'hec00, 16'hec01, 16'hec02, 16'hec03, 16'hec04, 16'hec05, 16'hec06, 16'hec07 	:	val_out <= 16'h43a9;
         16'hec08, 16'hec09, 16'hec0a, 16'hec0b, 16'hec0c, 16'hec0d, 16'hec0e, 16'hec0f 	:	val_out <= 16'h43bf;
         16'hec10, 16'hec11, 16'hec12, 16'hec13, 16'hec14, 16'hec15, 16'hec16, 16'hec17 	:	val_out <= 16'h43d5;
         16'hec18, 16'hec19, 16'hec1a, 16'hec1b, 16'hec1c, 16'hec1d, 16'hec1e, 16'hec1f 	:	val_out <= 16'h43eb;
         16'hec20, 16'hec21, 16'hec22, 16'hec23, 16'hec24, 16'hec25, 16'hec26, 16'hec27 	:	val_out <= 16'h4402;
         16'hec28, 16'hec29, 16'hec2a, 16'hec2b, 16'hec2c, 16'hec2d, 16'hec2e, 16'hec2f 	:	val_out <= 16'h4418;
         16'hec30, 16'hec31, 16'hec32, 16'hec33, 16'hec34, 16'hec35, 16'hec36, 16'hec37 	:	val_out <= 16'h442e;
         16'hec38, 16'hec39, 16'hec3a, 16'hec3b, 16'hec3c, 16'hec3d, 16'hec3e, 16'hec3f 	:	val_out <= 16'h4444;
         16'hec40, 16'hec41, 16'hec42, 16'hec43, 16'hec44, 16'hec45, 16'hec46, 16'hec47 	:	val_out <= 16'h445a;
         16'hec48, 16'hec49, 16'hec4a, 16'hec4b, 16'hec4c, 16'hec4d, 16'hec4e, 16'hec4f 	:	val_out <= 16'h4471;
         16'hec50, 16'hec51, 16'hec52, 16'hec53, 16'hec54, 16'hec55, 16'hec56, 16'hec57 	:	val_out <= 16'h4487;
         16'hec58, 16'hec59, 16'hec5a, 16'hec5b, 16'hec5c, 16'hec5d, 16'hec5e, 16'hec5f 	:	val_out <= 16'h449d;
         16'hec60, 16'hec61, 16'hec62, 16'hec63, 16'hec64, 16'hec65, 16'hec66, 16'hec67 	:	val_out <= 16'h44b3;
         16'hec68, 16'hec69, 16'hec6a, 16'hec6b, 16'hec6c, 16'hec6d, 16'hec6e, 16'hec6f 	:	val_out <= 16'h44ca;
         16'hec70, 16'hec71, 16'hec72, 16'hec73, 16'hec74, 16'hec75, 16'hec76, 16'hec77 	:	val_out <= 16'h44e0;
         16'hec78, 16'hec79, 16'hec7a, 16'hec7b, 16'hec7c, 16'hec7d, 16'hec7e, 16'hec7f 	:	val_out <= 16'h44f6;
         16'hec80, 16'hec81, 16'hec82, 16'hec83, 16'hec84, 16'hec85, 16'hec86, 16'hec87 	:	val_out <= 16'h450d;
         16'hec88, 16'hec89, 16'hec8a, 16'hec8b, 16'hec8c, 16'hec8d, 16'hec8e, 16'hec8f 	:	val_out <= 16'h4523;
         16'hec90, 16'hec91, 16'hec92, 16'hec93, 16'hec94, 16'hec95, 16'hec96, 16'hec97 	:	val_out <= 16'h4539;
         16'hec98, 16'hec99, 16'hec9a, 16'hec9b, 16'hec9c, 16'hec9d, 16'hec9e, 16'hec9f 	:	val_out <= 16'h4550;
         16'heca0, 16'heca1, 16'heca2, 16'heca3, 16'heca4, 16'heca5, 16'heca6, 16'heca7 	:	val_out <= 16'h4566;
         16'heca8, 16'heca9, 16'hecaa, 16'hecab, 16'hecac, 16'hecad, 16'hecae, 16'hecaf 	:	val_out <= 16'h457c;
         16'hecb0, 16'hecb1, 16'hecb2, 16'hecb3, 16'hecb4, 16'hecb5, 16'hecb6, 16'hecb7 	:	val_out <= 16'h4593;
         16'hecb8, 16'hecb9, 16'hecba, 16'hecbb, 16'hecbc, 16'hecbd, 16'hecbe, 16'hecbf 	:	val_out <= 16'h45a9;
         16'hecc0, 16'hecc1, 16'hecc2, 16'hecc3, 16'hecc4, 16'hecc5, 16'hecc6, 16'hecc7 	:	val_out <= 16'h45bf;
         16'hecc8, 16'hecc9, 16'hecca, 16'heccb, 16'heccc, 16'heccd, 16'hecce, 16'heccf 	:	val_out <= 16'h45d6;
         16'hecd0, 16'hecd1, 16'hecd2, 16'hecd3, 16'hecd4, 16'hecd5, 16'hecd6, 16'hecd7 	:	val_out <= 16'h45ec;
         16'hecd8, 16'hecd9, 16'hecda, 16'hecdb, 16'hecdc, 16'hecdd, 16'hecde, 16'hecdf 	:	val_out <= 16'h4602;
         16'hece0, 16'hece1, 16'hece2, 16'hece3, 16'hece4, 16'hece5, 16'hece6, 16'hece7 	:	val_out <= 16'h4619;
         16'hece8, 16'hece9, 16'hecea, 16'heceb, 16'hecec, 16'heced, 16'hecee, 16'hecef 	:	val_out <= 16'h462f;
         16'hecf0, 16'hecf1, 16'hecf2, 16'hecf3, 16'hecf4, 16'hecf5, 16'hecf6, 16'hecf7 	:	val_out <= 16'h4646;
         16'hecf8, 16'hecf9, 16'hecfa, 16'hecfb, 16'hecfc, 16'hecfd, 16'hecfe, 16'hecff 	:	val_out <= 16'h465c;
         16'hed00, 16'hed01, 16'hed02, 16'hed03, 16'hed04, 16'hed05, 16'hed06, 16'hed07 	:	val_out <= 16'h4673;
         16'hed08, 16'hed09, 16'hed0a, 16'hed0b, 16'hed0c, 16'hed0d, 16'hed0e, 16'hed0f 	:	val_out <= 16'h4689;
         16'hed10, 16'hed11, 16'hed12, 16'hed13, 16'hed14, 16'hed15, 16'hed16, 16'hed17 	:	val_out <= 16'h46a0;
         16'hed18, 16'hed19, 16'hed1a, 16'hed1b, 16'hed1c, 16'hed1d, 16'hed1e, 16'hed1f 	:	val_out <= 16'h46b6;
         16'hed20, 16'hed21, 16'hed22, 16'hed23, 16'hed24, 16'hed25, 16'hed26, 16'hed27 	:	val_out <= 16'h46cd;
         16'hed28, 16'hed29, 16'hed2a, 16'hed2b, 16'hed2c, 16'hed2d, 16'hed2e, 16'hed2f 	:	val_out <= 16'h46e3;
         16'hed30, 16'hed31, 16'hed32, 16'hed33, 16'hed34, 16'hed35, 16'hed36, 16'hed37 	:	val_out <= 16'h46f9;
         16'hed38, 16'hed39, 16'hed3a, 16'hed3b, 16'hed3c, 16'hed3d, 16'hed3e, 16'hed3f 	:	val_out <= 16'h4710;
         16'hed40, 16'hed41, 16'hed42, 16'hed43, 16'hed44, 16'hed45, 16'hed46, 16'hed47 	:	val_out <= 16'h4727;
         16'hed48, 16'hed49, 16'hed4a, 16'hed4b, 16'hed4c, 16'hed4d, 16'hed4e, 16'hed4f 	:	val_out <= 16'h473d;
         16'hed50, 16'hed51, 16'hed52, 16'hed53, 16'hed54, 16'hed55, 16'hed56, 16'hed57 	:	val_out <= 16'h4754;
         16'hed58, 16'hed59, 16'hed5a, 16'hed5b, 16'hed5c, 16'hed5d, 16'hed5e, 16'hed5f 	:	val_out <= 16'h476a;
         16'hed60, 16'hed61, 16'hed62, 16'hed63, 16'hed64, 16'hed65, 16'hed66, 16'hed67 	:	val_out <= 16'h4781;
         16'hed68, 16'hed69, 16'hed6a, 16'hed6b, 16'hed6c, 16'hed6d, 16'hed6e, 16'hed6f 	:	val_out <= 16'h4797;
         16'hed70, 16'hed71, 16'hed72, 16'hed73, 16'hed74, 16'hed75, 16'hed76, 16'hed77 	:	val_out <= 16'h47ae;
         16'hed78, 16'hed79, 16'hed7a, 16'hed7b, 16'hed7c, 16'hed7d, 16'hed7e, 16'hed7f 	:	val_out <= 16'h47c4;
         16'hed80, 16'hed81, 16'hed82, 16'hed83, 16'hed84, 16'hed85, 16'hed86, 16'hed87 	:	val_out <= 16'h47db;
         16'hed88, 16'hed89, 16'hed8a, 16'hed8b, 16'hed8c, 16'hed8d, 16'hed8e, 16'hed8f 	:	val_out <= 16'h47f2;
         16'hed90, 16'hed91, 16'hed92, 16'hed93, 16'hed94, 16'hed95, 16'hed96, 16'hed97 	:	val_out <= 16'h4808;
         16'hed98, 16'hed99, 16'hed9a, 16'hed9b, 16'hed9c, 16'hed9d, 16'hed9e, 16'hed9f 	:	val_out <= 16'h481f;
         16'heda0, 16'heda1, 16'heda2, 16'heda3, 16'heda4, 16'heda5, 16'heda6, 16'heda7 	:	val_out <= 16'h4835;
         16'heda8, 16'heda9, 16'hedaa, 16'hedab, 16'hedac, 16'hedad, 16'hedae, 16'hedaf 	:	val_out <= 16'h484c;
         16'hedb0, 16'hedb1, 16'hedb2, 16'hedb3, 16'hedb4, 16'hedb5, 16'hedb6, 16'hedb7 	:	val_out <= 16'h4863;
         16'hedb8, 16'hedb9, 16'hedba, 16'hedbb, 16'hedbc, 16'hedbd, 16'hedbe, 16'hedbf 	:	val_out <= 16'h4879;
         16'hedc0, 16'hedc1, 16'hedc2, 16'hedc3, 16'hedc4, 16'hedc5, 16'hedc6, 16'hedc7 	:	val_out <= 16'h4890;
         16'hedc8, 16'hedc9, 16'hedca, 16'hedcb, 16'hedcc, 16'hedcd, 16'hedce, 16'hedcf 	:	val_out <= 16'h48a7;
         16'hedd0, 16'hedd1, 16'hedd2, 16'hedd3, 16'hedd4, 16'hedd5, 16'hedd6, 16'hedd7 	:	val_out <= 16'h48bd;
         16'hedd8, 16'hedd9, 16'hedda, 16'heddb, 16'heddc, 16'heddd, 16'hedde, 16'heddf 	:	val_out <= 16'h48d4;
         16'hede0, 16'hede1, 16'hede2, 16'hede3, 16'hede4, 16'hede5, 16'hede6, 16'hede7 	:	val_out <= 16'h48eb;
         16'hede8, 16'hede9, 16'hedea, 16'hedeb, 16'hedec, 16'heded, 16'hedee, 16'hedef 	:	val_out <= 16'h4901;
         16'hedf0, 16'hedf1, 16'hedf2, 16'hedf3, 16'hedf4, 16'hedf5, 16'hedf6, 16'hedf7 	:	val_out <= 16'h4918;
         16'hedf8, 16'hedf9, 16'hedfa, 16'hedfb, 16'hedfc, 16'hedfd, 16'hedfe, 16'hedff 	:	val_out <= 16'h492f;
         16'hee00, 16'hee01, 16'hee02, 16'hee03, 16'hee04, 16'hee05, 16'hee06, 16'hee07 	:	val_out <= 16'h4945;
         16'hee08, 16'hee09, 16'hee0a, 16'hee0b, 16'hee0c, 16'hee0d, 16'hee0e, 16'hee0f 	:	val_out <= 16'h495c;
         16'hee10, 16'hee11, 16'hee12, 16'hee13, 16'hee14, 16'hee15, 16'hee16, 16'hee17 	:	val_out <= 16'h4973;
         16'hee18, 16'hee19, 16'hee1a, 16'hee1b, 16'hee1c, 16'hee1d, 16'hee1e, 16'hee1f 	:	val_out <= 16'h498a;
         16'hee20, 16'hee21, 16'hee22, 16'hee23, 16'hee24, 16'hee25, 16'hee26, 16'hee27 	:	val_out <= 16'h49a0;
         16'hee28, 16'hee29, 16'hee2a, 16'hee2b, 16'hee2c, 16'hee2d, 16'hee2e, 16'hee2f 	:	val_out <= 16'h49b7;
         16'hee30, 16'hee31, 16'hee32, 16'hee33, 16'hee34, 16'hee35, 16'hee36, 16'hee37 	:	val_out <= 16'h49ce;
         16'hee38, 16'hee39, 16'hee3a, 16'hee3b, 16'hee3c, 16'hee3d, 16'hee3e, 16'hee3f 	:	val_out <= 16'h49e5;
         16'hee40, 16'hee41, 16'hee42, 16'hee43, 16'hee44, 16'hee45, 16'hee46, 16'hee47 	:	val_out <= 16'h49fb;
         16'hee48, 16'hee49, 16'hee4a, 16'hee4b, 16'hee4c, 16'hee4d, 16'hee4e, 16'hee4f 	:	val_out <= 16'h4a12;
         16'hee50, 16'hee51, 16'hee52, 16'hee53, 16'hee54, 16'hee55, 16'hee56, 16'hee57 	:	val_out <= 16'h4a29;
         16'hee58, 16'hee59, 16'hee5a, 16'hee5b, 16'hee5c, 16'hee5d, 16'hee5e, 16'hee5f 	:	val_out <= 16'h4a40;
         16'hee60, 16'hee61, 16'hee62, 16'hee63, 16'hee64, 16'hee65, 16'hee66, 16'hee67 	:	val_out <= 16'h4a57;
         16'hee68, 16'hee69, 16'hee6a, 16'hee6b, 16'hee6c, 16'hee6d, 16'hee6e, 16'hee6f 	:	val_out <= 16'h4a6d;
         16'hee70, 16'hee71, 16'hee72, 16'hee73, 16'hee74, 16'hee75, 16'hee76, 16'hee77 	:	val_out <= 16'h4a84;
         16'hee78, 16'hee79, 16'hee7a, 16'hee7b, 16'hee7c, 16'hee7d, 16'hee7e, 16'hee7f 	:	val_out <= 16'h4a9b;
         16'hee80, 16'hee81, 16'hee82, 16'hee83, 16'hee84, 16'hee85, 16'hee86, 16'hee87 	:	val_out <= 16'h4ab2;
         16'hee88, 16'hee89, 16'hee8a, 16'hee8b, 16'hee8c, 16'hee8d, 16'hee8e, 16'hee8f 	:	val_out <= 16'h4ac9;
         16'hee90, 16'hee91, 16'hee92, 16'hee93, 16'hee94, 16'hee95, 16'hee96, 16'hee97 	:	val_out <= 16'h4ae0;
         16'hee98, 16'hee99, 16'hee9a, 16'hee9b, 16'hee9c, 16'hee9d, 16'hee9e, 16'hee9f 	:	val_out <= 16'h4af7;
         16'heea0, 16'heea1, 16'heea2, 16'heea3, 16'heea4, 16'heea5, 16'heea6, 16'heea7 	:	val_out <= 16'h4b0d;
         16'heea8, 16'heea9, 16'heeaa, 16'heeab, 16'heeac, 16'heead, 16'heeae, 16'heeaf 	:	val_out <= 16'h4b24;
         16'heeb0, 16'heeb1, 16'heeb2, 16'heeb3, 16'heeb4, 16'heeb5, 16'heeb6, 16'heeb7 	:	val_out <= 16'h4b3b;
         16'heeb8, 16'heeb9, 16'heeba, 16'heebb, 16'heebc, 16'heebd, 16'heebe, 16'heebf 	:	val_out <= 16'h4b52;
         16'heec0, 16'heec1, 16'heec2, 16'heec3, 16'heec4, 16'heec5, 16'heec6, 16'heec7 	:	val_out <= 16'h4b69;
         16'heec8, 16'heec9, 16'heeca, 16'heecb, 16'heecc, 16'heecd, 16'heece, 16'heecf 	:	val_out <= 16'h4b80;
         16'heed0, 16'heed1, 16'heed2, 16'heed3, 16'heed4, 16'heed5, 16'heed6, 16'heed7 	:	val_out <= 16'h4b97;
         16'heed8, 16'heed9, 16'heeda, 16'heedb, 16'heedc, 16'heedd, 16'heede, 16'heedf 	:	val_out <= 16'h4bae;
         16'heee0, 16'heee1, 16'heee2, 16'heee3, 16'heee4, 16'heee5, 16'heee6, 16'heee7 	:	val_out <= 16'h4bc5;
         16'heee8, 16'heee9, 16'heeea, 16'heeeb, 16'heeec, 16'heeed, 16'heeee, 16'heeef 	:	val_out <= 16'h4bdc;
         16'heef0, 16'heef1, 16'heef2, 16'heef3, 16'heef4, 16'heef5, 16'heef6, 16'heef7 	:	val_out <= 16'h4bf3;
         16'heef8, 16'heef9, 16'heefa, 16'heefb, 16'heefc, 16'heefd, 16'heefe, 16'heeff 	:	val_out <= 16'h4c0a;
         16'hef00, 16'hef01, 16'hef02, 16'hef03, 16'hef04, 16'hef05, 16'hef06, 16'hef07 	:	val_out <= 16'h4c21;
         16'hef08, 16'hef09, 16'hef0a, 16'hef0b, 16'hef0c, 16'hef0d, 16'hef0e, 16'hef0f 	:	val_out <= 16'h4c38;
         16'hef10, 16'hef11, 16'hef12, 16'hef13, 16'hef14, 16'hef15, 16'hef16, 16'hef17 	:	val_out <= 16'h4c4f;
         16'hef18, 16'hef19, 16'hef1a, 16'hef1b, 16'hef1c, 16'hef1d, 16'hef1e, 16'hef1f 	:	val_out <= 16'h4c66;
         16'hef20, 16'hef21, 16'hef22, 16'hef23, 16'hef24, 16'hef25, 16'hef26, 16'hef27 	:	val_out <= 16'h4c7d;
         16'hef28, 16'hef29, 16'hef2a, 16'hef2b, 16'hef2c, 16'hef2d, 16'hef2e, 16'hef2f 	:	val_out <= 16'h4c94;
         16'hef30, 16'hef31, 16'hef32, 16'hef33, 16'hef34, 16'hef35, 16'hef36, 16'hef37 	:	val_out <= 16'h4cab;
         16'hef38, 16'hef39, 16'hef3a, 16'hef3b, 16'hef3c, 16'hef3d, 16'hef3e, 16'hef3f 	:	val_out <= 16'h4cc2;
         16'hef40, 16'hef41, 16'hef42, 16'hef43, 16'hef44, 16'hef45, 16'hef46, 16'hef47 	:	val_out <= 16'h4cd9;
         16'hef48, 16'hef49, 16'hef4a, 16'hef4b, 16'hef4c, 16'hef4d, 16'hef4e, 16'hef4f 	:	val_out <= 16'h4cf0;
         16'hef50, 16'hef51, 16'hef52, 16'hef53, 16'hef54, 16'hef55, 16'hef56, 16'hef57 	:	val_out <= 16'h4d07;
         16'hef58, 16'hef59, 16'hef5a, 16'hef5b, 16'hef5c, 16'hef5d, 16'hef5e, 16'hef5f 	:	val_out <= 16'h4d1e;
         16'hef60, 16'hef61, 16'hef62, 16'hef63, 16'hef64, 16'hef65, 16'hef66, 16'hef67 	:	val_out <= 16'h4d35;
         16'hef68, 16'hef69, 16'hef6a, 16'hef6b, 16'hef6c, 16'hef6d, 16'hef6e, 16'hef6f 	:	val_out <= 16'h4d4c;
         16'hef70, 16'hef71, 16'hef72, 16'hef73, 16'hef74, 16'hef75, 16'hef76, 16'hef77 	:	val_out <= 16'h4d63;
         16'hef78, 16'hef79, 16'hef7a, 16'hef7b, 16'hef7c, 16'hef7d, 16'hef7e, 16'hef7f 	:	val_out <= 16'h4d7a;
         16'hef80, 16'hef81, 16'hef82, 16'hef83, 16'hef84, 16'hef85, 16'hef86, 16'hef87 	:	val_out <= 16'h4d91;
         16'hef88, 16'hef89, 16'hef8a, 16'hef8b, 16'hef8c, 16'hef8d, 16'hef8e, 16'hef8f 	:	val_out <= 16'h4da8;
         16'hef90, 16'hef91, 16'hef92, 16'hef93, 16'hef94, 16'hef95, 16'hef96, 16'hef97 	:	val_out <= 16'h4dbf;
         16'hef98, 16'hef99, 16'hef9a, 16'hef9b, 16'hef9c, 16'hef9d, 16'hef9e, 16'hef9f 	:	val_out <= 16'h4dd7;
         16'hefa0, 16'hefa1, 16'hefa2, 16'hefa3, 16'hefa4, 16'hefa5, 16'hefa6, 16'hefa7 	:	val_out <= 16'h4dee;
         16'hefa8, 16'hefa9, 16'hefaa, 16'hefab, 16'hefac, 16'hefad, 16'hefae, 16'hefaf 	:	val_out <= 16'h4e05;
         16'hefb0, 16'hefb1, 16'hefb2, 16'hefb3, 16'hefb4, 16'hefb5, 16'hefb6, 16'hefb7 	:	val_out <= 16'h4e1c;
         16'hefb8, 16'hefb9, 16'hefba, 16'hefbb, 16'hefbc, 16'hefbd, 16'hefbe, 16'hefbf 	:	val_out <= 16'h4e33;
         16'hefc0, 16'hefc1, 16'hefc2, 16'hefc3, 16'hefc4, 16'hefc5, 16'hefc6, 16'hefc7 	:	val_out <= 16'h4e4a;
         16'hefc8, 16'hefc9, 16'hefca, 16'hefcb, 16'hefcc, 16'hefcd, 16'hefce, 16'hefcf 	:	val_out <= 16'h4e61;
         16'hefd0, 16'hefd1, 16'hefd2, 16'hefd3, 16'hefd4, 16'hefd5, 16'hefd6, 16'hefd7 	:	val_out <= 16'h4e79;
         16'hefd8, 16'hefd9, 16'hefda, 16'hefdb, 16'hefdc, 16'hefdd, 16'hefde, 16'hefdf 	:	val_out <= 16'h4e90;
         16'hefe0, 16'hefe1, 16'hefe2, 16'hefe3, 16'hefe4, 16'hefe5, 16'hefe6, 16'hefe7 	:	val_out <= 16'h4ea7;
         16'hefe8, 16'hefe9, 16'hefea, 16'hefeb, 16'hefec, 16'hefed, 16'hefee, 16'hefef 	:	val_out <= 16'h4ebe;
         16'heff0, 16'heff1, 16'heff2, 16'heff3, 16'heff4, 16'heff5, 16'heff6, 16'heff7 	:	val_out <= 16'h4ed5;
         16'heff8, 16'heff9, 16'heffa, 16'heffb, 16'heffc, 16'heffd, 16'heffe, 16'hefff 	:	val_out <= 16'h4eed;
         16'hf000, 16'hf001, 16'hf002, 16'hf003, 16'hf004, 16'hf005, 16'hf006, 16'hf007 	:	val_out <= 16'h4f04;
         16'hf008, 16'hf009, 16'hf00a, 16'hf00b, 16'hf00c, 16'hf00d, 16'hf00e, 16'hf00f 	:	val_out <= 16'h4f1b;
         16'hf010, 16'hf011, 16'hf012, 16'hf013, 16'hf014, 16'hf015, 16'hf016, 16'hf017 	:	val_out <= 16'h4f32;
         16'hf018, 16'hf019, 16'hf01a, 16'hf01b, 16'hf01c, 16'hf01d, 16'hf01e, 16'hf01f 	:	val_out <= 16'h4f49;
         16'hf020, 16'hf021, 16'hf022, 16'hf023, 16'hf024, 16'hf025, 16'hf026, 16'hf027 	:	val_out <= 16'h4f61;
         16'hf028, 16'hf029, 16'hf02a, 16'hf02b, 16'hf02c, 16'hf02d, 16'hf02e, 16'hf02f 	:	val_out <= 16'h4f78;
         16'hf030, 16'hf031, 16'hf032, 16'hf033, 16'hf034, 16'hf035, 16'hf036, 16'hf037 	:	val_out <= 16'h4f8f;
         16'hf038, 16'hf039, 16'hf03a, 16'hf03b, 16'hf03c, 16'hf03d, 16'hf03e, 16'hf03f 	:	val_out <= 16'h4fa6;
         16'hf040, 16'hf041, 16'hf042, 16'hf043, 16'hf044, 16'hf045, 16'hf046, 16'hf047 	:	val_out <= 16'h4fbe;
         16'hf048, 16'hf049, 16'hf04a, 16'hf04b, 16'hf04c, 16'hf04d, 16'hf04e, 16'hf04f 	:	val_out <= 16'h4fd5;
         16'hf050, 16'hf051, 16'hf052, 16'hf053, 16'hf054, 16'hf055, 16'hf056, 16'hf057 	:	val_out <= 16'h4fec;
         16'hf058, 16'hf059, 16'hf05a, 16'hf05b, 16'hf05c, 16'hf05d, 16'hf05e, 16'hf05f 	:	val_out <= 16'h5004;
         16'hf060, 16'hf061, 16'hf062, 16'hf063, 16'hf064, 16'hf065, 16'hf066, 16'hf067 	:	val_out <= 16'h501b;
         16'hf068, 16'hf069, 16'hf06a, 16'hf06b, 16'hf06c, 16'hf06d, 16'hf06e, 16'hf06f 	:	val_out <= 16'h5032;
         16'hf070, 16'hf071, 16'hf072, 16'hf073, 16'hf074, 16'hf075, 16'hf076, 16'hf077 	:	val_out <= 16'h504a;
         16'hf078, 16'hf079, 16'hf07a, 16'hf07b, 16'hf07c, 16'hf07d, 16'hf07e, 16'hf07f 	:	val_out <= 16'h5061;
         16'hf080, 16'hf081, 16'hf082, 16'hf083, 16'hf084, 16'hf085, 16'hf086, 16'hf087 	:	val_out <= 16'h5078;
         16'hf088, 16'hf089, 16'hf08a, 16'hf08b, 16'hf08c, 16'hf08d, 16'hf08e, 16'hf08f 	:	val_out <= 16'h5090;
         16'hf090, 16'hf091, 16'hf092, 16'hf093, 16'hf094, 16'hf095, 16'hf096, 16'hf097 	:	val_out <= 16'h50a7;
         16'hf098, 16'hf099, 16'hf09a, 16'hf09b, 16'hf09c, 16'hf09d, 16'hf09e, 16'hf09f 	:	val_out <= 16'h50be;
         16'hf0a0, 16'hf0a1, 16'hf0a2, 16'hf0a3, 16'hf0a4, 16'hf0a5, 16'hf0a6, 16'hf0a7 	:	val_out <= 16'h50d6;
         16'hf0a8, 16'hf0a9, 16'hf0aa, 16'hf0ab, 16'hf0ac, 16'hf0ad, 16'hf0ae, 16'hf0af 	:	val_out <= 16'h50ed;
         16'hf0b0, 16'hf0b1, 16'hf0b2, 16'hf0b3, 16'hf0b4, 16'hf0b5, 16'hf0b6, 16'hf0b7 	:	val_out <= 16'h5104;
         16'hf0b8, 16'hf0b9, 16'hf0ba, 16'hf0bb, 16'hf0bc, 16'hf0bd, 16'hf0be, 16'hf0bf 	:	val_out <= 16'h511c;
         16'hf0c0, 16'hf0c1, 16'hf0c2, 16'hf0c3, 16'hf0c4, 16'hf0c5, 16'hf0c6, 16'hf0c7 	:	val_out <= 16'h5133;
         16'hf0c8, 16'hf0c9, 16'hf0ca, 16'hf0cb, 16'hf0cc, 16'hf0cd, 16'hf0ce, 16'hf0cf 	:	val_out <= 16'h514a;
         16'hf0d0, 16'hf0d1, 16'hf0d2, 16'hf0d3, 16'hf0d4, 16'hf0d5, 16'hf0d6, 16'hf0d7 	:	val_out <= 16'h5162;
         16'hf0d8, 16'hf0d9, 16'hf0da, 16'hf0db, 16'hf0dc, 16'hf0dd, 16'hf0de, 16'hf0df 	:	val_out <= 16'h5179;
         16'hf0e0, 16'hf0e1, 16'hf0e2, 16'hf0e3, 16'hf0e4, 16'hf0e5, 16'hf0e6, 16'hf0e7 	:	val_out <= 16'h5191;
         16'hf0e8, 16'hf0e9, 16'hf0ea, 16'hf0eb, 16'hf0ec, 16'hf0ed, 16'hf0ee, 16'hf0ef 	:	val_out <= 16'h51a8;
         16'hf0f0, 16'hf0f1, 16'hf0f2, 16'hf0f3, 16'hf0f4, 16'hf0f5, 16'hf0f6, 16'hf0f7 	:	val_out <= 16'h51c0;
         16'hf0f8, 16'hf0f9, 16'hf0fa, 16'hf0fb, 16'hf0fc, 16'hf0fd, 16'hf0fe, 16'hf0ff 	:	val_out <= 16'h51d7;
         16'hf100, 16'hf101, 16'hf102, 16'hf103, 16'hf104, 16'hf105, 16'hf106, 16'hf107 	:	val_out <= 16'h51ee;
         16'hf108, 16'hf109, 16'hf10a, 16'hf10b, 16'hf10c, 16'hf10d, 16'hf10e, 16'hf10f 	:	val_out <= 16'h5206;
         16'hf110, 16'hf111, 16'hf112, 16'hf113, 16'hf114, 16'hf115, 16'hf116, 16'hf117 	:	val_out <= 16'h521d;
         16'hf118, 16'hf119, 16'hf11a, 16'hf11b, 16'hf11c, 16'hf11d, 16'hf11e, 16'hf11f 	:	val_out <= 16'h5235;
         16'hf120, 16'hf121, 16'hf122, 16'hf123, 16'hf124, 16'hf125, 16'hf126, 16'hf127 	:	val_out <= 16'h524c;
         16'hf128, 16'hf129, 16'hf12a, 16'hf12b, 16'hf12c, 16'hf12d, 16'hf12e, 16'hf12f 	:	val_out <= 16'h5264;
         16'hf130, 16'hf131, 16'hf132, 16'hf133, 16'hf134, 16'hf135, 16'hf136, 16'hf137 	:	val_out <= 16'h527b;
         16'hf138, 16'hf139, 16'hf13a, 16'hf13b, 16'hf13c, 16'hf13d, 16'hf13e, 16'hf13f 	:	val_out <= 16'h5293;
         16'hf140, 16'hf141, 16'hf142, 16'hf143, 16'hf144, 16'hf145, 16'hf146, 16'hf147 	:	val_out <= 16'h52aa;
         16'hf148, 16'hf149, 16'hf14a, 16'hf14b, 16'hf14c, 16'hf14d, 16'hf14e, 16'hf14f 	:	val_out <= 16'h52c2;
         16'hf150, 16'hf151, 16'hf152, 16'hf153, 16'hf154, 16'hf155, 16'hf156, 16'hf157 	:	val_out <= 16'h52d9;
         16'hf158, 16'hf159, 16'hf15a, 16'hf15b, 16'hf15c, 16'hf15d, 16'hf15e, 16'hf15f 	:	val_out <= 16'h52f1;
         16'hf160, 16'hf161, 16'hf162, 16'hf163, 16'hf164, 16'hf165, 16'hf166, 16'hf167 	:	val_out <= 16'h5308;
         16'hf168, 16'hf169, 16'hf16a, 16'hf16b, 16'hf16c, 16'hf16d, 16'hf16e, 16'hf16f 	:	val_out <= 16'h5320;
         16'hf170, 16'hf171, 16'hf172, 16'hf173, 16'hf174, 16'hf175, 16'hf176, 16'hf177 	:	val_out <= 16'h5337;
         16'hf178, 16'hf179, 16'hf17a, 16'hf17b, 16'hf17c, 16'hf17d, 16'hf17e, 16'hf17f 	:	val_out <= 16'h534f;
         16'hf180, 16'hf181, 16'hf182, 16'hf183, 16'hf184, 16'hf185, 16'hf186, 16'hf187 	:	val_out <= 16'h5367;
         16'hf188, 16'hf189, 16'hf18a, 16'hf18b, 16'hf18c, 16'hf18d, 16'hf18e, 16'hf18f 	:	val_out <= 16'h537e;
         16'hf190, 16'hf191, 16'hf192, 16'hf193, 16'hf194, 16'hf195, 16'hf196, 16'hf197 	:	val_out <= 16'h5396;
         16'hf198, 16'hf199, 16'hf19a, 16'hf19b, 16'hf19c, 16'hf19d, 16'hf19e, 16'hf19f 	:	val_out <= 16'h53ad;
         16'hf1a0, 16'hf1a1, 16'hf1a2, 16'hf1a3, 16'hf1a4, 16'hf1a5, 16'hf1a6, 16'hf1a7 	:	val_out <= 16'h53c5;
         16'hf1a8, 16'hf1a9, 16'hf1aa, 16'hf1ab, 16'hf1ac, 16'hf1ad, 16'hf1ae, 16'hf1af 	:	val_out <= 16'h53dc;
         16'hf1b0, 16'hf1b1, 16'hf1b2, 16'hf1b3, 16'hf1b4, 16'hf1b5, 16'hf1b6, 16'hf1b7 	:	val_out <= 16'h53f4;
         16'hf1b8, 16'hf1b9, 16'hf1ba, 16'hf1bb, 16'hf1bc, 16'hf1bd, 16'hf1be, 16'hf1bf 	:	val_out <= 16'h540c;
         16'hf1c0, 16'hf1c1, 16'hf1c2, 16'hf1c3, 16'hf1c4, 16'hf1c5, 16'hf1c6, 16'hf1c7 	:	val_out <= 16'h5423;
         16'hf1c8, 16'hf1c9, 16'hf1ca, 16'hf1cb, 16'hf1cc, 16'hf1cd, 16'hf1ce, 16'hf1cf 	:	val_out <= 16'h543b;
         16'hf1d0, 16'hf1d1, 16'hf1d2, 16'hf1d3, 16'hf1d4, 16'hf1d5, 16'hf1d6, 16'hf1d7 	:	val_out <= 16'h5452;
         16'hf1d8, 16'hf1d9, 16'hf1da, 16'hf1db, 16'hf1dc, 16'hf1dd, 16'hf1de, 16'hf1df 	:	val_out <= 16'h546a;
         16'hf1e0, 16'hf1e1, 16'hf1e2, 16'hf1e3, 16'hf1e4, 16'hf1e5, 16'hf1e6, 16'hf1e7 	:	val_out <= 16'h5482;
         16'hf1e8, 16'hf1e9, 16'hf1ea, 16'hf1eb, 16'hf1ec, 16'hf1ed, 16'hf1ee, 16'hf1ef 	:	val_out <= 16'h5499;
         16'hf1f0, 16'hf1f1, 16'hf1f2, 16'hf1f3, 16'hf1f4, 16'hf1f5, 16'hf1f6, 16'hf1f7 	:	val_out <= 16'h54b1;
         16'hf1f8, 16'hf1f9, 16'hf1fa, 16'hf1fb, 16'hf1fc, 16'hf1fd, 16'hf1fe, 16'hf1ff 	:	val_out <= 16'h54c9;
         16'hf200, 16'hf201, 16'hf202, 16'hf203, 16'hf204, 16'hf205, 16'hf206, 16'hf207 	:	val_out <= 16'h54e0;
         16'hf208, 16'hf209, 16'hf20a, 16'hf20b, 16'hf20c, 16'hf20d, 16'hf20e, 16'hf20f 	:	val_out <= 16'h54f8;
         16'hf210, 16'hf211, 16'hf212, 16'hf213, 16'hf214, 16'hf215, 16'hf216, 16'hf217 	:	val_out <= 16'h5510;
         16'hf218, 16'hf219, 16'hf21a, 16'hf21b, 16'hf21c, 16'hf21d, 16'hf21e, 16'hf21f 	:	val_out <= 16'h5527;
         16'hf220, 16'hf221, 16'hf222, 16'hf223, 16'hf224, 16'hf225, 16'hf226, 16'hf227 	:	val_out <= 16'h553f;
         16'hf228, 16'hf229, 16'hf22a, 16'hf22b, 16'hf22c, 16'hf22d, 16'hf22e, 16'hf22f 	:	val_out <= 16'h5557;
         16'hf230, 16'hf231, 16'hf232, 16'hf233, 16'hf234, 16'hf235, 16'hf236, 16'hf237 	:	val_out <= 16'h556e;
         16'hf238, 16'hf239, 16'hf23a, 16'hf23b, 16'hf23c, 16'hf23d, 16'hf23e, 16'hf23f 	:	val_out <= 16'h5586;
         16'hf240, 16'hf241, 16'hf242, 16'hf243, 16'hf244, 16'hf245, 16'hf246, 16'hf247 	:	val_out <= 16'h559e;
         16'hf248, 16'hf249, 16'hf24a, 16'hf24b, 16'hf24c, 16'hf24d, 16'hf24e, 16'hf24f 	:	val_out <= 16'h55b6;
         16'hf250, 16'hf251, 16'hf252, 16'hf253, 16'hf254, 16'hf255, 16'hf256, 16'hf257 	:	val_out <= 16'h55cd;
         16'hf258, 16'hf259, 16'hf25a, 16'hf25b, 16'hf25c, 16'hf25d, 16'hf25e, 16'hf25f 	:	val_out <= 16'h55e5;
         16'hf260, 16'hf261, 16'hf262, 16'hf263, 16'hf264, 16'hf265, 16'hf266, 16'hf267 	:	val_out <= 16'h55fd;
         16'hf268, 16'hf269, 16'hf26a, 16'hf26b, 16'hf26c, 16'hf26d, 16'hf26e, 16'hf26f 	:	val_out <= 16'h5614;
         16'hf270, 16'hf271, 16'hf272, 16'hf273, 16'hf274, 16'hf275, 16'hf276, 16'hf277 	:	val_out <= 16'h562c;
         16'hf278, 16'hf279, 16'hf27a, 16'hf27b, 16'hf27c, 16'hf27d, 16'hf27e, 16'hf27f 	:	val_out <= 16'h5644;
         16'hf280, 16'hf281, 16'hf282, 16'hf283, 16'hf284, 16'hf285, 16'hf286, 16'hf287 	:	val_out <= 16'h565c;
         16'hf288, 16'hf289, 16'hf28a, 16'hf28b, 16'hf28c, 16'hf28d, 16'hf28e, 16'hf28f 	:	val_out <= 16'h5674;
         16'hf290, 16'hf291, 16'hf292, 16'hf293, 16'hf294, 16'hf295, 16'hf296, 16'hf297 	:	val_out <= 16'h568b;
         16'hf298, 16'hf299, 16'hf29a, 16'hf29b, 16'hf29c, 16'hf29d, 16'hf29e, 16'hf29f 	:	val_out <= 16'h56a3;
         16'hf2a0, 16'hf2a1, 16'hf2a2, 16'hf2a3, 16'hf2a4, 16'hf2a5, 16'hf2a6, 16'hf2a7 	:	val_out <= 16'h56bb;
         16'hf2a8, 16'hf2a9, 16'hf2aa, 16'hf2ab, 16'hf2ac, 16'hf2ad, 16'hf2ae, 16'hf2af 	:	val_out <= 16'h56d3;
         16'hf2b0, 16'hf2b1, 16'hf2b2, 16'hf2b3, 16'hf2b4, 16'hf2b5, 16'hf2b6, 16'hf2b7 	:	val_out <= 16'h56ea;
         16'hf2b8, 16'hf2b9, 16'hf2ba, 16'hf2bb, 16'hf2bc, 16'hf2bd, 16'hf2be, 16'hf2bf 	:	val_out <= 16'h5702;
         16'hf2c0, 16'hf2c1, 16'hf2c2, 16'hf2c3, 16'hf2c4, 16'hf2c5, 16'hf2c6, 16'hf2c7 	:	val_out <= 16'h571a;
         16'hf2c8, 16'hf2c9, 16'hf2ca, 16'hf2cb, 16'hf2cc, 16'hf2cd, 16'hf2ce, 16'hf2cf 	:	val_out <= 16'h5732;
         16'hf2d0, 16'hf2d1, 16'hf2d2, 16'hf2d3, 16'hf2d4, 16'hf2d5, 16'hf2d6, 16'hf2d7 	:	val_out <= 16'h574a;
         16'hf2d8, 16'hf2d9, 16'hf2da, 16'hf2db, 16'hf2dc, 16'hf2dd, 16'hf2de, 16'hf2df 	:	val_out <= 16'h5762;
         16'hf2e0, 16'hf2e1, 16'hf2e2, 16'hf2e3, 16'hf2e4, 16'hf2e5, 16'hf2e6, 16'hf2e7 	:	val_out <= 16'h5779;
         16'hf2e8, 16'hf2e9, 16'hf2ea, 16'hf2eb, 16'hf2ec, 16'hf2ed, 16'hf2ee, 16'hf2ef 	:	val_out <= 16'h5791;
         16'hf2f0, 16'hf2f1, 16'hf2f2, 16'hf2f3, 16'hf2f4, 16'hf2f5, 16'hf2f6, 16'hf2f7 	:	val_out <= 16'h57a9;
         16'hf2f8, 16'hf2f9, 16'hf2fa, 16'hf2fb, 16'hf2fc, 16'hf2fd, 16'hf2fe, 16'hf2ff 	:	val_out <= 16'h57c1;
         16'hf300, 16'hf301, 16'hf302, 16'hf303, 16'hf304, 16'hf305, 16'hf306, 16'hf307 	:	val_out <= 16'h57d9;
         16'hf308, 16'hf309, 16'hf30a, 16'hf30b, 16'hf30c, 16'hf30d, 16'hf30e, 16'hf30f 	:	val_out <= 16'h57f1;
         16'hf310, 16'hf311, 16'hf312, 16'hf313, 16'hf314, 16'hf315, 16'hf316, 16'hf317 	:	val_out <= 16'h5809;
         16'hf318, 16'hf319, 16'hf31a, 16'hf31b, 16'hf31c, 16'hf31d, 16'hf31e, 16'hf31f 	:	val_out <= 16'h5820;
         16'hf320, 16'hf321, 16'hf322, 16'hf323, 16'hf324, 16'hf325, 16'hf326, 16'hf327 	:	val_out <= 16'h5838;
         16'hf328, 16'hf329, 16'hf32a, 16'hf32b, 16'hf32c, 16'hf32d, 16'hf32e, 16'hf32f 	:	val_out <= 16'h5850;
         16'hf330, 16'hf331, 16'hf332, 16'hf333, 16'hf334, 16'hf335, 16'hf336, 16'hf337 	:	val_out <= 16'h5868;
         16'hf338, 16'hf339, 16'hf33a, 16'hf33b, 16'hf33c, 16'hf33d, 16'hf33e, 16'hf33f 	:	val_out <= 16'h5880;
         16'hf340, 16'hf341, 16'hf342, 16'hf343, 16'hf344, 16'hf345, 16'hf346, 16'hf347 	:	val_out <= 16'h5898;
         16'hf348, 16'hf349, 16'hf34a, 16'hf34b, 16'hf34c, 16'hf34d, 16'hf34e, 16'hf34f 	:	val_out <= 16'h58b0;
         16'hf350, 16'hf351, 16'hf352, 16'hf353, 16'hf354, 16'hf355, 16'hf356, 16'hf357 	:	val_out <= 16'h58c8;
         16'hf358, 16'hf359, 16'hf35a, 16'hf35b, 16'hf35c, 16'hf35d, 16'hf35e, 16'hf35f 	:	val_out <= 16'h58e0;
         16'hf360, 16'hf361, 16'hf362, 16'hf363, 16'hf364, 16'hf365, 16'hf366, 16'hf367 	:	val_out <= 16'h58f8;
         16'hf368, 16'hf369, 16'hf36a, 16'hf36b, 16'hf36c, 16'hf36d, 16'hf36e, 16'hf36f 	:	val_out <= 16'h5910;
         16'hf370, 16'hf371, 16'hf372, 16'hf373, 16'hf374, 16'hf375, 16'hf376, 16'hf377 	:	val_out <= 16'h5927;
         16'hf378, 16'hf379, 16'hf37a, 16'hf37b, 16'hf37c, 16'hf37d, 16'hf37e, 16'hf37f 	:	val_out <= 16'h593f;
         16'hf380, 16'hf381, 16'hf382, 16'hf383, 16'hf384, 16'hf385, 16'hf386, 16'hf387 	:	val_out <= 16'h5957;
         16'hf388, 16'hf389, 16'hf38a, 16'hf38b, 16'hf38c, 16'hf38d, 16'hf38e, 16'hf38f 	:	val_out <= 16'h596f;
         16'hf390, 16'hf391, 16'hf392, 16'hf393, 16'hf394, 16'hf395, 16'hf396, 16'hf397 	:	val_out <= 16'h5987;
         16'hf398, 16'hf399, 16'hf39a, 16'hf39b, 16'hf39c, 16'hf39d, 16'hf39e, 16'hf39f 	:	val_out <= 16'h599f;
         16'hf3a0, 16'hf3a1, 16'hf3a2, 16'hf3a3, 16'hf3a4, 16'hf3a5, 16'hf3a6, 16'hf3a7 	:	val_out <= 16'h59b7;
         16'hf3a8, 16'hf3a9, 16'hf3aa, 16'hf3ab, 16'hf3ac, 16'hf3ad, 16'hf3ae, 16'hf3af 	:	val_out <= 16'h59cf;
         16'hf3b0, 16'hf3b1, 16'hf3b2, 16'hf3b3, 16'hf3b4, 16'hf3b5, 16'hf3b6, 16'hf3b7 	:	val_out <= 16'h59e7;
         16'hf3b8, 16'hf3b9, 16'hf3ba, 16'hf3bb, 16'hf3bc, 16'hf3bd, 16'hf3be, 16'hf3bf 	:	val_out <= 16'h59ff;
         16'hf3c0, 16'hf3c1, 16'hf3c2, 16'hf3c3, 16'hf3c4, 16'hf3c5, 16'hf3c6, 16'hf3c7 	:	val_out <= 16'h5a17;
         16'hf3c8, 16'hf3c9, 16'hf3ca, 16'hf3cb, 16'hf3cc, 16'hf3cd, 16'hf3ce, 16'hf3cf 	:	val_out <= 16'h5a2f;
         16'hf3d0, 16'hf3d1, 16'hf3d2, 16'hf3d3, 16'hf3d4, 16'hf3d5, 16'hf3d6, 16'hf3d7 	:	val_out <= 16'h5a47;
         16'hf3d8, 16'hf3d9, 16'hf3da, 16'hf3db, 16'hf3dc, 16'hf3dd, 16'hf3de, 16'hf3df 	:	val_out <= 16'h5a5f;
         16'hf3e0, 16'hf3e1, 16'hf3e2, 16'hf3e3, 16'hf3e4, 16'hf3e5, 16'hf3e6, 16'hf3e7 	:	val_out <= 16'h5a77;
         16'hf3e8, 16'hf3e9, 16'hf3ea, 16'hf3eb, 16'hf3ec, 16'hf3ed, 16'hf3ee, 16'hf3ef 	:	val_out <= 16'h5a8f;
         16'hf3f0, 16'hf3f1, 16'hf3f2, 16'hf3f3, 16'hf3f4, 16'hf3f5, 16'hf3f6, 16'hf3f7 	:	val_out <= 16'h5aa7;
         16'hf3f8, 16'hf3f9, 16'hf3fa, 16'hf3fb, 16'hf3fc, 16'hf3fd, 16'hf3fe, 16'hf3ff 	:	val_out <= 16'h5abf;
         16'hf400, 16'hf401, 16'hf402, 16'hf403, 16'hf404, 16'hf405, 16'hf406, 16'hf407 	:	val_out <= 16'h5ad7;
         16'hf408, 16'hf409, 16'hf40a, 16'hf40b, 16'hf40c, 16'hf40d, 16'hf40e, 16'hf40f 	:	val_out <= 16'h5af0;
         16'hf410, 16'hf411, 16'hf412, 16'hf413, 16'hf414, 16'hf415, 16'hf416, 16'hf417 	:	val_out <= 16'h5b08;
         16'hf418, 16'hf419, 16'hf41a, 16'hf41b, 16'hf41c, 16'hf41d, 16'hf41e, 16'hf41f 	:	val_out <= 16'h5b20;
         16'hf420, 16'hf421, 16'hf422, 16'hf423, 16'hf424, 16'hf425, 16'hf426, 16'hf427 	:	val_out <= 16'h5b38;
         16'hf428, 16'hf429, 16'hf42a, 16'hf42b, 16'hf42c, 16'hf42d, 16'hf42e, 16'hf42f 	:	val_out <= 16'h5b50;
         16'hf430, 16'hf431, 16'hf432, 16'hf433, 16'hf434, 16'hf435, 16'hf436, 16'hf437 	:	val_out <= 16'h5b68;
         16'hf438, 16'hf439, 16'hf43a, 16'hf43b, 16'hf43c, 16'hf43d, 16'hf43e, 16'hf43f 	:	val_out <= 16'h5b80;
         16'hf440, 16'hf441, 16'hf442, 16'hf443, 16'hf444, 16'hf445, 16'hf446, 16'hf447 	:	val_out <= 16'h5b98;
         16'hf448, 16'hf449, 16'hf44a, 16'hf44b, 16'hf44c, 16'hf44d, 16'hf44e, 16'hf44f 	:	val_out <= 16'h5bb0;
         16'hf450, 16'hf451, 16'hf452, 16'hf453, 16'hf454, 16'hf455, 16'hf456, 16'hf457 	:	val_out <= 16'h5bc8;
         16'hf458, 16'hf459, 16'hf45a, 16'hf45b, 16'hf45c, 16'hf45d, 16'hf45e, 16'hf45f 	:	val_out <= 16'h5be0;
         16'hf460, 16'hf461, 16'hf462, 16'hf463, 16'hf464, 16'hf465, 16'hf466, 16'hf467 	:	val_out <= 16'h5bf8;
         16'hf468, 16'hf469, 16'hf46a, 16'hf46b, 16'hf46c, 16'hf46d, 16'hf46e, 16'hf46f 	:	val_out <= 16'h5c11;
         16'hf470, 16'hf471, 16'hf472, 16'hf473, 16'hf474, 16'hf475, 16'hf476, 16'hf477 	:	val_out <= 16'h5c29;
         16'hf478, 16'hf479, 16'hf47a, 16'hf47b, 16'hf47c, 16'hf47d, 16'hf47e, 16'hf47f 	:	val_out <= 16'h5c41;
         16'hf480, 16'hf481, 16'hf482, 16'hf483, 16'hf484, 16'hf485, 16'hf486, 16'hf487 	:	val_out <= 16'h5c59;
         16'hf488, 16'hf489, 16'hf48a, 16'hf48b, 16'hf48c, 16'hf48d, 16'hf48e, 16'hf48f 	:	val_out <= 16'h5c71;
         16'hf490, 16'hf491, 16'hf492, 16'hf493, 16'hf494, 16'hf495, 16'hf496, 16'hf497 	:	val_out <= 16'h5c89;
         16'hf498, 16'hf499, 16'hf49a, 16'hf49b, 16'hf49c, 16'hf49d, 16'hf49e, 16'hf49f 	:	val_out <= 16'h5ca1;
         16'hf4a0, 16'hf4a1, 16'hf4a2, 16'hf4a3, 16'hf4a4, 16'hf4a5, 16'hf4a6, 16'hf4a7 	:	val_out <= 16'h5cba;
         16'hf4a8, 16'hf4a9, 16'hf4aa, 16'hf4ab, 16'hf4ac, 16'hf4ad, 16'hf4ae, 16'hf4af 	:	val_out <= 16'h5cd2;
         16'hf4b0, 16'hf4b1, 16'hf4b2, 16'hf4b3, 16'hf4b4, 16'hf4b5, 16'hf4b6, 16'hf4b7 	:	val_out <= 16'h5cea;
         16'hf4b8, 16'hf4b9, 16'hf4ba, 16'hf4bb, 16'hf4bc, 16'hf4bd, 16'hf4be, 16'hf4bf 	:	val_out <= 16'h5d02;
         16'hf4c0, 16'hf4c1, 16'hf4c2, 16'hf4c3, 16'hf4c4, 16'hf4c5, 16'hf4c6, 16'hf4c7 	:	val_out <= 16'h5d1a;
         16'hf4c8, 16'hf4c9, 16'hf4ca, 16'hf4cb, 16'hf4cc, 16'hf4cd, 16'hf4ce, 16'hf4cf 	:	val_out <= 16'h5d32;
         16'hf4d0, 16'hf4d1, 16'hf4d2, 16'hf4d3, 16'hf4d4, 16'hf4d5, 16'hf4d6, 16'hf4d7 	:	val_out <= 16'h5d4b;
         16'hf4d8, 16'hf4d9, 16'hf4da, 16'hf4db, 16'hf4dc, 16'hf4dd, 16'hf4de, 16'hf4df 	:	val_out <= 16'h5d63;
         16'hf4e0, 16'hf4e1, 16'hf4e2, 16'hf4e3, 16'hf4e4, 16'hf4e5, 16'hf4e6, 16'hf4e7 	:	val_out <= 16'h5d7b;
         16'hf4e8, 16'hf4e9, 16'hf4ea, 16'hf4eb, 16'hf4ec, 16'hf4ed, 16'hf4ee, 16'hf4ef 	:	val_out <= 16'h5d93;
         16'hf4f0, 16'hf4f1, 16'hf4f2, 16'hf4f3, 16'hf4f4, 16'hf4f5, 16'hf4f6, 16'hf4f7 	:	val_out <= 16'h5dab;
         16'hf4f8, 16'hf4f9, 16'hf4fa, 16'hf4fb, 16'hf4fc, 16'hf4fd, 16'hf4fe, 16'hf4ff 	:	val_out <= 16'h5dc4;
         16'hf500, 16'hf501, 16'hf502, 16'hf503, 16'hf504, 16'hf505, 16'hf506, 16'hf507 	:	val_out <= 16'h5ddc;
         16'hf508, 16'hf509, 16'hf50a, 16'hf50b, 16'hf50c, 16'hf50d, 16'hf50e, 16'hf50f 	:	val_out <= 16'h5df4;
         16'hf510, 16'hf511, 16'hf512, 16'hf513, 16'hf514, 16'hf515, 16'hf516, 16'hf517 	:	val_out <= 16'h5e0c;
         16'hf518, 16'hf519, 16'hf51a, 16'hf51b, 16'hf51c, 16'hf51d, 16'hf51e, 16'hf51f 	:	val_out <= 16'h5e25;
         16'hf520, 16'hf521, 16'hf522, 16'hf523, 16'hf524, 16'hf525, 16'hf526, 16'hf527 	:	val_out <= 16'h5e3d;
         16'hf528, 16'hf529, 16'hf52a, 16'hf52b, 16'hf52c, 16'hf52d, 16'hf52e, 16'hf52f 	:	val_out <= 16'h5e55;
         16'hf530, 16'hf531, 16'hf532, 16'hf533, 16'hf534, 16'hf535, 16'hf536, 16'hf537 	:	val_out <= 16'h5e6d;
         16'hf538, 16'hf539, 16'hf53a, 16'hf53b, 16'hf53c, 16'hf53d, 16'hf53e, 16'hf53f 	:	val_out <= 16'h5e86;
         16'hf540, 16'hf541, 16'hf542, 16'hf543, 16'hf544, 16'hf545, 16'hf546, 16'hf547 	:	val_out <= 16'h5e9e;
         16'hf548, 16'hf549, 16'hf54a, 16'hf54b, 16'hf54c, 16'hf54d, 16'hf54e, 16'hf54f 	:	val_out <= 16'h5eb6;
         16'hf550, 16'hf551, 16'hf552, 16'hf553, 16'hf554, 16'hf555, 16'hf556, 16'hf557 	:	val_out <= 16'h5ece;
         16'hf558, 16'hf559, 16'hf55a, 16'hf55b, 16'hf55c, 16'hf55d, 16'hf55e, 16'hf55f 	:	val_out <= 16'h5ee7;
         16'hf560, 16'hf561, 16'hf562, 16'hf563, 16'hf564, 16'hf565, 16'hf566, 16'hf567 	:	val_out <= 16'h5eff;
         16'hf568, 16'hf569, 16'hf56a, 16'hf56b, 16'hf56c, 16'hf56d, 16'hf56e, 16'hf56f 	:	val_out <= 16'h5f17;
         16'hf570, 16'hf571, 16'hf572, 16'hf573, 16'hf574, 16'hf575, 16'hf576, 16'hf577 	:	val_out <= 16'h5f2f;
         16'hf578, 16'hf579, 16'hf57a, 16'hf57b, 16'hf57c, 16'hf57d, 16'hf57e, 16'hf57f 	:	val_out <= 16'h5f48;
         16'hf580, 16'hf581, 16'hf582, 16'hf583, 16'hf584, 16'hf585, 16'hf586, 16'hf587 	:	val_out <= 16'h5f60;
         16'hf588, 16'hf589, 16'hf58a, 16'hf58b, 16'hf58c, 16'hf58d, 16'hf58e, 16'hf58f 	:	val_out <= 16'h5f78;
         16'hf590, 16'hf591, 16'hf592, 16'hf593, 16'hf594, 16'hf595, 16'hf596, 16'hf597 	:	val_out <= 16'h5f91;
         16'hf598, 16'hf599, 16'hf59a, 16'hf59b, 16'hf59c, 16'hf59d, 16'hf59e, 16'hf59f 	:	val_out <= 16'h5fa9;
         16'hf5a0, 16'hf5a1, 16'hf5a2, 16'hf5a3, 16'hf5a4, 16'hf5a5, 16'hf5a6, 16'hf5a7 	:	val_out <= 16'h5fc1;
         16'hf5a8, 16'hf5a9, 16'hf5aa, 16'hf5ab, 16'hf5ac, 16'hf5ad, 16'hf5ae, 16'hf5af 	:	val_out <= 16'h5fda;
         16'hf5b0, 16'hf5b1, 16'hf5b2, 16'hf5b3, 16'hf5b4, 16'hf5b5, 16'hf5b6, 16'hf5b7 	:	val_out <= 16'h5ff2;
         16'hf5b8, 16'hf5b9, 16'hf5ba, 16'hf5bb, 16'hf5bc, 16'hf5bd, 16'hf5be, 16'hf5bf 	:	val_out <= 16'h600a;
         16'hf5c0, 16'hf5c1, 16'hf5c2, 16'hf5c3, 16'hf5c4, 16'hf5c5, 16'hf5c6, 16'hf5c7 	:	val_out <= 16'h6023;
         16'hf5c8, 16'hf5c9, 16'hf5ca, 16'hf5cb, 16'hf5cc, 16'hf5cd, 16'hf5ce, 16'hf5cf 	:	val_out <= 16'h603b;
         16'hf5d0, 16'hf5d1, 16'hf5d2, 16'hf5d3, 16'hf5d4, 16'hf5d5, 16'hf5d6, 16'hf5d7 	:	val_out <= 16'h6053;
         16'hf5d8, 16'hf5d9, 16'hf5da, 16'hf5db, 16'hf5dc, 16'hf5dd, 16'hf5de, 16'hf5df 	:	val_out <= 16'h606c;
         16'hf5e0, 16'hf5e1, 16'hf5e2, 16'hf5e3, 16'hf5e4, 16'hf5e5, 16'hf5e6, 16'hf5e7 	:	val_out <= 16'h6084;
         16'hf5e8, 16'hf5e9, 16'hf5ea, 16'hf5eb, 16'hf5ec, 16'hf5ed, 16'hf5ee, 16'hf5ef 	:	val_out <= 16'h609c;
         16'hf5f0, 16'hf5f1, 16'hf5f2, 16'hf5f3, 16'hf5f4, 16'hf5f5, 16'hf5f6, 16'hf5f7 	:	val_out <= 16'h60b5;
         16'hf5f8, 16'hf5f9, 16'hf5fa, 16'hf5fb, 16'hf5fc, 16'hf5fd, 16'hf5fe, 16'hf5ff 	:	val_out <= 16'h60cd;
         16'hf600, 16'hf601, 16'hf602, 16'hf603, 16'hf604, 16'hf605, 16'hf606, 16'hf607 	:	val_out <= 16'h60e6;
         16'hf608, 16'hf609, 16'hf60a, 16'hf60b, 16'hf60c, 16'hf60d, 16'hf60e, 16'hf60f 	:	val_out <= 16'h60fe;
         16'hf610, 16'hf611, 16'hf612, 16'hf613, 16'hf614, 16'hf615, 16'hf616, 16'hf617 	:	val_out <= 16'h6116;
         16'hf618, 16'hf619, 16'hf61a, 16'hf61b, 16'hf61c, 16'hf61d, 16'hf61e, 16'hf61f 	:	val_out <= 16'h612f;
         16'hf620, 16'hf621, 16'hf622, 16'hf623, 16'hf624, 16'hf625, 16'hf626, 16'hf627 	:	val_out <= 16'h6147;
         16'hf628, 16'hf629, 16'hf62a, 16'hf62b, 16'hf62c, 16'hf62d, 16'hf62e, 16'hf62f 	:	val_out <= 16'h615f;
         16'hf630, 16'hf631, 16'hf632, 16'hf633, 16'hf634, 16'hf635, 16'hf636, 16'hf637 	:	val_out <= 16'h6178;
         16'hf638, 16'hf639, 16'hf63a, 16'hf63b, 16'hf63c, 16'hf63d, 16'hf63e, 16'hf63f 	:	val_out <= 16'h6190;
         16'hf640, 16'hf641, 16'hf642, 16'hf643, 16'hf644, 16'hf645, 16'hf646, 16'hf647 	:	val_out <= 16'h61a9;
         16'hf648, 16'hf649, 16'hf64a, 16'hf64b, 16'hf64c, 16'hf64d, 16'hf64e, 16'hf64f 	:	val_out <= 16'h61c1;
         16'hf650, 16'hf651, 16'hf652, 16'hf653, 16'hf654, 16'hf655, 16'hf656, 16'hf657 	:	val_out <= 16'h61da;
         16'hf658, 16'hf659, 16'hf65a, 16'hf65b, 16'hf65c, 16'hf65d, 16'hf65e, 16'hf65f 	:	val_out <= 16'h61f2;
         16'hf660, 16'hf661, 16'hf662, 16'hf663, 16'hf664, 16'hf665, 16'hf666, 16'hf667 	:	val_out <= 16'h620a;
         16'hf668, 16'hf669, 16'hf66a, 16'hf66b, 16'hf66c, 16'hf66d, 16'hf66e, 16'hf66f 	:	val_out <= 16'h6223;
         16'hf670, 16'hf671, 16'hf672, 16'hf673, 16'hf674, 16'hf675, 16'hf676, 16'hf677 	:	val_out <= 16'h623b;
         16'hf678, 16'hf679, 16'hf67a, 16'hf67b, 16'hf67c, 16'hf67d, 16'hf67e, 16'hf67f 	:	val_out <= 16'h6254;
         16'hf680, 16'hf681, 16'hf682, 16'hf683, 16'hf684, 16'hf685, 16'hf686, 16'hf687 	:	val_out <= 16'h626c;
         16'hf688, 16'hf689, 16'hf68a, 16'hf68b, 16'hf68c, 16'hf68d, 16'hf68e, 16'hf68f 	:	val_out <= 16'h6285;
         16'hf690, 16'hf691, 16'hf692, 16'hf693, 16'hf694, 16'hf695, 16'hf696, 16'hf697 	:	val_out <= 16'h629d;
         16'hf698, 16'hf699, 16'hf69a, 16'hf69b, 16'hf69c, 16'hf69d, 16'hf69e, 16'hf69f 	:	val_out <= 16'h62b6;
         16'hf6a0, 16'hf6a1, 16'hf6a2, 16'hf6a3, 16'hf6a4, 16'hf6a5, 16'hf6a6, 16'hf6a7 	:	val_out <= 16'h62ce;
         16'hf6a8, 16'hf6a9, 16'hf6aa, 16'hf6ab, 16'hf6ac, 16'hf6ad, 16'hf6ae, 16'hf6af 	:	val_out <= 16'h62e7;
         16'hf6b0, 16'hf6b1, 16'hf6b2, 16'hf6b3, 16'hf6b4, 16'hf6b5, 16'hf6b6, 16'hf6b7 	:	val_out <= 16'h62ff;
         16'hf6b8, 16'hf6b9, 16'hf6ba, 16'hf6bb, 16'hf6bc, 16'hf6bd, 16'hf6be, 16'hf6bf 	:	val_out <= 16'h6317;
         16'hf6c0, 16'hf6c1, 16'hf6c2, 16'hf6c3, 16'hf6c4, 16'hf6c5, 16'hf6c6, 16'hf6c7 	:	val_out <= 16'h6330;
         16'hf6c8, 16'hf6c9, 16'hf6ca, 16'hf6cb, 16'hf6cc, 16'hf6cd, 16'hf6ce, 16'hf6cf 	:	val_out <= 16'h6348;
         16'hf6d0, 16'hf6d1, 16'hf6d2, 16'hf6d3, 16'hf6d4, 16'hf6d5, 16'hf6d6, 16'hf6d7 	:	val_out <= 16'h6361;
         16'hf6d8, 16'hf6d9, 16'hf6da, 16'hf6db, 16'hf6dc, 16'hf6dd, 16'hf6de, 16'hf6df 	:	val_out <= 16'h6379;
         16'hf6e0, 16'hf6e1, 16'hf6e2, 16'hf6e3, 16'hf6e4, 16'hf6e5, 16'hf6e6, 16'hf6e7 	:	val_out <= 16'h6392;
         16'hf6e8, 16'hf6e9, 16'hf6ea, 16'hf6eb, 16'hf6ec, 16'hf6ed, 16'hf6ee, 16'hf6ef 	:	val_out <= 16'h63aa;
         16'hf6f0, 16'hf6f1, 16'hf6f2, 16'hf6f3, 16'hf6f4, 16'hf6f5, 16'hf6f6, 16'hf6f7 	:	val_out <= 16'h63c3;
         16'hf6f8, 16'hf6f9, 16'hf6fa, 16'hf6fb, 16'hf6fc, 16'hf6fd, 16'hf6fe, 16'hf6ff 	:	val_out <= 16'h63db;
         16'hf700, 16'hf701, 16'hf702, 16'hf703, 16'hf704, 16'hf705, 16'hf706, 16'hf707 	:	val_out <= 16'h63f4;
         16'hf708, 16'hf709, 16'hf70a, 16'hf70b, 16'hf70c, 16'hf70d, 16'hf70e, 16'hf70f 	:	val_out <= 16'h640d;
         16'hf710, 16'hf711, 16'hf712, 16'hf713, 16'hf714, 16'hf715, 16'hf716, 16'hf717 	:	val_out <= 16'h6425;
         16'hf718, 16'hf719, 16'hf71a, 16'hf71b, 16'hf71c, 16'hf71d, 16'hf71e, 16'hf71f 	:	val_out <= 16'h643e;
         16'hf720, 16'hf721, 16'hf722, 16'hf723, 16'hf724, 16'hf725, 16'hf726, 16'hf727 	:	val_out <= 16'h6456;
         16'hf728, 16'hf729, 16'hf72a, 16'hf72b, 16'hf72c, 16'hf72d, 16'hf72e, 16'hf72f 	:	val_out <= 16'h646f;
         16'hf730, 16'hf731, 16'hf732, 16'hf733, 16'hf734, 16'hf735, 16'hf736, 16'hf737 	:	val_out <= 16'h6487;
         16'hf738, 16'hf739, 16'hf73a, 16'hf73b, 16'hf73c, 16'hf73d, 16'hf73e, 16'hf73f 	:	val_out <= 16'h64a0;
         16'hf740, 16'hf741, 16'hf742, 16'hf743, 16'hf744, 16'hf745, 16'hf746, 16'hf747 	:	val_out <= 16'h64b8;
         16'hf748, 16'hf749, 16'hf74a, 16'hf74b, 16'hf74c, 16'hf74d, 16'hf74e, 16'hf74f 	:	val_out <= 16'h64d1;
         16'hf750, 16'hf751, 16'hf752, 16'hf753, 16'hf754, 16'hf755, 16'hf756, 16'hf757 	:	val_out <= 16'h64e9;
         16'hf758, 16'hf759, 16'hf75a, 16'hf75b, 16'hf75c, 16'hf75d, 16'hf75e, 16'hf75f 	:	val_out <= 16'h6502;
         16'hf760, 16'hf761, 16'hf762, 16'hf763, 16'hf764, 16'hf765, 16'hf766, 16'hf767 	:	val_out <= 16'h651b;
         16'hf768, 16'hf769, 16'hf76a, 16'hf76b, 16'hf76c, 16'hf76d, 16'hf76e, 16'hf76f 	:	val_out <= 16'h6533;
         16'hf770, 16'hf771, 16'hf772, 16'hf773, 16'hf774, 16'hf775, 16'hf776, 16'hf777 	:	val_out <= 16'h654c;
         16'hf778, 16'hf779, 16'hf77a, 16'hf77b, 16'hf77c, 16'hf77d, 16'hf77e, 16'hf77f 	:	val_out <= 16'h6564;
         16'hf780, 16'hf781, 16'hf782, 16'hf783, 16'hf784, 16'hf785, 16'hf786, 16'hf787 	:	val_out <= 16'h657d;
         16'hf788, 16'hf789, 16'hf78a, 16'hf78b, 16'hf78c, 16'hf78d, 16'hf78e, 16'hf78f 	:	val_out <= 16'h6595;
         16'hf790, 16'hf791, 16'hf792, 16'hf793, 16'hf794, 16'hf795, 16'hf796, 16'hf797 	:	val_out <= 16'h65ae;
         16'hf798, 16'hf799, 16'hf79a, 16'hf79b, 16'hf79c, 16'hf79d, 16'hf79e, 16'hf79f 	:	val_out <= 16'h65c7;
         16'hf7a0, 16'hf7a1, 16'hf7a2, 16'hf7a3, 16'hf7a4, 16'hf7a5, 16'hf7a6, 16'hf7a7 	:	val_out <= 16'h65df;
         16'hf7a8, 16'hf7a9, 16'hf7aa, 16'hf7ab, 16'hf7ac, 16'hf7ad, 16'hf7ae, 16'hf7af 	:	val_out <= 16'h65f8;
         16'hf7b0, 16'hf7b1, 16'hf7b2, 16'hf7b3, 16'hf7b4, 16'hf7b5, 16'hf7b6, 16'hf7b7 	:	val_out <= 16'h6610;
         16'hf7b8, 16'hf7b9, 16'hf7ba, 16'hf7bb, 16'hf7bc, 16'hf7bd, 16'hf7be, 16'hf7bf 	:	val_out <= 16'h6629;
         16'hf7c0, 16'hf7c1, 16'hf7c2, 16'hf7c3, 16'hf7c4, 16'hf7c5, 16'hf7c6, 16'hf7c7 	:	val_out <= 16'h6642;
         16'hf7c8, 16'hf7c9, 16'hf7ca, 16'hf7cb, 16'hf7cc, 16'hf7cd, 16'hf7ce, 16'hf7cf 	:	val_out <= 16'h665a;
         16'hf7d0, 16'hf7d1, 16'hf7d2, 16'hf7d3, 16'hf7d4, 16'hf7d5, 16'hf7d6, 16'hf7d7 	:	val_out <= 16'h6673;
         16'hf7d8, 16'hf7d9, 16'hf7da, 16'hf7db, 16'hf7dc, 16'hf7dd, 16'hf7de, 16'hf7df 	:	val_out <= 16'h668c;
         16'hf7e0, 16'hf7e1, 16'hf7e2, 16'hf7e3, 16'hf7e4, 16'hf7e5, 16'hf7e6, 16'hf7e7 	:	val_out <= 16'h66a4;
         16'hf7e8, 16'hf7e9, 16'hf7ea, 16'hf7eb, 16'hf7ec, 16'hf7ed, 16'hf7ee, 16'hf7ef 	:	val_out <= 16'h66bd;
         16'hf7f0, 16'hf7f1, 16'hf7f2, 16'hf7f3, 16'hf7f4, 16'hf7f5, 16'hf7f6, 16'hf7f7 	:	val_out <= 16'h66d5;
         16'hf7f8, 16'hf7f9, 16'hf7fa, 16'hf7fb, 16'hf7fc, 16'hf7fd, 16'hf7fe, 16'hf7ff 	:	val_out <= 16'h66ee;
         16'hf800, 16'hf801, 16'hf802, 16'hf803, 16'hf804, 16'hf805, 16'hf806, 16'hf807 	:	val_out <= 16'h6707;
         16'hf808, 16'hf809, 16'hf80a, 16'hf80b, 16'hf80c, 16'hf80d, 16'hf80e, 16'hf80f 	:	val_out <= 16'h671f;
         16'hf810, 16'hf811, 16'hf812, 16'hf813, 16'hf814, 16'hf815, 16'hf816, 16'hf817 	:	val_out <= 16'h6738;
         16'hf818, 16'hf819, 16'hf81a, 16'hf81b, 16'hf81c, 16'hf81d, 16'hf81e, 16'hf81f 	:	val_out <= 16'h6751;
         16'hf820, 16'hf821, 16'hf822, 16'hf823, 16'hf824, 16'hf825, 16'hf826, 16'hf827 	:	val_out <= 16'h6769;
         16'hf828, 16'hf829, 16'hf82a, 16'hf82b, 16'hf82c, 16'hf82d, 16'hf82e, 16'hf82f 	:	val_out <= 16'h6782;
         16'hf830, 16'hf831, 16'hf832, 16'hf833, 16'hf834, 16'hf835, 16'hf836, 16'hf837 	:	val_out <= 16'h679b;
         16'hf838, 16'hf839, 16'hf83a, 16'hf83b, 16'hf83c, 16'hf83d, 16'hf83e, 16'hf83f 	:	val_out <= 16'h67b3;
         16'hf840, 16'hf841, 16'hf842, 16'hf843, 16'hf844, 16'hf845, 16'hf846, 16'hf847 	:	val_out <= 16'h67cc;
         16'hf848, 16'hf849, 16'hf84a, 16'hf84b, 16'hf84c, 16'hf84d, 16'hf84e, 16'hf84f 	:	val_out <= 16'h67e5;
         16'hf850, 16'hf851, 16'hf852, 16'hf853, 16'hf854, 16'hf855, 16'hf856, 16'hf857 	:	val_out <= 16'h67fd;
         16'hf858, 16'hf859, 16'hf85a, 16'hf85b, 16'hf85c, 16'hf85d, 16'hf85e, 16'hf85f 	:	val_out <= 16'h6816;
         16'hf860, 16'hf861, 16'hf862, 16'hf863, 16'hf864, 16'hf865, 16'hf866, 16'hf867 	:	val_out <= 16'h682f;
         16'hf868, 16'hf869, 16'hf86a, 16'hf86b, 16'hf86c, 16'hf86d, 16'hf86e, 16'hf86f 	:	val_out <= 16'h6848;
         16'hf870, 16'hf871, 16'hf872, 16'hf873, 16'hf874, 16'hf875, 16'hf876, 16'hf877 	:	val_out <= 16'h6860;
         16'hf878, 16'hf879, 16'hf87a, 16'hf87b, 16'hf87c, 16'hf87d, 16'hf87e, 16'hf87f 	:	val_out <= 16'h6879;
         16'hf880, 16'hf881, 16'hf882, 16'hf883, 16'hf884, 16'hf885, 16'hf886, 16'hf887 	:	val_out <= 16'h6892;
         16'hf888, 16'hf889, 16'hf88a, 16'hf88b, 16'hf88c, 16'hf88d, 16'hf88e, 16'hf88f 	:	val_out <= 16'h68aa;
         16'hf890, 16'hf891, 16'hf892, 16'hf893, 16'hf894, 16'hf895, 16'hf896, 16'hf897 	:	val_out <= 16'h68c3;
         16'hf898, 16'hf899, 16'hf89a, 16'hf89b, 16'hf89c, 16'hf89d, 16'hf89e, 16'hf89f 	:	val_out <= 16'h68dc;
         16'hf8a0, 16'hf8a1, 16'hf8a2, 16'hf8a3, 16'hf8a4, 16'hf8a5, 16'hf8a6, 16'hf8a7 	:	val_out <= 16'h68f5;
         16'hf8a8, 16'hf8a9, 16'hf8aa, 16'hf8ab, 16'hf8ac, 16'hf8ad, 16'hf8ae, 16'hf8af 	:	val_out <= 16'h690d;
         16'hf8b0, 16'hf8b1, 16'hf8b2, 16'hf8b3, 16'hf8b4, 16'hf8b5, 16'hf8b6, 16'hf8b7 	:	val_out <= 16'h6926;
         16'hf8b8, 16'hf8b9, 16'hf8ba, 16'hf8bb, 16'hf8bc, 16'hf8bd, 16'hf8be, 16'hf8bf 	:	val_out <= 16'h693f;
         16'hf8c0, 16'hf8c1, 16'hf8c2, 16'hf8c3, 16'hf8c4, 16'hf8c5, 16'hf8c6, 16'hf8c7 	:	val_out <= 16'h6957;
         16'hf8c8, 16'hf8c9, 16'hf8ca, 16'hf8cb, 16'hf8cc, 16'hf8cd, 16'hf8ce, 16'hf8cf 	:	val_out <= 16'h6970;
         16'hf8d0, 16'hf8d1, 16'hf8d2, 16'hf8d3, 16'hf8d4, 16'hf8d5, 16'hf8d6, 16'hf8d7 	:	val_out <= 16'h6989;
         16'hf8d8, 16'hf8d9, 16'hf8da, 16'hf8db, 16'hf8dc, 16'hf8dd, 16'hf8de, 16'hf8df 	:	val_out <= 16'h69a2;
         16'hf8e0, 16'hf8e1, 16'hf8e2, 16'hf8e3, 16'hf8e4, 16'hf8e5, 16'hf8e6, 16'hf8e7 	:	val_out <= 16'h69ba;
         16'hf8e8, 16'hf8e9, 16'hf8ea, 16'hf8eb, 16'hf8ec, 16'hf8ed, 16'hf8ee, 16'hf8ef 	:	val_out <= 16'h69d3;
         16'hf8f0, 16'hf8f1, 16'hf8f2, 16'hf8f3, 16'hf8f4, 16'hf8f5, 16'hf8f6, 16'hf8f7 	:	val_out <= 16'h69ec;
         16'hf8f8, 16'hf8f9, 16'hf8fa, 16'hf8fb, 16'hf8fc, 16'hf8fd, 16'hf8fe, 16'hf8ff 	:	val_out <= 16'h6a05;
         16'hf900, 16'hf901, 16'hf902, 16'hf903, 16'hf904, 16'hf905, 16'hf906, 16'hf907 	:	val_out <= 16'h6a1d;
         16'hf908, 16'hf909, 16'hf90a, 16'hf90b, 16'hf90c, 16'hf90d, 16'hf90e, 16'hf90f 	:	val_out <= 16'h6a36;
         16'hf910, 16'hf911, 16'hf912, 16'hf913, 16'hf914, 16'hf915, 16'hf916, 16'hf917 	:	val_out <= 16'h6a4f;
         16'hf918, 16'hf919, 16'hf91a, 16'hf91b, 16'hf91c, 16'hf91d, 16'hf91e, 16'hf91f 	:	val_out <= 16'h6a68;
         16'hf920, 16'hf921, 16'hf922, 16'hf923, 16'hf924, 16'hf925, 16'hf926, 16'hf927 	:	val_out <= 16'h6a80;
         16'hf928, 16'hf929, 16'hf92a, 16'hf92b, 16'hf92c, 16'hf92d, 16'hf92e, 16'hf92f 	:	val_out <= 16'h6a99;
         16'hf930, 16'hf931, 16'hf932, 16'hf933, 16'hf934, 16'hf935, 16'hf936, 16'hf937 	:	val_out <= 16'h6ab2;
         16'hf938, 16'hf939, 16'hf93a, 16'hf93b, 16'hf93c, 16'hf93d, 16'hf93e, 16'hf93f 	:	val_out <= 16'h6acb;
         16'hf940, 16'hf941, 16'hf942, 16'hf943, 16'hf944, 16'hf945, 16'hf946, 16'hf947 	:	val_out <= 16'h6ae4;
         16'hf948, 16'hf949, 16'hf94a, 16'hf94b, 16'hf94c, 16'hf94d, 16'hf94e, 16'hf94f 	:	val_out <= 16'h6afc;
         16'hf950, 16'hf951, 16'hf952, 16'hf953, 16'hf954, 16'hf955, 16'hf956, 16'hf957 	:	val_out <= 16'h6b15;
         16'hf958, 16'hf959, 16'hf95a, 16'hf95b, 16'hf95c, 16'hf95d, 16'hf95e, 16'hf95f 	:	val_out <= 16'h6b2e;
         16'hf960, 16'hf961, 16'hf962, 16'hf963, 16'hf964, 16'hf965, 16'hf966, 16'hf967 	:	val_out <= 16'h6b47;
         16'hf968, 16'hf969, 16'hf96a, 16'hf96b, 16'hf96c, 16'hf96d, 16'hf96e, 16'hf96f 	:	val_out <= 16'h6b60;
         16'hf970, 16'hf971, 16'hf972, 16'hf973, 16'hf974, 16'hf975, 16'hf976, 16'hf977 	:	val_out <= 16'h6b78;
         16'hf978, 16'hf979, 16'hf97a, 16'hf97b, 16'hf97c, 16'hf97d, 16'hf97e, 16'hf97f 	:	val_out <= 16'h6b91;
         16'hf980, 16'hf981, 16'hf982, 16'hf983, 16'hf984, 16'hf985, 16'hf986, 16'hf987 	:	val_out <= 16'h6baa;
         16'hf988, 16'hf989, 16'hf98a, 16'hf98b, 16'hf98c, 16'hf98d, 16'hf98e, 16'hf98f 	:	val_out <= 16'h6bc3;
         16'hf990, 16'hf991, 16'hf992, 16'hf993, 16'hf994, 16'hf995, 16'hf996, 16'hf997 	:	val_out <= 16'h6bdc;
         16'hf998, 16'hf999, 16'hf99a, 16'hf99b, 16'hf99c, 16'hf99d, 16'hf99e, 16'hf99f 	:	val_out <= 16'h6bf4;
         16'hf9a0, 16'hf9a1, 16'hf9a2, 16'hf9a3, 16'hf9a4, 16'hf9a5, 16'hf9a6, 16'hf9a7 	:	val_out <= 16'h6c0d;
         16'hf9a8, 16'hf9a9, 16'hf9aa, 16'hf9ab, 16'hf9ac, 16'hf9ad, 16'hf9ae, 16'hf9af 	:	val_out <= 16'h6c26;
         16'hf9b0, 16'hf9b1, 16'hf9b2, 16'hf9b3, 16'hf9b4, 16'hf9b5, 16'hf9b6, 16'hf9b7 	:	val_out <= 16'h6c3f;
         16'hf9b8, 16'hf9b9, 16'hf9ba, 16'hf9bb, 16'hf9bc, 16'hf9bd, 16'hf9be, 16'hf9bf 	:	val_out <= 16'h6c58;
         16'hf9c0, 16'hf9c1, 16'hf9c2, 16'hf9c3, 16'hf9c4, 16'hf9c5, 16'hf9c6, 16'hf9c7 	:	val_out <= 16'h6c71;
         16'hf9c8, 16'hf9c9, 16'hf9ca, 16'hf9cb, 16'hf9cc, 16'hf9cd, 16'hf9ce, 16'hf9cf 	:	val_out <= 16'h6c89;
         16'hf9d0, 16'hf9d1, 16'hf9d2, 16'hf9d3, 16'hf9d4, 16'hf9d5, 16'hf9d6, 16'hf9d7 	:	val_out <= 16'h6ca2;
         16'hf9d8, 16'hf9d9, 16'hf9da, 16'hf9db, 16'hf9dc, 16'hf9dd, 16'hf9de, 16'hf9df 	:	val_out <= 16'h6cbb;
         16'hf9e0, 16'hf9e1, 16'hf9e2, 16'hf9e3, 16'hf9e4, 16'hf9e5, 16'hf9e6, 16'hf9e7 	:	val_out <= 16'h6cd4;
         16'hf9e8, 16'hf9e9, 16'hf9ea, 16'hf9eb, 16'hf9ec, 16'hf9ed, 16'hf9ee, 16'hf9ef 	:	val_out <= 16'h6ced;
         16'hf9f0, 16'hf9f1, 16'hf9f2, 16'hf9f3, 16'hf9f4, 16'hf9f5, 16'hf9f6, 16'hf9f7 	:	val_out <= 16'h6d06;
         16'hf9f8, 16'hf9f9, 16'hf9fa, 16'hf9fb, 16'hf9fc, 16'hf9fd, 16'hf9fe, 16'hf9ff 	:	val_out <= 16'h6d1f;
         16'hfa00, 16'hfa01, 16'hfa02, 16'hfa03, 16'hfa04, 16'hfa05, 16'hfa06, 16'hfa07 	:	val_out <= 16'h6d37;
         16'hfa08, 16'hfa09, 16'hfa0a, 16'hfa0b, 16'hfa0c, 16'hfa0d, 16'hfa0e, 16'hfa0f 	:	val_out <= 16'h6d50;
         16'hfa10, 16'hfa11, 16'hfa12, 16'hfa13, 16'hfa14, 16'hfa15, 16'hfa16, 16'hfa17 	:	val_out <= 16'h6d69;
         16'hfa18, 16'hfa19, 16'hfa1a, 16'hfa1b, 16'hfa1c, 16'hfa1d, 16'hfa1e, 16'hfa1f 	:	val_out <= 16'h6d82;
         16'hfa20, 16'hfa21, 16'hfa22, 16'hfa23, 16'hfa24, 16'hfa25, 16'hfa26, 16'hfa27 	:	val_out <= 16'h6d9b;
         16'hfa28, 16'hfa29, 16'hfa2a, 16'hfa2b, 16'hfa2c, 16'hfa2d, 16'hfa2e, 16'hfa2f 	:	val_out <= 16'h6db4;
         16'hfa30, 16'hfa31, 16'hfa32, 16'hfa33, 16'hfa34, 16'hfa35, 16'hfa36, 16'hfa37 	:	val_out <= 16'h6dcd;
         16'hfa38, 16'hfa39, 16'hfa3a, 16'hfa3b, 16'hfa3c, 16'hfa3d, 16'hfa3e, 16'hfa3f 	:	val_out <= 16'h6de6;
         16'hfa40, 16'hfa41, 16'hfa42, 16'hfa43, 16'hfa44, 16'hfa45, 16'hfa46, 16'hfa47 	:	val_out <= 16'h6dfe;
         16'hfa48, 16'hfa49, 16'hfa4a, 16'hfa4b, 16'hfa4c, 16'hfa4d, 16'hfa4e, 16'hfa4f 	:	val_out <= 16'h6e17;
         16'hfa50, 16'hfa51, 16'hfa52, 16'hfa53, 16'hfa54, 16'hfa55, 16'hfa56, 16'hfa57 	:	val_out <= 16'h6e30;
         16'hfa58, 16'hfa59, 16'hfa5a, 16'hfa5b, 16'hfa5c, 16'hfa5d, 16'hfa5e, 16'hfa5f 	:	val_out <= 16'h6e49;
         16'hfa60, 16'hfa61, 16'hfa62, 16'hfa63, 16'hfa64, 16'hfa65, 16'hfa66, 16'hfa67 	:	val_out <= 16'h6e62;
         16'hfa68, 16'hfa69, 16'hfa6a, 16'hfa6b, 16'hfa6c, 16'hfa6d, 16'hfa6e, 16'hfa6f 	:	val_out <= 16'h6e7b;
         16'hfa70, 16'hfa71, 16'hfa72, 16'hfa73, 16'hfa74, 16'hfa75, 16'hfa76, 16'hfa77 	:	val_out <= 16'h6e94;
         16'hfa78, 16'hfa79, 16'hfa7a, 16'hfa7b, 16'hfa7c, 16'hfa7d, 16'hfa7e, 16'hfa7f 	:	val_out <= 16'h6ead;
         16'hfa80, 16'hfa81, 16'hfa82, 16'hfa83, 16'hfa84, 16'hfa85, 16'hfa86, 16'hfa87 	:	val_out <= 16'h6ec6;
         16'hfa88, 16'hfa89, 16'hfa8a, 16'hfa8b, 16'hfa8c, 16'hfa8d, 16'hfa8e, 16'hfa8f 	:	val_out <= 16'h6ede;
         16'hfa90, 16'hfa91, 16'hfa92, 16'hfa93, 16'hfa94, 16'hfa95, 16'hfa96, 16'hfa97 	:	val_out <= 16'h6ef7;
         16'hfa98, 16'hfa99, 16'hfa9a, 16'hfa9b, 16'hfa9c, 16'hfa9d, 16'hfa9e, 16'hfa9f 	:	val_out <= 16'h6f10;
         16'hfaa0, 16'hfaa1, 16'hfaa2, 16'hfaa3, 16'hfaa4, 16'hfaa5, 16'hfaa6, 16'hfaa7 	:	val_out <= 16'h6f29;
         16'hfaa8, 16'hfaa9, 16'hfaaa, 16'hfaab, 16'hfaac, 16'hfaad, 16'hfaae, 16'hfaaf 	:	val_out <= 16'h6f42;
         16'hfab0, 16'hfab1, 16'hfab2, 16'hfab3, 16'hfab4, 16'hfab5, 16'hfab6, 16'hfab7 	:	val_out <= 16'h6f5b;
         16'hfab8, 16'hfab9, 16'hfaba, 16'hfabb, 16'hfabc, 16'hfabd, 16'hfabe, 16'hfabf 	:	val_out <= 16'h6f74;
         16'hfac0, 16'hfac1, 16'hfac2, 16'hfac3, 16'hfac4, 16'hfac5, 16'hfac6, 16'hfac7 	:	val_out <= 16'h6f8d;
         16'hfac8, 16'hfac9, 16'hfaca, 16'hfacb, 16'hfacc, 16'hfacd, 16'hface, 16'hfacf 	:	val_out <= 16'h6fa6;
         16'hfad0, 16'hfad1, 16'hfad2, 16'hfad3, 16'hfad4, 16'hfad5, 16'hfad6, 16'hfad7 	:	val_out <= 16'h6fbf;
         16'hfad8, 16'hfad9, 16'hfada, 16'hfadb, 16'hfadc, 16'hfadd, 16'hfade, 16'hfadf 	:	val_out <= 16'h6fd8;
         16'hfae0, 16'hfae1, 16'hfae2, 16'hfae3, 16'hfae4, 16'hfae5, 16'hfae6, 16'hfae7 	:	val_out <= 16'h6ff1;
         16'hfae8, 16'hfae9, 16'hfaea, 16'hfaeb, 16'hfaec, 16'hfaed, 16'hfaee, 16'hfaef 	:	val_out <= 16'h700a;
         16'hfaf0, 16'hfaf1, 16'hfaf2, 16'hfaf3, 16'hfaf4, 16'hfaf5, 16'hfaf6, 16'hfaf7 	:	val_out <= 16'h7022;
         16'hfaf8, 16'hfaf9, 16'hfafa, 16'hfafb, 16'hfafc, 16'hfafd, 16'hfafe, 16'hfaff 	:	val_out <= 16'h703b;
         16'hfb00, 16'hfb01, 16'hfb02, 16'hfb03, 16'hfb04, 16'hfb05, 16'hfb06, 16'hfb07 	:	val_out <= 16'h7054;
         16'hfb08, 16'hfb09, 16'hfb0a, 16'hfb0b, 16'hfb0c, 16'hfb0d, 16'hfb0e, 16'hfb0f 	:	val_out <= 16'h706d;
         16'hfb10, 16'hfb11, 16'hfb12, 16'hfb13, 16'hfb14, 16'hfb15, 16'hfb16, 16'hfb17 	:	val_out <= 16'h7086;
         16'hfb18, 16'hfb19, 16'hfb1a, 16'hfb1b, 16'hfb1c, 16'hfb1d, 16'hfb1e, 16'hfb1f 	:	val_out <= 16'h709f;
         16'hfb20, 16'hfb21, 16'hfb22, 16'hfb23, 16'hfb24, 16'hfb25, 16'hfb26, 16'hfb27 	:	val_out <= 16'h70b8;
         16'hfb28, 16'hfb29, 16'hfb2a, 16'hfb2b, 16'hfb2c, 16'hfb2d, 16'hfb2e, 16'hfb2f 	:	val_out <= 16'h70d1;
         16'hfb30, 16'hfb31, 16'hfb32, 16'hfb33, 16'hfb34, 16'hfb35, 16'hfb36, 16'hfb37 	:	val_out <= 16'h70ea;
         16'hfb38, 16'hfb39, 16'hfb3a, 16'hfb3b, 16'hfb3c, 16'hfb3d, 16'hfb3e, 16'hfb3f 	:	val_out <= 16'h7103;
         16'hfb40, 16'hfb41, 16'hfb42, 16'hfb43, 16'hfb44, 16'hfb45, 16'hfb46, 16'hfb47 	:	val_out <= 16'h711c;
         16'hfb48, 16'hfb49, 16'hfb4a, 16'hfb4b, 16'hfb4c, 16'hfb4d, 16'hfb4e, 16'hfb4f 	:	val_out <= 16'h7135;
         16'hfb50, 16'hfb51, 16'hfb52, 16'hfb53, 16'hfb54, 16'hfb55, 16'hfb56, 16'hfb57 	:	val_out <= 16'h714e;
         16'hfb58, 16'hfb59, 16'hfb5a, 16'hfb5b, 16'hfb5c, 16'hfb5d, 16'hfb5e, 16'hfb5f 	:	val_out <= 16'h7167;
         16'hfb60, 16'hfb61, 16'hfb62, 16'hfb63, 16'hfb64, 16'hfb65, 16'hfb66, 16'hfb67 	:	val_out <= 16'h7180;
         16'hfb68, 16'hfb69, 16'hfb6a, 16'hfb6b, 16'hfb6c, 16'hfb6d, 16'hfb6e, 16'hfb6f 	:	val_out <= 16'h7199;
         16'hfb70, 16'hfb71, 16'hfb72, 16'hfb73, 16'hfb74, 16'hfb75, 16'hfb76, 16'hfb77 	:	val_out <= 16'h71b2;
         16'hfb78, 16'hfb79, 16'hfb7a, 16'hfb7b, 16'hfb7c, 16'hfb7d, 16'hfb7e, 16'hfb7f 	:	val_out <= 16'h71cb;
         16'hfb80, 16'hfb81, 16'hfb82, 16'hfb83, 16'hfb84, 16'hfb85, 16'hfb86, 16'hfb87 	:	val_out <= 16'h71e4;
         16'hfb88, 16'hfb89, 16'hfb8a, 16'hfb8b, 16'hfb8c, 16'hfb8d, 16'hfb8e, 16'hfb8f 	:	val_out <= 16'h71fd;
         16'hfb90, 16'hfb91, 16'hfb92, 16'hfb93, 16'hfb94, 16'hfb95, 16'hfb96, 16'hfb97 	:	val_out <= 16'h7216;
         16'hfb98, 16'hfb99, 16'hfb9a, 16'hfb9b, 16'hfb9c, 16'hfb9d, 16'hfb9e, 16'hfb9f 	:	val_out <= 16'h722f;
         16'hfba0, 16'hfba1, 16'hfba2, 16'hfba3, 16'hfba4, 16'hfba5, 16'hfba6, 16'hfba7 	:	val_out <= 16'h7248;
         16'hfba8, 16'hfba9, 16'hfbaa, 16'hfbab, 16'hfbac, 16'hfbad, 16'hfbae, 16'hfbaf 	:	val_out <= 16'h7261;
         16'hfbb0, 16'hfbb1, 16'hfbb2, 16'hfbb3, 16'hfbb4, 16'hfbb5, 16'hfbb6, 16'hfbb7 	:	val_out <= 16'h727a;
         16'hfbb8, 16'hfbb9, 16'hfbba, 16'hfbbb, 16'hfbbc, 16'hfbbd, 16'hfbbe, 16'hfbbf 	:	val_out <= 16'h7293;
         16'hfbc0, 16'hfbc1, 16'hfbc2, 16'hfbc3, 16'hfbc4, 16'hfbc5, 16'hfbc6, 16'hfbc7 	:	val_out <= 16'h72ac;
         16'hfbc8, 16'hfbc9, 16'hfbca, 16'hfbcb, 16'hfbcc, 16'hfbcd, 16'hfbce, 16'hfbcf 	:	val_out <= 16'h72c5;
         16'hfbd0, 16'hfbd1, 16'hfbd2, 16'hfbd3, 16'hfbd4, 16'hfbd5, 16'hfbd6, 16'hfbd7 	:	val_out <= 16'h72de;
         16'hfbd8, 16'hfbd9, 16'hfbda, 16'hfbdb, 16'hfbdc, 16'hfbdd, 16'hfbde, 16'hfbdf 	:	val_out <= 16'h72f7;
         16'hfbe0, 16'hfbe1, 16'hfbe2, 16'hfbe3, 16'hfbe4, 16'hfbe5, 16'hfbe6, 16'hfbe7 	:	val_out <= 16'h7310;
         16'hfbe8, 16'hfbe9, 16'hfbea, 16'hfbeb, 16'hfbec, 16'hfbed, 16'hfbee, 16'hfbef 	:	val_out <= 16'h7329;
         16'hfbf0, 16'hfbf1, 16'hfbf2, 16'hfbf3, 16'hfbf4, 16'hfbf5, 16'hfbf6, 16'hfbf7 	:	val_out <= 16'h7342;
         16'hfbf8, 16'hfbf9, 16'hfbfa, 16'hfbfb, 16'hfbfc, 16'hfbfd, 16'hfbfe, 16'hfbff 	:	val_out <= 16'h735b;
         16'hfc00, 16'hfc01, 16'hfc02, 16'hfc03, 16'hfc04, 16'hfc05, 16'hfc06, 16'hfc07 	:	val_out <= 16'h7374;
         16'hfc08, 16'hfc09, 16'hfc0a, 16'hfc0b, 16'hfc0c, 16'hfc0d, 16'hfc0e, 16'hfc0f 	:	val_out <= 16'h738d;
         16'hfc10, 16'hfc11, 16'hfc12, 16'hfc13, 16'hfc14, 16'hfc15, 16'hfc16, 16'hfc17 	:	val_out <= 16'h73a6;
         16'hfc18, 16'hfc19, 16'hfc1a, 16'hfc1b, 16'hfc1c, 16'hfc1d, 16'hfc1e, 16'hfc1f 	:	val_out <= 16'h73bf;
         16'hfc20, 16'hfc21, 16'hfc22, 16'hfc23, 16'hfc24, 16'hfc25, 16'hfc26, 16'hfc27 	:	val_out <= 16'h73d8;
         16'hfc28, 16'hfc29, 16'hfc2a, 16'hfc2b, 16'hfc2c, 16'hfc2d, 16'hfc2e, 16'hfc2f 	:	val_out <= 16'h73f1;
         16'hfc30, 16'hfc31, 16'hfc32, 16'hfc33, 16'hfc34, 16'hfc35, 16'hfc36, 16'hfc37 	:	val_out <= 16'h740a;
         16'hfc38, 16'hfc39, 16'hfc3a, 16'hfc3b, 16'hfc3c, 16'hfc3d, 16'hfc3e, 16'hfc3f 	:	val_out <= 16'h7423;
         16'hfc40, 16'hfc41, 16'hfc42, 16'hfc43, 16'hfc44, 16'hfc45, 16'hfc46, 16'hfc47 	:	val_out <= 16'h743c;
         16'hfc48, 16'hfc49, 16'hfc4a, 16'hfc4b, 16'hfc4c, 16'hfc4d, 16'hfc4e, 16'hfc4f 	:	val_out <= 16'h7455;
         16'hfc50, 16'hfc51, 16'hfc52, 16'hfc53, 16'hfc54, 16'hfc55, 16'hfc56, 16'hfc57 	:	val_out <= 16'h746e;
         16'hfc58, 16'hfc59, 16'hfc5a, 16'hfc5b, 16'hfc5c, 16'hfc5d, 16'hfc5e, 16'hfc5f 	:	val_out <= 16'h7487;
         16'hfc60, 16'hfc61, 16'hfc62, 16'hfc63, 16'hfc64, 16'hfc65, 16'hfc66, 16'hfc67 	:	val_out <= 16'h74a0;
         16'hfc68, 16'hfc69, 16'hfc6a, 16'hfc6b, 16'hfc6c, 16'hfc6d, 16'hfc6e, 16'hfc6f 	:	val_out <= 16'h74b9;
         16'hfc70, 16'hfc71, 16'hfc72, 16'hfc73, 16'hfc74, 16'hfc75, 16'hfc76, 16'hfc77 	:	val_out <= 16'h74d2;
         16'hfc78, 16'hfc79, 16'hfc7a, 16'hfc7b, 16'hfc7c, 16'hfc7d, 16'hfc7e, 16'hfc7f 	:	val_out <= 16'h74eb;
         16'hfc80, 16'hfc81, 16'hfc82, 16'hfc83, 16'hfc84, 16'hfc85, 16'hfc86, 16'hfc87 	:	val_out <= 16'h7504;
         16'hfc88, 16'hfc89, 16'hfc8a, 16'hfc8b, 16'hfc8c, 16'hfc8d, 16'hfc8e, 16'hfc8f 	:	val_out <= 16'h751d;
         16'hfc90, 16'hfc91, 16'hfc92, 16'hfc93, 16'hfc94, 16'hfc95, 16'hfc96, 16'hfc97 	:	val_out <= 16'h7536;
         16'hfc98, 16'hfc99, 16'hfc9a, 16'hfc9b, 16'hfc9c, 16'hfc9d, 16'hfc9e, 16'hfc9f 	:	val_out <= 16'h754f;
         16'hfca0, 16'hfca1, 16'hfca2, 16'hfca3, 16'hfca4, 16'hfca5, 16'hfca6, 16'hfca7 	:	val_out <= 16'h7568;
         16'hfca8, 16'hfca9, 16'hfcaa, 16'hfcab, 16'hfcac, 16'hfcad, 16'hfcae, 16'hfcaf 	:	val_out <= 16'h7581;
         16'hfcb0, 16'hfcb1, 16'hfcb2, 16'hfcb3, 16'hfcb4, 16'hfcb5, 16'hfcb6, 16'hfcb7 	:	val_out <= 16'h759a;
         16'hfcb8, 16'hfcb9, 16'hfcba, 16'hfcbb, 16'hfcbc, 16'hfcbd, 16'hfcbe, 16'hfcbf 	:	val_out <= 16'h75b3;
         16'hfcc0, 16'hfcc1, 16'hfcc2, 16'hfcc3, 16'hfcc4, 16'hfcc5, 16'hfcc6, 16'hfcc7 	:	val_out <= 16'h75cc;
         16'hfcc8, 16'hfcc9, 16'hfcca, 16'hfccb, 16'hfccc, 16'hfccd, 16'hfcce, 16'hfccf 	:	val_out <= 16'h75e6;
         16'hfcd0, 16'hfcd1, 16'hfcd2, 16'hfcd3, 16'hfcd4, 16'hfcd5, 16'hfcd6, 16'hfcd7 	:	val_out <= 16'h75ff;
         16'hfcd8, 16'hfcd9, 16'hfcda, 16'hfcdb, 16'hfcdc, 16'hfcdd, 16'hfcde, 16'hfcdf 	:	val_out <= 16'h7618;
         16'hfce0, 16'hfce1, 16'hfce2, 16'hfce3, 16'hfce4, 16'hfce5, 16'hfce6, 16'hfce7 	:	val_out <= 16'h7631;
         16'hfce8, 16'hfce9, 16'hfcea, 16'hfceb, 16'hfcec, 16'hfced, 16'hfcee, 16'hfcef 	:	val_out <= 16'h764a;
         16'hfcf0, 16'hfcf1, 16'hfcf2, 16'hfcf3, 16'hfcf4, 16'hfcf5, 16'hfcf6, 16'hfcf7 	:	val_out <= 16'h7663;
         16'hfcf8, 16'hfcf9, 16'hfcfa, 16'hfcfb, 16'hfcfc, 16'hfcfd, 16'hfcfe, 16'hfcff 	:	val_out <= 16'h767c;
         16'hfd00, 16'hfd01, 16'hfd02, 16'hfd03, 16'hfd04, 16'hfd05, 16'hfd06, 16'hfd07 	:	val_out <= 16'h7695;
         16'hfd08, 16'hfd09, 16'hfd0a, 16'hfd0b, 16'hfd0c, 16'hfd0d, 16'hfd0e, 16'hfd0f 	:	val_out <= 16'h76ae;
         16'hfd10, 16'hfd11, 16'hfd12, 16'hfd13, 16'hfd14, 16'hfd15, 16'hfd16, 16'hfd17 	:	val_out <= 16'h76c7;
         16'hfd18, 16'hfd19, 16'hfd1a, 16'hfd1b, 16'hfd1c, 16'hfd1d, 16'hfd1e, 16'hfd1f 	:	val_out <= 16'h76e0;
         16'hfd20, 16'hfd21, 16'hfd22, 16'hfd23, 16'hfd24, 16'hfd25, 16'hfd26, 16'hfd27 	:	val_out <= 16'h76f9;
         16'hfd28, 16'hfd29, 16'hfd2a, 16'hfd2b, 16'hfd2c, 16'hfd2d, 16'hfd2e, 16'hfd2f 	:	val_out <= 16'h7712;
         16'hfd30, 16'hfd31, 16'hfd32, 16'hfd33, 16'hfd34, 16'hfd35, 16'hfd36, 16'hfd37 	:	val_out <= 16'h772b;
         16'hfd38, 16'hfd39, 16'hfd3a, 16'hfd3b, 16'hfd3c, 16'hfd3d, 16'hfd3e, 16'hfd3f 	:	val_out <= 16'h7744;
         16'hfd40, 16'hfd41, 16'hfd42, 16'hfd43, 16'hfd44, 16'hfd45, 16'hfd46, 16'hfd47 	:	val_out <= 16'h775d;
         16'hfd48, 16'hfd49, 16'hfd4a, 16'hfd4b, 16'hfd4c, 16'hfd4d, 16'hfd4e, 16'hfd4f 	:	val_out <= 16'h7777;
         16'hfd50, 16'hfd51, 16'hfd52, 16'hfd53, 16'hfd54, 16'hfd55, 16'hfd56, 16'hfd57 	:	val_out <= 16'h7790;
         16'hfd58, 16'hfd59, 16'hfd5a, 16'hfd5b, 16'hfd5c, 16'hfd5d, 16'hfd5e, 16'hfd5f 	:	val_out <= 16'h77a9;
         16'hfd60, 16'hfd61, 16'hfd62, 16'hfd63, 16'hfd64, 16'hfd65, 16'hfd66, 16'hfd67 	:	val_out <= 16'h77c2;
         16'hfd68, 16'hfd69, 16'hfd6a, 16'hfd6b, 16'hfd6c, 16'hfd6d, 16'hfd6e, 16'hfd6f 	:	val_out <= 16'h77db;
         16'hfd70, 16'hfd71, 16'hfd72, 16'hfd73, 16'hfd74, 16'hfd75, 16'hfd76, 16'hfd77 	:	val_out <= 16'h77f4;
         16'hfd78, 16'hfd79, 16'hfd7a, 16'hfd7b, 16'hfd7c, 16'hfd7d, 16'hfd7e, 16'hfd7f 	:	val_out <= 16'h780d;
         16'hfd80, 16'hfd81, 16'hfd82, 16'hfd83, 16'hfd84, 16'hfd85, 16'hfd86, 16'hfd87 	:	val_out <= 16'h7826;
         16'hfd88, 16'hfd89, 16'hfd8a, 16'hfd8b, 16'hfd8c, 16'hfd8d, 16'hfd8e, 16'hfd8f 	:	val_out <= 16'h783f;
         16'hfd90, 16'hfd91, 16'hfd92, 16'hfd93, 16'hfd94, 16'hfd95, 16'hfd96, 16'hfd97 	:	val_out <= 16'h7858;
         16'hfd98, 16'hfd99, 16'hfd9a, 16'hfd9b, 16'hfd9c, 16'hfd9d, 16'hfd9e, 16'hfd9f 	:	val_out <= 16'h7871;
         16'hfda0, 16'hfda1, 16'hfda2, 16'hfda3, 16'hfda4, 16'hfda5, 16'hfda6, 16'hfda7 	:	val_out <= 16'h788a;
         16'hfda8, 16'hfda9, 16'hfdaa, 16'hfdab, 16'hfdac, 16'hfdad, 16'hfdae, 16'hfdaf 	:	val_out <= 16'h78a4;
         16'hfdb0, 16'hfdb1, 16'hfdb2, 16'hfdb3, 16'hfdb4, 16'hfdb5, 16'hfdb6, 16'hfdb7 	:	val_out <= 16'h78bd;
         16'hfdb8, 16'hfdb9, 16'hfdba, 16'hfdbb, 16'hfdbc, 16'hfdbd, 16'hfdbe, 16'hfdbf 	:	val_out <= 16'h78d6;
         16'hfdc0, 16'hfdc1, 16'hfdc2, 16'hfdc3, 16'hfdc4, 16'hfdc5, 16'hfdc6, 16'hfdc7 	:	val_out <= 16'h78ef;
         16'hfdc8, 16'hfdc9, 16'hfdca, 16'hfdcb, 16'hfdcc, 16'hfdcd, 16'hfdce, 16'hfdcf 	:	val_out <= 16'h7908;
         16'hfdd0, 16'hfdd1, 16'hfdd2, 16'hfdd3, 16'hfdd4, 16'hfdd5, 16'hfdd6, 16'hfdd7 	:	val_out <= 16'h7921;
         16'hfdd8, 16'hfdd9, 16'hfdda, 16'hfddb, 16'hfddc, 16'hfddd, 16'hfdde, 16'hfddf 	:	val_out <= 16'h793a;
         16'hfde0, 16'hfde1, 16'hfde2, 16'hfde3, 16'hfde4, 16'hfde5, 16'hfde6, 16'hfde7 	:	val_out <= 16'h7953;
         16'hfde8, 16'hfde9, 16'hfdea, 16'hfdeb, 16'hfdec, 16'hfded, 16'hfdee, 16'hfdef 	:	val_out <= 16'h796c;
         16'hfdf0, 16'hfdf1, 16'hfdf2, 16'hfdf3, 16'hfdf4, 16'hfdf5, 16'hfdf6, 16'hfdf7 	:	val_out <= 16'h7985;
         16'hfdf8, 16'hfdf9, 16'hfdfa, 16'hfdfb, 16'hfdfc, 16'hfdfd, 16'hfdfe, 16'hfdff 	:	val_out <= 16'h799f;
         16'hfe00, 16'hfe01, 16'hfe02, 16'hfe03, 16'hfe04, 16'hfe05, 16'hfe06, 16'hfe07 	:	val_out <= 16'h79b8;
         16'hfe08, 16'hfe09, 16'hfe0a, 16'hfe0b, 16'hfe0c, 16'hfe0d, 16'hfe0e, 16'hfe0f 	:	val_out <= 16'h79d1;
         16'hfe10, 16'hfe11, 16'hfe12, 16'hfe13, 16'hfe14, 16'hfe15, 16'hfe16, 16'hfe17 	:	val_out <= 16'h79ea;
         16'hfe18, 16'hfe19, 16'hfe1a, 16'hfe1b, 16'hfe1c, 16'hfe1d, 16'hfe1e, 16'hfe1f 	:	val_out <= 16'h7a03;
         16'hfe20, 16'hfe21, 16'hfe22, 16'hfe23, 16'hfe24, 16'hfe25, 16'hfe26, 16'hfe27 	:	val_out <= 16'h7a1c;
         16'hfe28, 16'hfe29, 16'hfe2a, 16'hfe2b, 16'hfe2c, 16'hfe2d, 16'hfe2e, 16'hfe2f 	:	val_out <= 16'h7a35;
         16'hfe30, 16'hfe31, 16'hfe32, 16'hfe33, 16'hfe34, 16'hfe35, 16'hfe36, 16'hfe37 	:	val_out <= 16'h7a4e;
         16'hfe38, 16'hfe39, 16'hfe3a, 16'hfe3b, 16'hfe3c, 16'hfe3d, 16'hfe3e, 16'hfe3f 	:	val_out <= 16'h7a67;
         16'hfe40, 16'hfe41, 16'hfe42, 16'hfe43, 16'hfe44, 16'hfe45, 16'hfe46, 16'hfe47 	:	val_out <= 16'h7a80;
         16'hfe48, 16'hfe49, 16'hfe4a, 16'hfe4b, 16'hfe4c, 16'hfe4d, 16'hfe4e, 16'hfe4f 	:	val_out <= 16'h7a9a;
         16'hfe50, 16'hfe51, 16'hfe52, 16'hfe53, 16'hfe54, 16'hfe55, 16'hfe56, 16'hfe57 	:	val_out <= 16'h7ab3;
         16'hfe58, 16'hfe59, 16'hfe5a, 16'hfe5b, 16'hfe5c, 16'hfe5d, 16'hfe5e, 16'hfe5f 	:	val_out <= 16'h7acc;
         16'hfe60, 16'hfe61, 16'hfe62, 16'hfe63, 16'hfe64, 16'hfe65, 16'hfe66, 16'hfe67 	:	val_out <= 16'h7ae5;
         16'hfe68, 16'hfe69, 16'hfe6a, 16'hfe6b, 16'hfe6c, 16'hfe6d, 16'hfe6e, 16'hfe6f 	:	val_out <= 16'h7afe;
         16'hfe70, 16'hfe71, 16'hfe72, 16'hfe73, 16'hfe74, 16'hfe75, 16'hfe76, 16'hfe77 	:	val_out <= 16'h7b17;
         16'hfe78, 16'hfe79, 16'hfe7a, 16'hfe7b, 16'hfe7c, 16'hfe7d, 16'hfe7e, 16'hfe7f 	:	val_out <= 16'h7b30;
         16'hfe80, 16'hfe81, 16'hfe82, 16'hfe83, 16'hfe84, 16'hfe85, 16'hfe86, 16'hfe87 	:	val_out <= 16'h7b49;
         16'hfe88, 16'hfe89, 16'hfe8a, 16'hfe8b, 16'hfe8c, 16'hfe8d, 16'hfe8e, 16'hfe8f 	:	val_out <= 16'h7b63;
         16'hfe90, 16'hfe91, 16'hfe92, 16'hfe93, 16'hfe94, 16'hfe95, 16'hfe96, 16'hfe97 	:	val_out <= 16'h7b7c;
         16'hfe98, 16'hfe99, 16'hfe9a, 16'hfe9b, 16'hfe9c, 16'hfe9d, 16'hfe9e, 16'hfe9f 	:	val_out <= 16'h7b95;
         16'hfea0, 16'hfea1, 16'hfea2, 16'hfea3, 16'hfea4, 16'hfea5, 16'hfea6, 16'hfea7 	:	val_out <= 16'h7bae;
         16'hfea8, 16'hfea9, 16'hfeaa, 16'hfeab, 16'hfeac, 16'hfead, 16'hfeae, 16'hfeaf 	:	val_out <= 16'h7bc7;
         16'hfeb0, 16'hfeb1, 16'hfeb2, 16'hfeb3, 16'hfeb4, 16'hfeb5, 16'hfeb6, 16'hfeb7 	:	val_out <= 16'h7be0;
         16'hfeb8, 16'hfeb9, 16'hfeba, 16'hfebb, 16'hfebc, 16'hfebd, 16'hfebe, 16'hfebf 	:	val_out <= 16'h7bf9;
         16'hfec0, 16'hfec1, 16'hfec2, 16'hfec3, 16'hfec4, 16'hfec5, 16'hfec6, 16'hfec7 	:	val_out <= 16'h7c12;
         16'hfec8, 16'hfec9, 16'hfeca, 16'hfecb, 16'hfecc, 16'hfecd, 16'hfece, 16'hfecf 	:	val_out <= 16'h7c2b;
         16'hfed0, 16'hfed1, 16'hfed2, 16'hfed3, 16'hfed4, 16'hfed5, 16'hfed6, 16'hfed7 	:	val_out <= 16'h7c45;
         16'hfed8, 16'hfed9, 16'hfeda, 16'hfedb, 16'hfedc, 16'hfedd, 16'hfede, 16'hfedf 	:	val_out <= 16'h7c5e;
         16'hfee0, 16'hfee1, 16'hfee2, 16'hfee3, 16'hfee4, 16'hfee5, 16'hfee6, 16'hfee7 	:	val_out <= 16'h7c77;
         16'hfee8, 16'hfee9, 16'hfeea, 16'hfeeb, 16'hfeec, 16'hfeed, 16'hfeee, 16'hfeef 	:	val_out <= 16'h7c90;
         16'hfef0, 16'hfef1, 16'hfef2, 16'hfef3, 16'hfef4, 16'hfef5, 16'hfef6, 16'hfef7 	:	val_out <= 16'h7ca9;
         16'hfef8, 16'hfef9, 16'hfefa, 16'hfefb, 16'hfefc, 16'hfefd, 16'hfefe, 16'hfeff 	:	val_out <= 16'h7cc2;
         16'hff00, 16'hff01, 16'hff02, 16'hff03, 16'hff04, 16'hff05, 16'hff06, 16'hff07 	:	val_out <= 16'h7cdb;
         16'hff08, 16'hff09, 16'hff0a, 16'hff0b, 16'hff0c, 16'hff0d, 16'hff0e, 16'hff0f 	:	val_out <= 16'h7cf4;
         16'hff10, 16'hff11, 16'hff12, 16'hff13, 16'hff14, 16'hff15, 16'hff16, 16'hff17 	:	val_out <= 16'h7d0e;
         16'hff18, 16'hff19, 16'hff1a, 16'hff1b, 16'hff1c, 16'hff1d, 16'hff1e, 16'hff1f 	:	val_out <= 16'h7d27;
         16'hff20, 16'hff21, 16'hff22, 16'hff23, 16'hff24, 16'hff25, 16'hff26, 16'hff27 	:	val_out <= 16'h7d40;
         16'hff28, 16'hff29, 16'hff2a, 16'hff2b, 16'hff2c, 16'hff2d, 16'hff2e, 16'hff2f 	:	val_out <= 16'h7d59;
         16'hff30, 16'hff31, 16'hff32, 16'hff33, 16'hff34, 16'hff35, 16'hff36, 16'hff37 	:	val_out <= 16'h7d72;
         16'hff38, 16'hff39, 16'hff3a, 16'hff3b, 16'hff3c, 16'hff3d, 16'hff3e, 16'hff3f 	:	val_out <= 16'h7d8b;
         16'hff40, 16'hff41, 16'hff42, 16'hff43, 16'hff44, 16'hff45, 16'hff46, 16'hff47 	:	val_out <= 16'h7da4;
         16'hff48, 16'hff49, 16'hff4a, 16'hff4b, 16'hff4c, 16'hff4d, 16'hff4e, 16'hff4f 	:	val_out <= 16'h7dbd;
         16'hff50, 16'hff51, 16'hff52, 16'hff53, 16'hff54, 16'hff55, 16'hff56, 16'hff57 	:	val_out <= 16'h7dd7;
         16'hff58, 16'hff59, 16'hff5a, 16'hff5b, 16'hff5c, 16'hff5d, 16'hff5e, 16'hff5f 	:	val_out <= 16'h7df0;
         16'hff60, 16'hff61, 16'hff62, 16'hff63, 16'hff64, 16'hff65, 16'hff66, 16'hff67 	:	val_out <= 16'h7e09;
         16'hff68, 16'hff69, 16'hff6a, 16'hff6b, 16'hff6c, 16'hff6d, 16'hff6e, 16'hff6f 	:	val_out <= 16'h7e22;
         16'hff70, 16'hff71, 16'hff72, 16'hff73, 16'hff74, 16'hff75, 16'hff76, 16'hff77 	:	val_out <= 16'h7e3b;
         16'hff78, 16'hff79, 16'hff7a, 16'hff7b, 16'hff7c, 16'hff7d, 16'hff7e, 16'hff7f 	:	val_out <= 16'h7e54;
         16'hff80, 16'hff81, 16'hff82, 16'hff83, 16'hff84, 16'hff85, 16'hff86, 16'hff87 	:	val_out <= 16'h7e6d;
         16'hff88, 16'hff89, 16'hff8a, 16'hff8b, 16'hff8c, 16'hff8d, 16'hff8e, 16'hff8f 	:	val_out <= 16'h7e87;
         16'hff90, 16'hff91, 16'hff92, 16'hff93, 16'hff94, 16'hff95, 16'hff96, 16'hff97 	:	val_out <= 16'h7ea0;
         16'hff98, 16'hff99, 16'hff9a, 16'hff9b, 16'hff9c, 16'hff9d, 16'hff9e, 16'hff9f 	:	val_out <= 16'h7eb9;
         16'hffa0, 16'hffa1, 16'hffa2, 16'hffa3, 16'hffa4, 16'hffa5, 16'hffa6, 16'hffa7 	:	val_out <= 16'h7ed2;
         16'hffa8, 16'hffa9, 16'hffaa, 16'hffab, 16'hffac, 16'hffad, 16'hffae, 16'hffaf 	:	val_out <= 16'h7eeb;
         16'hffb0, 16'hffb1, 16'hffb2, 16'hffb3, 16'hffb4, 16'hffb5, 16'hffb6, 16'hffb7 	:	val_out <= 16'h7f04;
         16'hffb8, 16'hffb9, 16'hffba, 16'hffbb, 16'hffbc, 16'hffbd, 16'hffbe, 16'hffbf 	:	val_out <= 16'h7f1d;
         16'hffc0, 16'hffc1, 16'hffc2, 16'hffc3, 16'hffc4, 16'hffc5, 16'hffc6, 16'hffc7 	:	val_out <= 16'h7f36;
         16'hffc8, 16'hffc9, 16'hffca, 16'hffcb, 16'hffcc, 16'hffcd, 16'hffce, 16'hffcf 	:	val_out <= 16'h7f50;
         16'hffd0, 16'hffd1, 16'hffd2, 16'hffd3, 16'hffd4, 16'hffd5, 16'hffd6, 16'hffd7 	:	val_out <= 16'h7f69;
         16'hffd8, 16'hffd9, 16'hffda, 16'hffdb, 16'hffdc, 16'hffdd, 16'hffde, 16'hffdf 	:	val_out <= 16'h7f82;
         16'hffe0, 16'hffe1, 16'hffe2, 16'hffe3, 16'hffe4, 16'hffe5, 16'hffe6, 16'hffe7 	:	val_out <= 16'h7f9b;
         16'hffe8, 16'hffe9, 16'hffea, 16'hffeb, 16'hffec, 16'hffed, 16'hffee, 16'hffef 	:	val_out <= 16'h7fb4;
         16'hfff0, 16'hfff1, 16'hfff2, 16'hfff3, 16'hfff4, 16'hfff5, 16'hfff6, 16'hfff7 	:	val_out <= 16'h7fcd;
         16'hfff8, 16'hfff9, 16'hfffa, 16'hfffb, 16'hfffc, 16'hfffd, 16'hfffe, 16'hffff 	:	val_out <= 16'h7fe6;
			default	:	val_out <= 16'h0;
		endcase
	end
endmodule
