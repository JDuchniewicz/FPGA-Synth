// Pipelined State variable filter based on Andrew Simper's SVF whitepaper https://cytomic.com/files/dsp/SvfLinearTrapOptimised2.pdf

module state_variable_filter_iir_p(input clk,
											input clk_en,
											input rst,
											input[6:0] i_midi,
											output reg[6:0] o_midi,
											input signed[23:0] i_data,
											input i_valid,
											output reg o_valid,
											output reg signed[23:0] o_filtered // == v2
											);
	parameter NBANKS = 10;
	
	reg signed[39:0] v1[NBANKS-1:0];
	reg signed[39:0] v2[NBANKS-1:0];
	reg signed[39:0] v3[NBANKS-1:0];
	reg signed[39:0] ic1eq[NBANKS-1:0];
	reg signed[39:0] ic2eq[NBANKS-1:0];
	
	wire signed[39:0] w_a1, w_a2, w_a3;
	wire signed[79:0] mR_0, mR_1, mR_2, mR_3;
	
	reg signed[39:0] r_m_a1, r_m_a2, r_m_a3, r_m_ic1eq, r_m_v3;
	
	// for buffering values
	reg valid[1:0];
	reg[6:0] midi[1:0];
	
	wire signed[39:0] w_extended_i_data;
	
	coefficients_lut lut(.i_midi(i_midi), 
								.o_a1(w_a1),
								.o_a2(w_a2), 
								.o_a3(w_a3));
								
	lpm_multiplier 
						mult0(.dataa(r_m_a1), // first try with higher precision, then decrease to 32 bits and try again?
								.datab(r_m_ic1eq),
								.result(mR_0)),
						mult1(.dataa(r_m_a2), 
								.datab(r_m_v3), 
								.result(mR_1)),
						mult2(.dataa(r_m_a2), 
								.datab(r_m_ic1eq), 
								.result(mR_2)),
						mult3(.dataa(r_m_a3), 
								.datab(r_m_v3), 
								.result(mR_3));
								
	integer v_idx;
	integer i;
	
	assign w_extended_i_data = {{3{i_data[23]}}, {i_data[22:0]}, 14'b0};

	initial begin
		for (i = 0; i < NBANKS; i = i + 1) begin
			v1[i] = 40'b0;
			v2[i] = 40'b0;
			v3[i] = 40'b0;
			ic1eq[i] = 40'b0;
			ic2eq[i] = 40'b0;
		end
		for (i = 0; i < 2; i = i + 1) begin
			valid[i] = 1'b0;
			midi[i] = 7'b0;
		end
		r_m_a1 = 40'b0;
		r_m_a2 = 40'b0;
		r_m_a3 = 40'b0;
		r_m_ic1eq = 40'b0;
		r_m_v3 = 40'b0;

		v_idx = 5;
	end
	
	always @(posedge clk or posedge rst) begin
		if (rst) begin // what about passthrough midi value?
			for (i = 0; i < NBANKS; i = i + 1) begin
				v1[i] <= 40'b0;
				v2[i] <= 40'b0;
				v3[i] <= 40'b0;
				ic1eq[i] <= 40'b0;
				ic2eq[i] <= 40'b0;		
			end
			for (i = 0; i < 2; i = i + 1) begin
				valid[i] <= 1'b0;
				midi[i] <= 7'b0;
			end
			r_m_a1 <= 40'b0;
			r_m_a2 <= 40'b0;
			r_m_a3 <= 40'b0;
			r_m_ic1eq <= 40'b0;
			r_m_v3 <= 40'b0;

			v_idx <= 5;
		end else if (clk_en) begin
			// three cycles of delay - sine-like solution
			// first cycle calc coefficients -> clear registers if midi 00
			if (i_midi == 7'b0) begin
				v1[v_idx] <= 40'b0;
				v2[v_idx] <= 40'b0;
				v3[v_idx] <= 40'b0;
				ic1eq[v_idx] <= 40'b0;
				ic2eq[v_idx] <= 40'b0;
				// fill the lpm_multiplier
				r_m_a1 <= 40'b0;
				r_m_a2 <= 40'b0;
				r_m_a3 <= 40'b0;
				r_m_ic1eq <= 40'b0;
				r_m_v3 <= 40'b0;
			end else begin
				// fill the lpm_multiplier
				r_m_a1 <= w_a1;
				r_m_a2 <= w_a2;
				r_m_a3 <= w_a3;
				r_m_ic1eq <= ic1eq[v_idx];
				r_m_v3 <= w_extended_i_data - ic2eq[v_idx]; // to prevent 1 cycle delay
				// filter step
				v3[v_idx] <= w_extended_i_data - ic2eq[v_idx];
			end
			
			// second cycle -> obtain multiplication results
			if (v_idx == 0) begin
				v1[NBANKS - 1] <= (mR_0 >>> 37) + (mR_1 >>> 37); // remove scaling factor due to multiplication  (probably need to take a slice out of it, truncates automatically)
				v2[NBANKS - 1] <= ic2eq[NBANKS - 1] + (mR_2 >>> 37) + (mR_3 >>> 37); // should this be a shift or (TODO: this could probably need a greater width...?)
			end else begin
				v1[v_idx - 1] <= (mR_0 >>> 37) + (mR_1 >>> 37);
				v2[v_idx - 1] <= ic2eq[v_idx - 1] + (mR_2 >>> 37) + (mR_3 >>> 37);
			end

			// third cycle -> last steps and output result
			if (v_idx == 0) begin
				ic1eq[NBANKS - 2] <= (v1[NBANKS - 2] <<< 1) - ic1eq[NBANKS - 2];
				ic2eq[NBANKS - 2] <= (v2[NBANKS - 2] <<< 1) - ic2eq[NBANKS - 2];
				o_filtered <= {v2[NBANKS - 2][39], v2[NBANKS - 2][36:14]};		
			end else if (v_idx == 1) begin
				ic1eq[NBANKS - 1] <= (v1[NBANKS - 1] <<< 1) - ic1eq[NBANKS - 1];
				ic2eq[NBANKS - 1] <= (v2[NBANKS - 1] <<< 1) - ic2eq[NBANKS - 1];
				o_filtered <= {v2[NBANKS - 1][39], v2[NBANKS - 1][36:14]};
			end else begin
				ic1eq[v_idx - 2] <= (v1[v_idx - 2] <<< 1) - ic1eq[v_idx - 2];
				ic2eq[v_idx - 2] <= (v2[v_idx - 2] <<< 1) - ic2eq[v_idx - 2];
				o_filtered <= {v2[v_idx - 2][39], v2[v_idx - 2][36:14]};				
			end
			
			// move valid value
			valid[0] <= i_valid;
			valid[1] <= valid[0];
			o_valid <= valid[1];
			
			// move midi value
			midi[0] <= i_midi;
			midi[1] <= midi[0];
			o_midi <= midi[1];
			
			if (v_idx == NBANKS - 1)
				v_idx <= 0;
			else
				v_idx <= v_idx + 1;
		end
	end

endmodule

// Q2.37 format
module coefficients_lut(input[6:0] i_midi,
								output reg signed[39:0] o_a1,
								output reg signed[39:0] o_a2,
								output reg signed[39:0] o_a3); // q format needed here check maths if are proper, addition substraction and multiplication have to be done
										// check required precision for calculating the output signal etc, when to convert and how v2 -> output signal, input should be rescaled to -1 - 1 range? and to q format?
	initial begin
		o_a1 = 40'b0;
		o_a2 = 40'b0;
		o_a3 = 40'b0;
	end
	
	always @(i_midi) begin
		case (i_midi)
            7'h00 	:	 begin 
                o_a1 <= 40'b0000000000000000000000000000000000000000;
                o_a2 <= 40'b0000000000000000000000000000000000000000;
                o_a3 <= 40'b0000000000000000000000000000000000000000;
                end
            7'h01 	:	 begin 
                o_a1 <= 40'b0001111111100001100101010011110110110001;
                o_a2 <= 40'b0000000000001111001100011100001000111100;
                o_a3 <= 40'b0000000000000000000001110011110111010101;
                end
            7'h02 	:	 begin 
                o_a1 <= 40'b0001111111000010101111000011010111101000;
                o_a2 <= 40'b0000000000011110100100110010110110010001;
                o_a3 <= 40'b0000000000000000000111010110111011110100;
                end
            7'h03 	:	 begin 
                o_a1 <= 40'b0001111110100011011101000001100011111010;
                o_a2 <= 40'b0000000000101110001001000100110111101110;
                o_a3 <= 40'b0000000000000000010000110100101100100111;
                end
            7'h04 	:	 begin 
                o_a1 <= 40'b0001111110000011101111000001110000111001;
                o_a2 <= 40'b0000000000111101111001010010100111001110;
                o_a3 <= 40'b0000000000000000011110011001000000101001;
                end
            7'h05 	:	 begin 
                o_a1 <= 40'b0001111101100011100100110111101000110001;
                o_a2 <= 40'b0000000001001101110101011100001000000111;
                o_a3 <= 40'b0000000000000000110000010000000111000000;
                end
            7'h06 	:	 begin 
                o_a1 <= 40'b0001111101000010111110010111001011100101;
                o_a2 <= 40'b0000000001011101111101100001000110011010;
                o_a3 <= 40'b0000000000000001000110100110100111100101;
                end
            7'h07 	:	 begin 
                o_a1 <= 40'b0001111100100001111011010100110000010001;
                o_a2 <= 40'b0000000001101110010001100000110110000111;
                o_a3 <= 40'b0000000000000001100001101001100011011111;
                end
            7'h08 	:	 begin 
                o_a1 <= 40'b0001111100000000011011100101000101100100;
                o_a2 <= 40'b0000000001111110110001011010010010011011;
                o_a3 <= 40'b0000000000000010000001100110010101100101;
                end
            7'h09 	:	 begin 
                o_a1 <= 40'b0001111011011110011110111101010011000001;
                o_a2 <= 40'b0000000010001111011101001011111100111110;
                o_a3 <= 40'b0000000000000010100110101010110011000000;
                end
            7'h0a 	:	 begin 
                o_a1 <= 40'b0001111010111100000101010010111001111111;
                o_a2 <= 40'b0000000010100000010100110011111101001000;
                o_a3 <= 40'b0000000000000011010001000101001011101111;
                end
            7'h0b 	:	 begin 
                o_a1 <= 40'b0001111010011001001110011011110110101001;
                o_a2 <= 40'b0000000010110001011000001111111111001010;
                o_a3 <= 40'b0000000000000100000001000100001011000001;
                end
            7'h0c 	:	 begin 
                o_a1 <= 40'b0001111001110101111010001110100000111010;
                o_a2 <= 40'b0000000011000010100111011101010011100101;
                o_a3 <= 40'b0000000000000100110110110110110111111011;
                end
            7'h0d 	:	 begin 
                o_a1 <= 40'b0001111001010010001000100001101101100000;
                o_a2 <= 40'b0000000011010100000010011000101110010011;
                o_a3 <= 40'b0000000000000101110010101100110101111000;
                end
            7'h0e 	:	 begin 
                o_a1 <= 40'b0001111000101101111001001100101110111000;
                o_a2 <= 40'b0000000011100101101000111110100101111110;
                o_a3 <= 40'b0000000000000110110100110110000101001011;
                end
            7'h0f 	:	 begin 
                o_a1 <= 40'b0001111000001001001100000111010110001110;
                o_a2 <= 40'b0000000011110111011011001010110011001001;
                o_a3 <= 40'b0000000000000111111101100011000011011110;
                end
            7'h10 	:	 begin 
                o_a1 <= 40'b0001110111100100000001001001110100011101;
                o_a2 <= 40'b0000000100001001011000111000101111101000;
                o_a3 <= 40'b0000000000001001001101000100101100010001;
                end
            7'h11 	:	 begin 
                o_a1 <= 40'b0001110110111110011000001100111011001011;
                o_a2 <= 40'b0000000100011011100010000011010101101000;
                o_a3 <= 40'b0000000000001010100011101100011001100011;
                end
            7'h12 	:	 begin 
                o_a1 <= 40'b0001110110011000010001001001111101100100;
                o_a2 <= 40'b0000000100101101110110100100111111001001;
                o_a3 <= 40'b0000000000001100000001101100000100000111;
                end
            7'h13 	:	 begin 
                o_a1 <= 40'b0001110101110001101011111010110001011100;
                o_a2 <= 40'b0000000101000000010110010111100101001001;
                o_a3 <= 40'b0000000000001101100111010110000100010000;
                end
            7'h14 	:	 begin 
                o_a1 <= 40'b0001110101001010101000011001110000000100;
                o_a2 <= 40'b0000000101010011000001010100011110111001;
                o_a3 <= 40'b0000000000001111010100111101010010001001;
                end
            7'h15 	:	 begin 
                o_a1 <= 40'b0001110100100011000110100001110111001001;
                o_a2 <= 40'b0000000101100101110111010100100001001110;
                o_a3 <= 40'b0000000000010001001010110101000110011001;
                end
            7'h16 	:	 begin 
                o_a1 <= 40'b0001110011111011000110001110101001101011;
                o_a2 <= 40'b0000000101111000111000001111111101110111;
                o_a3 <= 40'b0000000000010011001001010001011010100100;
                end
            7'h17 	:	 begin 
                o_a1 <= 40'b0001110011010010100111011100010000110110;
                o_a2 <= 40'b0000000110001100000011111110100010101111;
                o_a3 <= 40'b0000000000010101010000100110101001101001;
                end
            7'h18 	:	 begin 
                o_a1 <= 40'b0001110010101001101010000111011100110111;
                o_a2 <= 40'b0000000110011111011010010111011001010001;
                o_a3 <= 40'b0000000000010111100001001001110000100100;
                end
            7'h19 	:	 begin 
                o_a1 <= 40'b0001110010000000001110001101100101110001;
                o_a2 <= 40'b0000000110110010111011010001000101110000;
                o_a3 <= 40'b0000000000011001111011010000001110101101;
                end
            7'h1a 	:	 begin 
                o_a1 <= 40'b0001110001010110010011101100101100010010;
                o_a2 <= 40'b0000000111000110100110100001100110101011;
                o_a3 <= 40'b0000000000011100011111010000000110010111;
                end
            7'h1b 	:	 begin 
                o_a1 <= 40'b0001110000101011111010100011011010011111;
                o_a2 <= 40'b0000000111011010011011111110010100000110;
                o_a3 <= 40'b0000000000011111001101011111111101010011;
                end
            7'h1c 	:	 begin 
                o_a1 <= 40'b0001110000000001000010110001000100101010;
                o_a2 <= 40'b0000000111101110011011011011111111000100;
                o_a3 <= 40'b0000000000100010000110010110111101001100;
                end
            7'h1d 	:	 begin 
                o_a1 <= 40'b0001101111010101101100010101101001111000;
                o_a2 <= 40'b0000001000000010100100101110110000111110;
                o_a3 <= 40'b0000000000100101001010001100110100001001;
                end
            7'h1e 	:	 begin 
                o_a1 <= 40'b0001101110101001110111010001110100101111;
                o_a2 <= 40'b0000001000010110110111101010001011000000;
                o_a3 <= 40'b0000000000101000011001011001110101001111;
                end
            7'h1f 	:	 begin 
                o_a1 <= 40'b0001101101111101100011100110111011111010;
                o_a2 <= 40'b0000001000101011010100000001000101100100;
                o_a3 <= 40'b0000000000101011110100010110111000111101;
                end
            7'h20 	:	 begin 
                o_a1 <= 40'b0001101101010000110001010111000010110100;
                o_a2 <= 40'b0000001000111111111001100101101111101111;
                o_a3 <= 40'b0000000000101111011011011101011101101101;
                end
            7'h21 	:	 begin 
                o_a1 <= 40'b0001101100100011100000100100111010000011;
                o_a2 <= 40'b0000001001010100101000001001101110110001;
                o_a3 <= 40'b0000000000110011001111000111101000011000;
                end
            7'h22 	:	 begin 
                o_a1 <= 40'b0001101011110101110001010011111111111010;
                o_a2 <= 40'b0000001001101001011111011101111101101000;
                o_a3 <= 40'b0000000000110111001111110000000100110100;
                end
            7'h23 	:	 begin 
                o_a1 <= 40'b0001101011000111100011101000100000110111;
                o_a2 <= 40'b0000001001111110011111010010101100011001;
                o_a3 <= 40'b0000000000111011011101110010000110010101;
                end
            7'h24 	:	 begin 
                o_a1 <= 40'b0001101010011000110111100111010111110100;
                o_a2 <= 40'b0000001010010011100111010111011111111101;
                o_a3 <= 40'b0000000000111111111001101001101000010001;
                end
            7'h25 	:	 begin 
                o_a1 <= 40'b0001101001101001101101010110001110100010;
                o_a2 <= 40'b0000001010101000110111011011010001011111;
                o_a3 <= 40'b0000000001000100100011110011001110011110;
                end
            7'h26 	:	 begin 
                o_a1 <= 40'b0001101000111010000100111011011101111000;
                o_a2 <= 40'b0000001010111110001111001100001110000101;
                o_a3 <= 40'b0000000001001001011100101100000101111101;
                end
            7'h27 	:	 begin 
                o_a1 <= 40'b0001101000001001111110011110001101111110;
                o_a2 <= 40'b0000001011010011101110010111110110010110;
                o_a3 <= 40'b0000000001001110100100110010000101010101;
                end
            7'h28 	:	 begin 
                o_a1 <= 40'b0001100111011001011010000110010110010101;
                o_a2 <= 40'b0000001011101001010100101010111110000101;
                o_a3 <= 40'b0000000001010011111100100011101101011110;
                end
            7'h29 	:	 begin 
                o_a1 <= 40'b0001100110101000010111111100011110000000;
                o_a2 <= 40'b0000001011111111000001110001101011111011;
                o_a3 <= 40'b0000000001011001100100100000001010000111;
                end
            7'h2a 	:	 begin 
                o_a1 <= 40'b0001100101110110111000001001111011011110;
                o_a2 <= 40'b0000001100010100110101010111011001000010;
                o_a3 <= 40'b0000000001011111011101000111010010011011;
                end
            7'h2b 	:	 begin 
                o_a1 <= 40'b0001100101000100111010111000110100101010;
                o_a2 <= 40'b0000001100101010101111000110110000110100;
                o_a3 <= 40'b0000000001100101100110111001101001101011;
                end
            7'h2c 	:	 begin 
                o_a1 <= 40'b0001100100010010100000010011111110101101;
                o_a2 <= 40'b0000001101000000101110101001110000101010;
                o_a3 <= 40'b0000000001101100000010011000011111111110;
                end
            7'h2d 	:	 begin 
                o_a1 <= 40'b0001100011011111101000100110111101110011;
                o_a2 <= 40'b0000001101010110110011101001100111101010;
                o_a3 <= 40'b0000000001110010110000000101110010110111;
                end
            7'h2e 	:	 begin 
                o_a1 <= 40'b0001100010101100010011111110000100110111;
                o_a2 <= 40'b0000001101101100111101101110110110011111;
                o_a3 <= 40'b0000000001111001110000100100001110001010;
                end
            7'h2f 	:	 begin 
                o_a1 <= 40'b0001100001111000100010100110010101001001;
                o_a2 <= 40'b0000001110000011001100100001001111000100;
                o_a3 <= 40'b0000000010000001000100010111001100101100;
                end
            7'h30 	:	 begin 
                o_a1 <= 40'b0001100001000100010100101101011101110010;
                o_a2 <= 40'b0000001110011001011111100111110100100000;
                o_a3 <= 40'b0000000010001000101100000010111001001011;
                end
            7'h31 	:	 begin 
                o_a1 <= 40'b0001100000001111101010100001111011001110;
                o_a2 <= 40'b0000001110101111110110101000111010110110;
                o_a3 <= 40'b0000000010010000101000001100001111000011;
                end
            7'h32 	:	 begin 
                o_a1 <= 40'b0001011111011010100100010010110110100101;
                o_a2 <= 40'b0000001111000110010001001010000110111101;
                o_a3 <= 40'b0000000010011000111001011000111011011111;
                end
            7'h33 	:	 begin 
                o_a1 <= 40'b0001011110100101000010010000000100111100;
                o_a2 <= 40'b0000001111011100101110110000001110010111;
                o_a3 <= 40'b0000000010100001100000001111011110010101;
                end
            7'h34 	:	 begin 
                o_a1 <= 40'b0001011101101111000100101010000110011110;
                o_a2 <= 40'b0000001111110011001110111111010111001000;
                o_a3 <= 40'b0000000010101010011101010111001011010000;
                end
            7'h35 	:	 begin 
                o_a1 <= 40'b0001011100111000101011110010000101101000;
                o_a2 <= 40'b0000010000001001110001011010110111110000;
                o_a3 <= 40'b0000000010110011110001011000001010110101;
                end
            7'h36 	:	 begin 
                o_a1 <= 40'b0001011100000001110111111001110110000000;
                o_a2 <= 40'b0000010000100000010101100101010111000010;
                o_a3 <= 40'b0000000010111101011100111011011011111010;
                end
            7'h37 	:	 begin 
                o_a1 <= 40'b0001011011001010101001010011110011011000;
                o_a2 <= 40'b0000010000110110111011000000101011111000;
                o_a3 <= 40'b0000000011000111100000101010110100110110;
                end
            7'h38 	:	 begin 
                o_a1 <= 40'b0001011010010011000000010011000000011001;
                o_a2 <= 40'b0000010001001101100001001101111101010010;
                o_a3 <= 40'b0000000011010001111101010001000101000000;
                end
            7'h39 	:	 begin 
                o_a1 <= 40'b0001011001011010111101001011000101010110;
                o_a2 <= 40'b0000010001100100000111101101100010001001;
                o_a3 <= 40'b0000000011011100110011011001110110010101;
                end
            7'h3a 	:	 begin 
                o_a1 <= 40'b0001011000100010100000010000001110110001;
                o_a2 <= 40'b0000010001111010101101111111000001000101;
                o_a3 <= 40'b0000000011101000000011110001101111000010;
                end
            7'h3b 	:	 begin 
                o_a1 <= 40'b0001010111101001101001110111001011111101;
                o_a2 <= 40'b0000010010010001010011100001010000010011;
                o_a3 <= 40'b0000000011110011101111000110010011011011;
                end
            7'h3c 	:	 begin 
                o_a1 <= 40'b0001010110110000011010010101001101011001;
                o_a2 <= 40'b0000010010100111110111110010010101010110;
                o_a3 <= 40'b0000000011111111110110000110000111111010;
                end
            7'h3d 	:	 begin 
                o_a1 <= 40'b0001010101110110110010000000000011000001;
                o_a2 <= 40'b0000010010111110011010001111100100111011;
                o_a3 <= 40'b0000000100001100011001100000110011001000;
                end
            7'h3e 	:	 begin 
                o_a1 <= 40'b0001010100111100110001001101111010100011;
                o_a2 <= 40'b0000010011010100111010010101100010100100;
                o_a3 <= 40'b0000000100011001011010000111000000010100;
                end
            7'h3f 	:	 begin 
                o_a1 <= 40'b0001010100000010011000010101011101100000;
                o_a2 <= 40'b0000010011101011010111100000000000010101;
                o_a3 <= 40'b0000000100100110111000101010100001110011;
                end
            7'h40 	:	 begin 
                o_a1 <= 40'b0001010011000111100111101101101111010100;
                o_a2 <= 40'b0000010100000001110001001001111110011100;
                o_a3 <= 40'b0000000100110100110101111110010011110010;
                end
            7'h41 	:	 begin 
                o_a1 <= 40'b0001010010001100011111101110001011001110;
                o_a2 <= 40'b0000010100011000000110101101101010101111;
                o_a3 <= 40'b0000000101000011010010110110011111010001;
                end
            7'h42 	:	 begin 
                o_a1 <= 40'b0001010001010001000000101110100010001000;
                o_a2 <= 40'b0000010100101110010111100100100000010000;
                o_a3 <= 40'b0000000101010010010000001000011101010101;
                end
            7'h43 	:	 begin 
                o_a1 <= 40'b0001010000010101001011000110111000010011;
                o_a2 <= 40'b0000010101000100100011000111000110100001;
                o_a3 <= 40'b0000000101100001101110101010111010101001;
                end
            7'h44 	:	 begin 
                o_a1 <= 40'b0001001111011000111111001111100011001001;
                o_a2 <= 40'b0000010101011010101000101101010000110101;
                o_a3 <= 40'b0000000101110001101111010101111011001011;
                end
            7'h45 	:	 begin 
                o_a1 <= 40'b0001001110011100011101100001000110101010;
                o_a2 <= 40'b0000010101110000100111101101111101011011;
                o_a3 <= 40'b0000000110000010010011000010111110011110;
                end
            7'h46 	:	 begin 
                o_a1 <= 40'b0001001101011111100110010100010010111111;
                o_a2 <= 40'b0000010110000110011111011111010100011111;
                o_a3 <= 40'b0000000110010011011010101101000100000001;
                end
            7'h47 	:	 begin 
                o_a1 <= 40'b0001001100100010011010000010000001110001;
                o_a2 <= 40'b0000010110011100001111010110100111000011;
                o_a3 <= 40'b0000000110100101000111010000110000000110;
                end
            7'h48 	:	 begin 
                o_a1 <= 40'b0001001011100100111001000011010011100001;
                o_a2 <= 40'b0000010110110001110110101000001101101001;
                o_a3 <= 40'b0000000110110111011001101100010001001010;
                end
            7'h49 	:	 begin 
                o_a1 <= 40'b0001001010100111000011110001001100110100;
                o_a2 <= 40'b0000010111000111010100100111100110110111;
                o_a3 <= 40'b0000000111001010010010111111100101011100;
                end
            7'h4a 	:	 begin 
                o_a1 <= 40'b0001001001101000111010100100110011100001;
                o_a2 <= 40'b0000010111011100101000100111010101101001;
                o_a3 <= 40'b0000000111011101110100001100100001001011;
                end
            7'h4b 	:	 begin 
                o_a1 <= 40'b0001001000101010011101110111001011110110;
                o_a2 <= 40'b0000010111110001110001111000111111010111;
                o_a3 <= 40'b0000000111110001111110010110110101011001;
                end
            7'h4c 	:	 begin 
                o_a1 <= 40'b0001000111101011101110000001010101011010;
                o_a2 <= 40'b0000011000000110101111101101001001101101;
                o_a3 <= 40'b0000001000000110110010100100010111001011;
                end
            7'h4d 	:	 begin 
                o_a1 <= 40'b0001000110101100101011011100001000001101;
                o_a2 <= 40'b0000011000011011100001010011011000001000;
                o_a3 <= 40'b0000001000011100010001111101000111100010;
                end
            7'h4e 	:	 begin 
                o_a1 <= 40'b0001000101101101010110100000010001100010;
                o_a2 <= 40'b0000011000110000000101111010001001001100;
                o_a3 <= 40'b0000001000110010011101101011011100000100;
                end
            7'h4f 	:	 begin 
                o_a1 <= 40'b0001000100101101101111100110010000111010;
                o_a2 <= 40'b0000011001000100011100101110110011011001;
                o_a3 <= 40'b0000001001001001010110111100001000010010;
                end
            7'h50 	:	 begin 
                o_a1 <= 40'b0001000011101101110111000110010100110111;
                o_a2 <= 40'b0000011001011000100100111101100001101111;
                o_a3 <= 40'b0000001001100000111110111110100111101001;
                end
            7'h51 	:	 begin 
                o_a1 <= 40'b0001000010101101101101011000010111110001;
                o_a2 <= 40'b0000011001101100011101110001001111110011;
                o_a3 <= 40'b0000001001111001010111000101001000100111;
                end
            7'h52 	:	 begin 
                o_a1 <= 40'b0001000001101101010010110011111100101010;
                o_a2 <= 40'b0000011010000000000110010011100101011001;
                o_a3 <= 40'b0000001010010010100000100100111000100001;
                end
            7'h53 	:	 begin 
                o_a1 <= 40'b0001000000101100100111110000001011111111;
                o_a2 <= 40'b0000011010010011011101101100110001101110;
                o_a3 <= 40'b0000001010101100011100110110010000100011;
                end
            7'h54 	:	 begin 
                o_a1 <= 40'b0000111111101011101100100011110000010111;
                o_a2 <= 40'b0000011010100110100011000011100101111101;
                o_a3 <= 40'b0000001011000111001101010101000011101101;
                end
            7'h55 	:	 begin 
                o_a1 <= 40'b0000111110101010100001100100110011011100;
                o_a2 <= 40'b0000011010111001010101011101001111001100;
                o_a3 <= 40'b0000001011100010110011100000101110001010;
                end
            7'h56 	:	 begin 
                o_a1 <= 40'b0000111101101001000111001000111010101010;
                o_a2 <= 40'b0000011011001011110011111101001111110010;
                o_a3 <= 40'b0000001011111111010000111100100101110000;
                end
            7'h57 	:	 begin 
                o_a1 <= 40'b0000111100100111011101100101000100000100;
                o_a2 <= 40'b0000011011011101111101100101010111111011;
                o_a3 <= 40'b0000001100011100100111010000001100000101;
                end
            7'h58 	:	 begin 
                o_a1 <= 40'b0000111011100101100101001101100011010101;
                o_a2 <= 40'b0000011011101111110001010101011101010011;
                o_a3 <= 40'b0000001100111010111000000111100010000010;
                end
            7'h59 	:	 begin 
                o_a1 <= 40'b0000111010100011011110010101111110101010;
                o_a2 <= 40'b0000011100000001001110001011010010000011;
                o_a3 <= 40'b0000001101011010000101010011011101001101;
                end
            7'h5a 	:	 begin 
                o_a1 <= 40'b0000111001100001001001010001001011111010;
                o_a2 <= 40'b0000011100010010010011000010011010100000;
                o_a3 <= 40'b0000001101111010010000101001111111000011;
                end
            7'h5b 	:	 begin 
                o_a1 <= 40'b0000111000011110100110010001001101110010;
                o_a2 <= 40'b0000011100100010111110110100000001111111;
                o_a3 <= 40'b0000001110011011011100000110101110001110;
                end
            7'h5c 	:	 begin 
                o_a1 <= 40'b0000110111011011110101100111010001001101;
                o_a2 <= 40'b0000011100110011010000010110101110010101;
                o_a3 <= 40'b0000001110111101101001101011010010000111;
                end
            7'h5d 	:	 begin 
                o_a1 <= 40'b0000110110011000110111100011101010110111;
                o_a2 <= 40'b0000011101000011000110011110010010000010;
                o_a3 <= 40'b0000001111100000111011011111110001000011;
                end
            7'h5e 	:	 begin 
                o_a1 <= 40'b0000110101010101101100010101110100111111;
                o_a2 <= 40'b0000011101010010011111111011011100111110;
                o_a3 <= 40'b0000010000000101010011110011010001000100;
                end
            7'h5f 	:	 begin 
                o_a1 <= 40'b0000110100010010010100001100001101010110;
                o_a2 <= 40'b0000011101100001011011011011101011011010;
                o_a3 <= 40'b0000010000101010110100111100011011110011;
                end
            7'h60 	:	 begin 
                o_a1 <= 40'b0000110011001110101111010100010011101010;
                o_a2 <= 40'b0000011101101111110111101000110011001110;
                o_a3 <= 40'b0000010001010001100001011010000101111000;
                end
            7'h61 	:	 begin 
                o_a1 <= 40'b0000110010001010111101111010101000001101;
                o_a2 <= 40'b0000011101111101110011001000101110111110;
                o_a3 <= 40'b0000010001111001011011110011111001110100;
                end
            7'h62 	:	 begin 
                o_a1 <= 40'b0000110001000111000000001010101011000100;
                o_a2 <= 40'b0000011110001011001100011101000110110111;
                o_a3 <= 40'b0000010010100010100110111011000111001100;
                end
            7'h63 	:	 begin 
                o_a1 <= 40'b0000110000000010110110001110111011101110;
                o_a2 <= 40'b0000011110011000000010000010110110111100;
                o_a3 <= 40'b0000010011001101000101101011010110011000;
                end
            7'h64 	:	 begin 
                o_a1 <= 40'b0000101110111110100000010000111001010011;
                o_a2 <= 40'b0000011110100100010010010001110010101011;
                o_a3 <= 40'b0000010011111000111011001011100001010101;
                end
            7'h65 	:	 begin 
                o_a1 <= 40'b0000101101111001111110011001000011100010;
                o_a2 <= 40'b0000011110101111111011011100000101001100;
                o_a3 <= 40'b0000010100100110001010101110110010000100;
                end
            7'h66 	:	 begin 
                o_a1 <= 40'b0000101100110101010000101110111100100001;
                o_a2 <= 40'b0000011110111010111011101101101101111111;
                o_a3 <= 40'b0000010101010100110111110101100111100000;
                end
            7'h67 	:	 begin 
                o_a1 <= 40'b0000101011110000010111011001001011011010;
                o_a2 <= 40'b0000011111000101010001001011111001101000;
                o_a3 <= 40'b0000010110000101000110001111000001010011;
                end
            7'h68 	:	 begin 
                o_a1 <= 40'b0000101010101011010010011101100000010001;
                o_a2 <= 40'b0000011111001110111001110100010110000000;
                o_a3 <= 40'b0000010110110110111001111001110011101100;
                end
            7'h69 	:	 begin 
                o_a1 <= 40'b0000101001100110000010000000111001001101;
                o_a2 <= 40'b0000011111010111110011011100100001010100;
                o_a3 <= 40'b0000010111101010010111000110000100001001;
                end
            7'h6a 	:	 begin 
                o_a1 <= 40'b0000101000100000100110000111101001000001;
                o_a2 <= 40'b0000011111011111111011110000110011011110;
                o_a3 <= 40'b0000011000011111100010010110110000000010;
                end
            7'h6b 	:	 begin 
                o_a1 <= 40'b0000100111011010111110110101011111101110;
                o_a2 <= 40'b0000011111100111010000010011100000110111;
                o_a3 <= 40'b0000011001010110100000100011011110100011;
                end
            7'h6c 	:	 begin 
                o_a1 <= 40'b0000100110010101001100001101110101000110;
                o_a2 <= 40'b0000011111101101101110011011110101110011;
                o_a3 <= 40'b0000011010001111010110111010011111010011;
                end
            7'h6d 	:	 begin 
                o_a1 <= 40'b0000100101001111001110010011110101110010;
                o_a2 <= 40'b0000011111110011010011010100101001011101;
                o_a3 <= 40'b0000011011001010001011000010110111010010;
                end
            7'h6e 	:	 begin 
                o_a1 <= 40'b0000100100001001000101001010110011010100;
                o_a2 <= 40'b0000011111110111111011111011000111001111;
                o_a3 <= 40'b0000011100000111000010111110111110001100;
                end
            7'h6f 	:	 begin 
                o_a1 <= 40'b0000100011000010110000110110010111100010;
                o_a2 <= 40'b0000011111111011100100111101001101001011;
                o_a3 <= 40'b0000011101000110000101001111001110000110;
                end
            7'h70 	:	 begin 
                o_a1 <= 40'b0000100001111100010001011010111100001111;
                o_a2 <= 40'b0000011111111110001010110111111101101101;
                o_a3 <= 40'b0000011110000111011000110101001000010110;
                end
            7'h71 	:	 begin 
                o_a1 <= 40'b0000100000110101100110111110000111011111;
                o_a2 <= 40'b0000011111111111101001110101100011000000;
                o_a3 <= 40'b0000011111001011000101010110110010011111;
                end
            7'h72 	:	 begin 
                o_a1 <= 40'b0000011111101110110001100111001101110111;
                o_a2 <= 40'b0000011111111111111101101011000001101010;
                o_a3 <= 40'b0000100000010001010011000010101110110011;
                end
            7'h73 	:	 begin 
                o_a1 <= 40'b0000011110100111110001011111111011011101;
                o_a2 <= 40'b0000011111111111000001110101111000000100;
                o_a3 <= 40'b0000100001011010001010110100010100011001;
                end
            7'h74 	:	 begin 
                o_a1 <= 40'b0000011101100000100110110101000100111101;
                o_a2 <= 40'b0000011111111100110001011001000111100100;
                o_a3 <= 40'b0000100010100101110110011000101011111000;
                end
            7'h75 	:	 begin 
                o_a1 <= 40'b0000011100011001010001110111100010101011;
                o_a2 <= 40'b0000011111111001000110111010000011101001;
                o_a3 <= 40'b0000100011110100100000010100010110000001;
                end
            7'h76 	:	 begin 
                o_a1 <= 40'b0000011011010001110010111101010111000001;
                o_a2 <= 40'b0000011111110011111100011100100010111100;
                o_a3 <= 40'b0000100101000110010100001001100011000100;
                end
            7'h77 	:	 begin 
                o_a1 <= 40'b0000011010001010001010100011000011001010;
                o_a2 <= 40'b0000011111101101001011011110101100111101;
                o_a3 <= 40'b0000100110011011011110011111100010111001;
                end
            7'h78 	:	 begin 
                o_a1 <= 40'b0000011001000010011001001101001100100001;
                o_a2 <= 40'b0000011111100100101100110011111110010111;
                o_a3 <= 40'b0000100111110100001101001010110110101111;
                end
            7'h79 	:	 begin 
                o_a1 <= 40'b0000010111111010011111101010010110101010;
                o_a2 <= 40'b0000011111011010011000011111011100011111;
                o_a3 <= 40'b0000101001010000101111010110110000010110;
                end
            7'h7a 	:	 begin 
                o_a1 <= 40'b0000010110110010011110110101010101110111;
                o_a2 <= 40'b0000011111001110000101101101001111011000;
                o_a3 <= 40'b0000101010110001010101110000001011010110;
                end
            7'h7b 	:	 begin 
                o_a1 <= 40'b0000010101101010010111110111111111110111;
                o_a2 <= 40'b0000011110111111101010101010110111011100;
                o_a3 <= 40'b0000101100010110010010110010010001001111;
                end
            7'h7c 	:	 begin 
                o_a1 <= 40'b0000010100100010001100001110100001001000;
                o_a2 <= 40'b0000011110101110111100011110010001110111;
                o_a3 <= 40'b0000101101111111111010110100111011001000;
                end
            7'h7d 	:	 begin 
                o_a1 <= 40'b0000010011011001111101101011011111000001;
                o_a2 <= 40'b0000011110011011101110111011011100000100;
                o_a3 <= 40'b0000101111101110100100011101101000110101;
                end
            7'h7e 	:	 begin 
                o_a1 <= 40'b0000010010010001101110011100110001001000;
                o_a2 <= 40'b0000011110000101110100011000000010011100;
                o_a3 <= 40'b0000110001100010101000110011001001111110;
                end
            7'h7f 	:	 begin 
                o_a1 <= 40'b0000010001001001100001010001011110100111;
                o_a2 <= 40'b0000011101101100111101011101000010110000;
                o_a3 <= 40'b0000110011011100100011110100011011110111;
                end
        endcase
	end								
endmodule
