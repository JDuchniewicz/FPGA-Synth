module quarter_sine_lut(input[8:0] i_phase,
								output reg signed[15:0] o_val);
        initial o_val = 16'b0;

		always @(i_phase) begin
			case(i_phase)
                9'h000 	:	o_val <= 16'b0000000000110010;
                9'h001 	:	o_val <= 16'b0000000010010110;
                9'h002 	:	o_val <= 16'b0000000011111011;
                9'h003 	:	o_val <= 16'b0000000101011111;
                9'h004 	:	o_val <= 16'b0000000111000100;
                9'h005 	:	o_val <= 16'b0000001000101000;
                9'h006 	:	o_val <= 16'b0000001010001101;
                9'h007 	:	o_val <= 16'b0000001011110001;
                9'h008 	:	o_val <= 16'b0000001101010110;
                9'h009 	:	o_val <= 16'b0000001110111010;
                9'h00a 	:	o_val <= 16'b0000010000011111;
                9'h00b 	:	o_val <= 16'b0000010010000011;
                9'h00c 	:	o_val <= 16'b0000010011101000;
                9'h00d 	:	o_val <= 16'b0000010101001100;
                9'h00e 	:	o_val <= 16'b0000010110110001;
                9'h00f 	:	o_val <= 16'b0000011000010101;
                9'h010 	:	o_val <= 16'b0000011001111010;
                9'h011 	:	o_val <= 16'b0000011011011110;
                9'h012 	:	o_val <= 16'b0000011101000010;
                9'h013 	:	o_val <= 16'b0000011110100111;
                9'h014 	:	o_val <= 16'b0000100000001011;
                9'h015 	:	o_val <= 16'b0000100001101111;
                9'h016 	:	o_val <= 16'b0000100011010100;
                9'h017 	:	o_val <= 16'b0000100100111000;
                9'h018 	:	o_val <= 16'b0000100110011100;
                9'h019 	:	o_val <= 16'b0000101000000000;
                9'h01a 	:	o_val <= 16'b0000101001100101;
                9'h01b 	:	o_val <= 16'b0000101011001001;
                9'h01c 	:	o_val <= 16'b0000101100101101;
                9'h01d 	:	o_val <= 16'b0000101110010001;
                9'h01e 	:	o_val <= 16'b0000101111110101;
                9'h01f 	:	o_val <= 16'b0000110001011001;
                9'h020 	:	o_val <= 16'b0000110010111101;
                9'h021 	:	o_val <= 16'b0000110100100001;
                9'h022 	:	o_val <= 16'b0000110110000101;
                9'h023 	:	o_val <= 16'b0000110111101001;
                9'h024 	:	o_val <= 16'b0000111001001101;
                9'h025 	:	o_val <= 16'b0000111010110001;
                9'h026 	:	o_val <= 16'b0000111100010101;
                9'h027 	:	o_val <= 16'b0000111101111001;
                9'h028 	:	o_val <= 16'b0000111111011101;
                9'h029 	:	o_val <= 16'b0001000001000000;
                9'h02a 	:	o_val <= 16'b0001000010100100;
                9'h02b 	:	o_val <= 16'b0001000100001000;
                9'h02c 	:	o_val <= 16'b0001000101101011;
                9'h02d 	:	o_val <= 16'b0001000111001111;
                9'h02e 	:	o_val <= 16'b0001001000110010;
                9'h02f 	:	o_val <= 16'b0001001010010110;
                9'h030 	:	o_val <= 16'b0001001011111001;
                9'h031 	:	o_val <= 16'b0001001101011101;
                9'h032 	:	o_val <= 16'b0001001111000000;
                9'h033 	:	o_val <= 16'b0001010000100011;
                9'h034 	:	o_val <= 16'b0001010010000111;
                9'h035 	:	o_val <= 16'b0001010011101010;
                9'h036 	:	o_val <= 16'b0001010101001101;
                9'h037 	:	o_val <= 16'b0001010110110000;
                9'h038 	:	o_val <= 16'b0001011000010011;
                9'h039 	:	o_val <= 16'b0001011001110110;
                9'h03a 	:	o_val <= 16'b0001011011011001;
                9'h03b 	:	o_val <= 16'b0001011100111100;
                9'h03c 	:	o_val <= 16'b0001011110011111;
                9'h03d 	:	o_val <= 16'b0001100000000010;
                9'h03e 	:	o_val <= 16'b0001100001100100;
                9'h03f 	:	o_val <= 16'b0001100011000111;
                9'h040 	:	o_val <= 16'b0001100100101010;
                9'h041 	:	o_val <= 16'b0001100110001100;
                9'h042 	:	o_val <= 16'b0001100111101111;
                9'h043 	:	o_val <= 16'b0001101001010001;
                9'h044 	:	o_val <= 16'b0001101010110011;
                9'h045 	:	o_val <= 16'b0001101100010110;
                9'h046 	:	o_val <= 16'b0001101101111000;
                9'h047 	:	o_val <= 16'b0001101111011010;
                9'h048 	:	o_val <= 16'b0001110000111100;
                9'h049 	:	o_val <= 16'b0001110010011110;
                9'h04a 	:	o_val <= 16'b0001110100000000;
                9'h04b 	:	o_val <= 16'b0001110101100010;
                9'h04c 	:	o_val <= 16'b0001110111000100;
                9'h04d 	:	o_val <= 16'b0001111000100101;
                9'h04e 	:	o_val <= 16'b0001111010000111;
                9'h04f 	:	o_val <= 16'b0001111011101001;
                9'h050 	:	o_val <= 16'b0001111101001010;
                9'h051 	:	o_val <= 16'b0001111110101100;
                9'h052 	:	o_val <= 16'b0010000000001101;
                9'h053 	:	o_val <= 16'b0010000001101110;
                9'h054 	:	o_val <= 16'b0010000011010000;
                9'h055 	:	o_val <= 16'b0010000100110001;
                9'h056 	:	o_val <= 16'b0010000110010010;
                9'h057 	:	o_val <= 16'b0010000111110011;
                9'h058 	:	o_val <= 16'b0010001001010100;
                9'h059 	:	o_val <= 16'b0010001010110100;
                9'h05a 	:	o_val <= 16'b0010001100010101;
                9'h05b 	:	o_val <= 16'b0010001101110110;
                9'h05c 	:	o_val <= 16'b0010001111010110;
                9'h05d 	:	o_val <= 16'b0010010000110111;
                9'h05e 	:	o_val <= 16'b0010010010010111;
                9'h05f 	:	o_val <= 16'b0010010011110111;
                9'h060 	:	o_val <= 16'b0010010101011000;
                9'h061 	:	o_val <= 16'b0010010110111000;
                9'h062 	:	o_val <= 16'b0010011000011000;
                9'h063 	:	o_val <= 16'b0010011001111000;
                9'h064 	:	o_val <= 16'b0010011011011000;
                9'h065 	:	o_val <= 16'b0010011100110111;
                9'h066 	:	o_val <= 16'b0010011110010111;
                9'h067 	:	o_val <= 16'b0010011111110110;
                9'h068 	:	o_val <= 16'b0010100001010110;
                9'h069 	:	o_val <= 16'b0010100010110101;
                9'h06a 	:	o_val <= 16'b0010100100010101;
                9'h06b 	:	o_val <= 16'b0010100101110100;
                9'h06c 	:	o_val <= 16'b0010100111010011;
                9'h06d 	:	o_val <= 16'b0010101000110010;
                9'h06e 	:	o_val <= 16'b0010101010010001;
                9'h06f 	:	o_val <= 16'b0010101011101111;
                9'h070 	:	o_val <= 16'b0010101101001110;
                9'h071 	:	o_val <= 16'b0010101110101101;
                9'h072 	:	o_val <= 16'b0010110000001011;
                9'h073 	:	o_val <= 16'b0010110001101001;
                9'h074 	:	o_val <= 16'b0010110011001000;
                9'h075 	:	o_val <= 16'b0010110100100110;
                9'h076 	:	o_val <= 16'b0010110110000100;
                9'h077 	:	o_val <= 16'b0010110111100010;
                9'h078 	:	o_val <= 16'b0010111000111111;
                9'h079 	:	o_val <= 16'b0010111010011101;
                9'h07a 	:	o_val <= 16'b0010111011111011;
                9'h07b 	:	o_val <= 16'b0010111101011000;
                9'h07c 	:	o_val <= 16'b0010111110110101;
                9'h07d 	:	o_val <= 16'b0011000000010011;
                9'h07e 	:	o_val <= 16'b0011000001110000;
                9'h07f 	:	o_val <= 16'b0011000011001101;
                9'h080 	:	o_val <= 16'b0011000100101010;
                9'h081 	:	o_val <= 16'b0011000110000110;
                9'h082 	:	o_val <= 16'b0011000111100011;
                9'h083 	:	o_val <= 16'b0011001001000000;
                9'h084 	:	o_val <= 16'b0011001010011100;
                9'h085 	:	o_val <= 16'b0011001011111000;
                9'h086 	:	o_val <= 16'b0011001101010100;
                9'h087 	:	o_val <= 16'b0011001110110000;
                9'h088 	:	o_val <= 16'b0011010000001100;
                9'h089 	:	o_val <= 16'b0011010001101000;
                9'h08a 	:	o_val <= 16'b0011010011000100;
                9'h08b 	:	o_val <= 16'b0011010100011111;
                9'h08c 	:	o_val <= 16'b0011010101111011;
                9'h08d 	:	o_val <= 16'b0011010111010110;
                9'h08e 	:	o_val <= 16'b0011011000110001;
                9'h08f 	:	o_val <= 16'b0011011010001100;
                9'h090 	:	o_val <= 16'b0011011011100111;
                9'h091 	:	o_val <= 16'b0011011101000010;
                9'h092 	:	o_val <= 16'b0011011110011100;
                9'h093 	:	o_val <= 16'b0011011111110111;
                9'h094 	:	o_val <= 16'b0011100001010001;
                9'h095 	:	o_val <= 16'b0011100010101011;
                9'h096 	:	o_val <= 16'b0011100100000110;
                9'h097 	:	o_val <= 16'b0011100101011111;
                9'h098 	:	o_val <= 16'b0011100110111001;
                9'h099 	:	o_val <= 16'b0011101000010011;
                9'h09a 	:	o_val <= 16'b0011101001101100;
                9'h09b 	:	o_val <= 16'b0011101011000110;
                9'h09c 	:	o_val <= 16'b0011101100011111;
                9'h09d 	:	o_val <= 16'b0011101101111000;
                9'h09e 	:	o_val <= 16'b0011101111010001;
                9'h09f 	:	o_val <= 16'b0011110000101010;
                9'h0a0 	:	o_val <= 16'b0011110010000011;
                9'h0a1 	:	o_val <= 16'b0011110011011011;
                9'h0a2 	:	o_val <= 16'b0011110100110011;
                9'h0a3 	:	o_val <= 16'b0011110110001100;
                9'h0a4 	:	o_val <= 16'b0011110111100100;
                9'h0a5 	:	o_val <= 16'b0011111000111100;
                9'h0a6 	:	o_val <= 16'b0011111010010011;
                9'h0a7 	:	o_val <= 16'b0011111011101011;
                9'h0a8 	:	o_val <= 16'b0011111101000011;
                9'h0a9 	:	o_val <= 16'b0011111110011010;
                9'h0aa 	:	o_val <= 16'b0011111111110001;
                9'h0ab 	:	o_val <= 16'b0100000001001000;
                9'h0ac 	:	o_val <= 16'b0100000010011111;
                9'h0ad 	:	o_val <= 16'b0100000011110110;
                9'h0ae 	:	o_val <= 16'b0100000101001100;
                9'h0af 	:	o_val <= 16'b0100000110100010;
                9'h0b0 	:	o_val <= 16'b0100000111111001;
                9'h0b1 	:	o_val <= 16'b0100001001001111;
                9'h0b2 	:	o_val <= 16'b0100001010100101;
                9'h0b3 	:	o_val <= 16'b0100001011111010;
                9'h0b4 	:	o_val <= 16'b0100001101010000;
                9'h0b5 	:	o_val <= 16'b0100001110100101;
                9'h0b6 	:	o_val <= 16'b0100001111111011;
                9'h0b7 	:	o_val <= 16'b0100010001010000;
                9'h0b8 	:	o_val <= 16'b0100010010100101;
                9'h0b9 	:	o_val <= 16'b0100010011111010;
                9'h0ba 	:	o_val <= 16'b0100010101001110;
                9'h0bb 	:	o_val <= 16'b0100010110100011;
                9'h0bc 	:	o_val <= 16'b0100010111110111;
                9'h0bd 	:	o_val <= 16'b0100011001001011;
                9'h0be 	:	o_val <= 16'b0100011010011111;
                9'h0bf 	:	o_val <= 16'b0100011011110011;
                9'h0c0 	:	o_val <= 16'b0100011101000110;
                9'h0c1 	:	o_val <= 16'b0100011110011010;
                9'h0c2 	:	o_val <= 16'b0100011111101101;
                9'h0c3 	:	o_val <= 16'b0100100001000000;
                9'h0c4 	:	o_val <= 16'b0100100010010011;
                9'h0c5 	:	o_val <= 16'b0100100011100110;
                9'h0c6 	:	o_val <= 16'b0100100100111000;
                9'h0c7 	:	o_val <= 16'b0100100110001010;
                9'h0c8 	:	o_val <= 16'b0100100111011101;
                9'h0c9 	:	o_val <= 16'b0100101000101111;
                9'h0ca 	:	o_val <= 16'b0100101010000001;
                9'h0cb 	:	o_val <= 16'b0100101011010010;
                9'h0cc 	:	o_val <= 16'b0100101100100100;
                9'h0cd 	:	o_val <= 16'b0100101101110101;
                9'h0ce 	:	o_val <= 16'b0100101111000110;
                9'h0cf 	:	o_val <= 16'b0100110000010111;
                9'h0d0 	:	o_val <= 16'b0100110001101000;
                9'h0d1 	:	o_val <= 16'b0100110010111000;
                9'h0d2 	:	o_val <= 16'b0100110100001001;
                9'h0d3 	:	o_val <= 16'b0100110101011001;
                9'h0d4 	:	o_val <= 16'b0100110110101001;
                9'h0d5 	:	o_val <= 16'b0100110111111001;
                9'h0d6 	:	o_val <= 16'b0100111001001000;
                9'h0d7 	:	o_val <= 16'b0100111010011000;
                9'h0d8 	:	o_val <= 16'b0100111011100111;
                9'h0d9 	:	o_val <= 16'b0100111100110110;
                9'h0da 	:	o_val <= 16'b0100111110000101;
                9'h0db 	:	o_val <= 16'b0100111111010100;
                9'h0dc 	:	o_val <= 16'b0101000000100010;
                9'h0dd 	:	o_val <= 16'b0101000001110000;
                9'h0de 	:	o_val <= 16'b0101000010111111;
                9'h0df 	:	o_val <= 16'b0101000100001100;
                9'h0e0 	:	o_val <= 16'b0101000101011010;
                9'h0e1 	:	o_val <= 16'b0101000110101000;
                9'h0e2 	:	o_val <= 16'b0101000111110101;
                9'h0e3 	:	o_val <= 16'b0101001001000010;
                9'h0e4 	:	o_val <= 16'b0101001010001111;
                9'h0e5 	:	o_val <= 16'b0101001011011100;
                9'h0e6 	:	o_val <= 16'b0101001100101000;
                9'h0e7 	:	o_val <= 16'b0101001101110101;
                9'h0e8 	:	o_val <= 16'b0101001111000001;
                9'h0e9 	:	o_val <= 16'b0101010000001101;
                9'h0ea 	:	o_val <= 16'b0101010001011000;
                9'h0eb 	:	o_val <= 16'b0101010010100100;
                9'h0ec 	:	o_val <= 16'b0101010011101111;
                9'h0ed 	:	o_val <= 16'b0101010100111010;
                9'h0ee 	:	o_val <= 16'b0101010110000101;
                9'h0ef 	:	o_val <= 16'b0101010111010000;
                9'h0f0 	:	o_val <= 16'b0101011000011010;
                9'h0f1 	:	o_val <= 16'b0101011001100101;
                9'h0f2 	:	o_val <= 16'b0101011010101111;
                9'h0f3 	:	o_val <= 16'b0101011011111001;
                9'h0f4 	:	o_val <= 16'b0101011101000010;
                9'h0f5 	:	o_val <= 16'b0101011110001100;
                9'h0f6 	:	o_val <= 16'b0101011111010101;
                9'h0f7 	:	o_val <= 16'b0101100000011110;
                9'h0f8 	:	o_val <= 16'b0101100001100111;
                9'h0f9 	:	o_val <= 16'b0101100010101111;
                9'h0fa 	:	o_val <= 16'b0101100011111000;
                9'h0fb 	:	o_val <= 16'b0101100101000000;
                9'h0fc 	:	o_val <= 16'b0101100110001000;
                9'h0fd 	:	o_val <= 16'b0101100111010000;
                9'h0fe 	:	o_val <= 16'b0101101000010111;
                9'h0ff 	:	o_val <= 16'b0101101001011110;
                9'h100 	:	o_val <= 16'b0101101010100101;
                9'h101 	:	o_val <= 16'b0101101011101100;
                9'h102 	:	o_val <= 16'b0101101100110011;
                9'h103 	:	o_val <= 16'b0101101101111001;
                9'h104 	:	o_val <= 16'b0101101111000000;
                9'h105 	:	o_val <= 16'b0101110000000110;
                9'h106 	:	o_val <= 16'b0101110001001011;
                9'h107 	:	o_val <= 16'b0101110010010001;
                9'h108 	:	o_val <= 16'b0101110011010110;
                9'h109 	:	o_val <= 16'b0101110100011011;
                9'h10a 	:	o_val <= 16'b0101110101100000;
                9'h10b 	:	o_val <= 16'b0101110110100101;
                9'h10c 	:	o_val <= 16'b0101110111101001;
                9'h10d 	:	o_val <= 16'b0101111000101101;
                9'h10e 	:	o_val <= 16'b0101111001110001;
                9'h10f 	:	o_val <= 16'b0101111010110101;
                9'h110 	:	o_val <= 16'b0101111011111001;
                9'h111 	:	o_val <= 16'b0101111100111100;
                9'h112 	:	o_val <= 16'b0101111101111111;
                9'h113 	:	o_val <= 16'b0101111111000010;
                9'h114 	:	o_val <= 16'b0110000000000100;
                9'h115 	:	o_val <= 16'b0110000001000111;
                9'h116 	:	o_val <= 16'b0110000010001001;
                9'h117 	:	o_val <= 16'b0110000011001011;
                9'h118 	:	o_val <= 16'b0110000100001101;
                9'h119 	:	o_val <= 16'b0110000101001110;
                9'h11a 	:	o_val <= 16'b0110000110001111;
                9'h11b 	:	o_val <= 16'b0110000111010000;
                9'h11c 	:	o_val <= 16'b0110001000010001;
                9'h11d 	:	o_val <= 16'b0110001001010001;
                9'h11e 	:	o_val <= 16'b0110001010010010;
                9'h11f 	:	o_val <= 16'b0110001011010010;
                9'h120 	:	o_val <= 16'b0110001100010001;
                9'h121 	:	o_val <= 16'b0110001101010001;
                9'h122 	:	o_val <= 16'b0110001110010000;
                9'h123 	:	o_val <= 16'b0110001111001111;
                9'h124 	:	o_val <= 16'b0110010000001110;
                9'h125 	:	o_val <= 16'b0110010001001101;
                9'h126 	:	o_val <= 16'b0110010010001011;
                9'h127 	:	o_val <= 16'b0110010011001001;
                9'h128 	:	o_val <= 16'b0110010100000111;
                9'h129 	:	o_val <= 16'b0110010101000101;
                9'h12a 	:	o_val <= 16'b0110010110000010;
                9'h12b 	:	o_val <= 16'b0110010110111111;
                9'h12c 	:	o_val <= 16'b0110010111111100;
                9'h12d 	:	o_val <= 16'b0110011000111001;
                9'h12e 	:	o_val <= 16'b0110011001110101;
                9'h12f 	:	o_val <= 16'b0110011010110001;
                9'h130 	:	o_val <= 16'b0110011011101101;
                9'h131 	:	o_val <= 16'b0110011100101001;
                9'h132 	:	o_val <= 16'b0110011101100100;
                9'h133 	:	o_val <= 16'b0110011110011111;
                9'h134 	:	o_val <= 16'b0110011111011010;
                9'h135 	:	o_val <= 16'b0110100000010101;
                9'h136 	:	o_val <= 16'b0110100001001111;
                9'h137 	:	o_val <= 16'b0110100010001001;
                9'h138 	:	o_val <= 16'b0110100011000011;
                9'h139 	:	o_val <= 16'b0110100011111101;
                9'h13a 	:	o_val <= 16'b0110100100110110;
                9'h13b 	:	o_val <= 16'b0110100101101111;
                9'h13c 	:	o_val <= 16'b0110100110101000;
                9'h13d 	:	o_val <= 16'b0110100111100001;
                9'h13e 	:	o_val <= 16'b0110101000011001;
                9'h13f 	:	o_val <= 16'b0110101001010001;
                9'h140 	:	o_val <= 16'b0110101010001001;
                9'h141 	:	o_val <= 16'b0110101011000001;
                9'h142 	:	o_val <= 16'b0110101011111000;
                9'h143 	:	o_val <= 16'b0110101100101111;
                9'h144 	:	o_val <= 16'b0110101101100110;
                9'h145 	:	o_val <= 16'b0110101110011100;
                9'h146 	:	o_val <= 16'b0110101111010011;
                9'h147 	:	o_val <= 16'b0110110000001001;
                9'h148 	:	o_val <= 16'b0110110000111111;
                9'h149 	:	o_val <= 16'b0110110001110100;
                9'h14a 	:	o_val <= 16'b0110110010101001;
                9'h14b 	:	o_val <= 16'b0110110011011110;
                9'h14c 	:	o_val <= 16'b0110110100010011;
                9'h14d 	:	o_val <= 16'b0110110101001000;
                9'h14e 	:	o_val <= 16'b0110110101111100;
                9'h14f 	:	o_val <= 16'b0110110110110000;
                9'h150 	:	o_val <= 16'b0110110111100011;
                9'h151 	:	o_val <= 16'b0110111000010111;
                9'h152 	:	o_val <= 16'b0110111001001010;
                9'h153 	:	o_val <= 16'b0110111001111101;
                9'h154 	:	o_val <= 16'b0110111010101111;
                9'h155 	:	o_val <= 16'b0110111011100010;
                9'h156 	:	o_val <= 16'b0110111100010100;
                9'h157 	:	o_val <= 16'b0110111101000110;
                9'h158 	:	o_val <= 16'b0110111101110111;
                9'h159 	:	o_val <= 16'b0110111110101001;
                9'h15a 	:	o_val <= 16'b0110111111011010;
                9'h15b 	:	o_val <= 16'b0111000000001010;
                9'h15c 	:	o_val <= 16'b0111000000111011;
                9'h15d 	:	o_val <= 16'b0111000001101011;
                9'h15e 	:	o_val <= 16'b0111000010011011;
                9'h15f 	:	o_val <= 16'b0111000011001011;
                9'h160 	:	o_val <= 16'b0111000011111010;
                9'h161 	:	o_val <= 16'b0111000100101001;
                9'h162 	:	o_val <= 16'b0111000101011000;
                9'h163 	:	o_val <= 16'b0111000110000110;
                9'h164 	:	o_val <= 16'b0111000110110101;
                9'h165 	:	o_val <= 16'b0111000111100011;
                9'h166 	:	o_val <= 16'b0111001000010001;
                9'h167 	:	o_val <= 16'b0111001000111110;
                9'h168 	:	o_val <= 16'b0111001001101011;
                9'h169 	:	o_val <= 16'b0111001010011000;
                9'h16a 	:	o_val <= 16'b0111001011000101;
                9'h16b 	:	o_val <= 16'b0111001011110001;
                9'h16c 	:	o_val <= 16'b0111001100011101;
                9'h16d 	:	o_val <= 16'b0111001101001001;
                9'h16e 	:	o_val <= 16'b0111001101110101;
                9'h16f 	:	o_val <= 16'b0111001110100000;
                9'h170 	:	o_val <= 16'b0111001111001011;
                9'h171 	:	o_val <= 16'b0111001111110110;
                9'h172 	:	o_val <= 16'b0111010000100000;
                9'h173 	:	o_val <= 16'b0111010001001010;
                9'h174 	:	o_val <= 16'b0111010001110100;
                9'h175 	:	o_val <= 16'b0111010010011110;
                9'h176 	:	o_val <= 16'b0111010011000111;
                9'h177 	:	o_val <= 16'b0111010011110000;
                9'h178 	:	o_val <= 16'b0111010100011001;
                9'h179 	:	o_val <= 16'b0111010101000001;
                9'h17a 	:	o_val <= 16'b0111010101101001;
                9'h17b 	:	o_val <= 16'b0111010110010001;
                9'h17c 	:	o_val <= 16'b0111010110111001;
                9'h17d 	:	o_val <= 16'b0111010111100000;
                9'h17e 	:	o_val <= 16'b0111011000000111;
                9'h17f 	:	o_val <= 16'b0111011000101110;
                9'h180 	:	o_val <= 16'b0111011001010100;
                9'h181 	:	o_val <= 16'b0111011001111011;
                9'h182 	:	o_val <= 16'b0111011010100000;
                9'h183 	:	o_val <= 16'b0111011011000110;
                9'h184 	:	o_val <= 16'b0111011011101011;
                9'h185 	:	o_val <= 16'b0111011100010000;
                9'h186 	:	o_val <= 16'b0111011100110101;
                9'h187 	:	o_val <= 16'b0111011101011010;
                9'h188 	:	o_val <= 16'b0111011101111110;
                9'h189 	:	o_val <= 16'b0111011110100010;
                9'h18a 	:	o_val <= 16'b0111011111000101;
                9'h18b 	:	o_val <= 16'b0111011111101001;
                9'h18c 	:	o_val <= 16'b0111100000001100;
                9'h18d 	:	o_val <= 16'b0111100000101110;
                9'h18e 	:	o_val <= 16'b0111100001010001;
                9'h18f 	:	o_val <= 16'b0111100001110011;
                9'h190 	:	o_val <= 16'b0111100010010101;
                9'h191 	:	o_val <= 16'b0111100010110110;
                9'h192 	:	o_val <= 16'b0111100011011000;
                9'h193 	:	o_val <= 16'b0111100011111001;
                9'h194 	:	o_val <= 16'b0111100100011001;
                9'h195 	:	o_val <= 16'b0111100100111010;
                9'h196 	:	o_val <= 16'b0111100101011010;
                9'h197 	:	o_val <= 16'b0111100101111010;
                9'h198 	:	o_val <= 16'b0111100110011001;
                9'h199 	:	o_val <= 16'b0111100110111001;
                9'h19a 	:	o_val <= 16'b0111100111011000;
                9'h19b 	:	o_val <= 16'b0111100111110110;
                9'h19c 	:	o_val <= 16'b0111101000010101;
                9'h19d 	:	o_val <= 16'b0111101000110011;
                9'h19e 	:	o_val <= 16'b0111101001010000;
                9'h19f 	:	o_val <= 16'b0111101001101110;
                9'h1a0 	:	o_val <= 16'b0111101010001011;
                9'h1a1 	:	o_val <= 16'b0111101010101000;
                9'h1a2 	:	o_val <= 16'b0111101011000101;
                9'h1a3 	:	o_val <= 16'b0111101011100001;
                9'h1a4 	:	o_val <= 16'b0111101011111101;
                9'h1a5 	:	o_val <= 16'b0111101100011001;
                9'h1a6 	:	o_val <= 16'b0111101100110100;
                9'h1a7 	:	o_val <= 16'b0111101101001111;
                9'h1a8 	:	o_val <= 16'b0111101101101010;
                9'h1a9 	:	o_val <= 16'b0111101110000100;
                9'h1aa 	:	o_val <= 16'b0111101110011111;
                9'h1ab 	:	o_val <= 16'b0111101110111001;
                9'h1ac 	:	o_val <= 16'b0111101111010010;
                9'h1ad 	:	o_val <= 16'b0111101111101011;
                9'h1ae 	:	o_val <= 16'b0111110000000101;
                9'h1af 	:	o_val <= 16'b0111110000011101;
                9'h1b0 	:	o_val <= 16'b0111110000110110;
                9'h1b1 	:	o_val <= 16'b0111110001001110;
                9'h1b2 	:	o_val <= 16'b0111110001100110;
                9'h1b3 	:	o_val <= 16'b0111110001111101;
                9'h1b4 	:	o_val <= 16'b0111110010010100;
                9'h1b5 	:	o_val <= 16'b0111110010101011;
                9'h1b6 	:	o_val <= 16'b0111110011000010;
                9'h1b7 	:	o_val <= 16'b0111110011011000;
                9'h1b8 	:	o_val <= 16'b0111110011101110;
                9'h1b9 	:	o_val <= 16'b0111110100000100;
                9'h1ba 	:	o_val <= 16'b0111110100011001;
                9'h1bb 	:	o_val <= 16'b0111110100101111;
                9'h1bc 	:	o_val <= 16'b0111110101000011;
                9'h1bd 	:	o_val <= 16'b0111110101011000;
                9'h1be 	:	o_val <= 16'b0111110101101100;
                9'h1bf 	:	o_val <= 16'b0111110110000000;
                9'h1c0 	:	o_val <= 16'b0111110110010100;
                9'h1c1 	:	o_val <= 16'b0111110110100111;
                9'h1c2 	:	o_val <= 16'b0111110110111010;
                9'h1c3 	:	o_val <= 16'b0111110111001101;
                9'h1c4 	:	o_val <= 16'b0111110111011111;
                9'h1c5 	:	o_val <= 16'b0111110111110001;
                9'h1c6 	:	o_val <= 16'b0111111000000011;
                9'h1c7 	:	o_val <= 16'b0111111000010100;
                9'h1c8 	:	o_val <= 16'b0111111000100110;
                9'h1c9 	:	o_val <= 16'b0111111000110111;
                9'h1ca 	:	o_val <= 16'b0111111001000111;
                9'h1cb 	:	o_val <= 16'b0111111001010111;
                9'h1cc 	:	o_val <= 16'b0111111001100111;
                9'h1cd 	:	o_val <= 16'b0111111001110111;
                9'h1ce 	:	o_val <= 16'b0111111010000110;
                9'h1cf 	:	o_val <= 16'b0111111010010101;
                9'h1d0 	:	o_val <= 16'b0111111010100100;
                9'h1d1 	:	o_val <= 16'b0111111010110011;
                9'h1d2 	:	o_val <= 16'b0111111011000001;
                9'h1d3 	:	o_val <= 16'b0111111011001111;
                9'h1d4 	:	o_val <= 16'b0111111011011100;
                9'h1d5 	:	o_val <= 16'b0111111011101001;
                9'h1d6 	:	o_val <= 16'b0111111011110110;
                9'h1d7 	:	o_val <= 16'b0111111100000011;
                9'h1d8 	:	o_val <= 16'b0111111100001111;
                9'h1d9 	:	o_val <= 16'b0111111100011011;
                9'h1da 	:	o_val <= 16'b0111111100100111;
                9'h1db 	:	o_val <= 16'b0111111100110010;
                9'h1dc 	:	o_val <= 16'b0111111100111101;
                9'h1dd 	:	o_val <= 16'b0111111101001000;
                9'h1de 	:	o_val <= 16'b0111111101010011;
                9'h1df 	:	o_val <= 16'b0111111101011101;
                9'h1e0 	:	o_val <= 16'b0111111101100111;
                9'h1e1 	:	o_val <= 16'b0111111101110000;
                9'h1e2 	:	o_val <= 16'b0111111101111001;
                9'h1e3 	:	o_val <= 16'b0111111110000010;
                9'h1e4 	:	o_val <= 16'b0111111110001011;
                9'h1e5 	:	o_val <= 16'b0111111110010011;
                9'h1e6 	:	o_val <= 16'b0111111110011011;
                9'h1e7 	:	o_val <= 16'b0111111110100011;
                9'h1e8 	:	o_val <= 16'b0111111110101010;
                9'h1e9 	:	o_val <= 16'b0111111110110001;
                9'h1ea 	:	o_val <= 16'b0111111110111000;
                9'h1eb 	:	o_val <= 16'b0111111110111111;
                9'h1ec 	:	o_val <= 16'b0111111111000101;
                9'h1ed 	:	o_val <= 16'b0111111111001011;
                9'h1ee 	:	o_val <= 16'b0111111111010000;
                9'h1ef 	:	o_val <= 16'b0111111111010110;
                9'h1f0 	:	o_val <= 16'b0111111111011010;
                9'h1f1 	:	o_val <= 16'b0111111111011111;
                9'h1f2 	:	o_val <= 16'b0111111111100011;
                9'h1f3 	:	o_val <= 16'b0111111111100111;
                9'h1f4 	:	o_val <= 16'b0111111111101011;
                9'h1f5 	:	o_val <= 16'b0111111111101110;
                9'h1f6 	:	o_val <= 16'b0111111111110010;
                9'h1f7 	:	o_val <= 16'b0111111111110100;
                9'h1f8 	:	o_val <= 16'b0111111111110111;
                9'h1f9 	:	o_val <= 16'b0111111111111001;
                9'h1fa 	:	o_val <= 16'b0111111111111011;
                9'h1fb 	:	o_val <= 16'b0111111111111100;
                9'h1fc 	:	o_val <= 16'b0111111111111110;
                9'h1fd 	:	o_val <= 16'b0111111111111111;
                9'h1fe 	:	o_val <= 16'b0111111111111111;
                9'h1ff 	:	o_val <= 16'b0111111111111111;
				 default		:	o_val <= 16'b0;
			endcase
		end
endmodule
                                        
