module quarter_sine_lut(input[13:0] i_phase,
								output reg signed[15:0] o_val);
		always @(i_phase) begin
			case(i_phase)
            14'h0000 	:	o_val <= 16'b0000000000000001;
            14'h0001 	:	o_val <= 16'b0000000000000100;
            14'h0002 	:	o_val <= 16'b0000000000000111;
            14'h0003 	:	o_val <= 16'b0000000000001010;
            14'h0004 	:	o_val <= 16'b0000000000001110;
            14'h0005 	:	o_val <= 16'b0000000000010001;
            14'h0006 	:	o_val <= 16'b0000000000010100;
            14'h0007 	:	o_val <= 16'b0000000000010111;
            14'h0008 	:	o_val <= 16'b0000000000011010;
            14'h0009 	:	o_val <= 16'b0000000000011101;
            14'h000a 	:	o_val <= 16'b0000000000100000;
            14'h000b 	:	o_val <= 16'b0000000000100100;
            14'h000c 	:	o_val <= 16'b0000000000100111;
            14'h000d 	:	o_val <= 16'b0000000000101010;
            14'h000e 	:	o_val <= 16'b0000000000101101;
            14'h000f 	:	o_val <= 16'b0000000000110000;
            14'h0010 	:	o_val <= 16'b0000000000110011;
            14'h0011 	:	o_val <= 16'b0000000000110110;
            14'h0012 	:	o_val <= 16'b0000000000111010;
            14'h0013 	:	o_val <= 16'b0000000000111101;
            14'h0014 	:	o_val <= 16'b0000000001000000;
            14'h0015 	:	o_val <= 16'b0000000001000011;
            14'h0016 	:	o_val <= 16'b0000000001000110;
            14'h0017 	:	o_val <= 16'b0000000001001001;
            14'h0018 	:	o_val <= 16'b0000000001001100;
            14'h0019 	:	o_val <= 16'b0000000001010000;
            14'h001a 	:	o_val <= 16'b0000000001010011;
            14'h001b 	:	o_val <= 16'b0000000001010110;
            14'h001c 	:	o_val <= 16'b0000000001011001;
            14'h001d 	:	o_val <= 16'b0000000001011100;
            14'h001e 	:	o_val <= 16'b0000000001011111;
            14'h001f 	:	o_val <= 16'b0000000001100010;
            14'h0020 	:	o_val <= 16'b0000000001100110;
            14'h0021 	:	o_val <= 16'b0000000001101001;
            14'h0022 	:	o_val <= 16'b0000000001101100;
            14'h0023 	:	o_val <= 16'b0000000001101111;
            14'h0024 	:	o_val <= 16'b0000000001110010;
            14'h0025 	:	o_val <= 16'b0000000001110101;
            14'h0026 	:	o_val <= 16'b0000000001111000;
            14'h0027 	:	o_val <= 16'b0000000001111100;
            14'h0028 	:	o_val <= 16'b0000000001111111;
            14'h0029 	:	o_val <= 16'b0000000010000010;
            14'h002a 	:	o_val <= 16'b0000000010000101;
            14'h002b 	:	o_val <= 16'b0000000010001000;
            14'h002c 	:	o_val <= 16'b0000000010001011;
            14'h002d 	:	o_val <= 16'b0000000010001110;
            14'h002e 	:	o_val <= 16'b0000000010010010;
            14'h002f 	:	o_val <= 16'b0000000010010101;
            14'h0030 	:	o_val <= 16'b0000000010011000;
            14'h0031 	:	o_val <= 16'b0000000010011011;
            14'h0032 	:	o_val <= 16'b0000000010011110;
            14'h0033 	:	o_val <= 16'b0000000010100001;
            14'h0034 	:	o_val <= 16'b0000000010100100;
            14'h0035 	:	o_val <= 16'b0000000010101000;
            14'h0036 	:	o_val <= 16'b0000000010101011;
            14'h0037 	:	o_val <= 16'b0000000010101110;
            14'h0038 	:	o_val <= 16'b0000000010110001;
            14'h0039 	:	o_val <= 16'b0000000010110100;
            14'h003a 	:	o_val <= 16'b0000000010110111;
            14'h003b 	:	o_val <= 16'b0000000010111010;
            14'h003c 	:	o_val <= 16'b0000000010111110;
            14'h003d 	:	o_val <= 16'b0000000011000001;
            14'h003e 	:	o_val <= 16'b0000000011000100;
            14'h003f 	:	o_val <= 16'b0000000011000111;
            14'h0040 	:	o_val <= 16'b0000000011001010;
            14'h0041 	:	o_val <= 16'b0000000011001101;
            14'h0042 	:	o_val <= 16'b0000000011010000;
            14'h0043 	:	o_val <= 16'b0000000011010100;
            14'h0044 	:	o_val <= 16'b0000000011010111;
            14'h0045 	:	o_val <= 16'b0000000011011010;
            14'h0046 	:	o_val <= 16'b0000000011011101;
            14'h0047 	:	o_val <= 16'b0000000011100000;
            14'h0048 	:	o_val <= 16'b0000000011100011;
            14'h0049 	:	o_val <= 16'b0000000011100110;
            14'h004a 	:	o_val <= 16'b0000000011101010;
            14'h004b 	:	o_val <= 16'b0000000011101101;
            14'h004c 	:	o_val <= 16'b0000000011110000;
            14'h004d 	:	o_val <= 16'b0000000011110011;
            14'h004e 	:	o_val <= 16'b0000000011110110;
            14'h004f 	:	o_val <= 16'b0000000011111001;
            14'h0050 	:	o_val <= 16'b0000000011111100;
            14'h0051 	:	o_val <= 16'b0000000100000000;
            14'h0052 	:	o_val <= 16'b0000000100000011;
            14'h0053 	:	o_val <= 16'b0000000100000110;
            14'h0054 	:	o_val <= 16'b0000000100001001;
            14'h0055 	:	o_val <= 16'b0000000100001100;
            14'h0056 	:	o_val <= 16'b0000000100001111;
            14'h0057 	:	o_val <= 16'b0000000100010010;
            14'h0058 	:	o_val <= 16'b0000000100010110;
            14'h0059 	:	o_val <= 16'b0000000100011001;
            14'h005a 	:	o_val <= 16'b0000000100011100;
            14'h005b 	:	o_val <= 16'b0000000100011111;
            14'h005c 	:	o_val <= 16'b0000000100100010;
            14'h005d 	:	o_val <= 16'b0000000100100101;
            14'h005e 	:	o_val <= 16'b0000000100101000;
            14'h005f 	:	o_val <= 16'b0000000100101100;
            14'h0060 	:	o_val <= 16'b0000000100101111;
            14'h0061 	:	o_val <= 16'b0000000100110010;
            14'h0062 	:	o_val <= 16'b0000000100110101;
            14'h0063 	:	o_val <= 16'b0000000100111000;
            14'h0064 	:	o_val <= 16'b0000000100111011;
            14'h0065 	:	o_val <= 16'b0000000100111110;
            14'h0066 	:	o_val <= 16'b0000000101000010;
            14'h0067 	:	o_val <= 16'b0000000101000101;
            14'h0068 	:	o_val <= 16'b0000000101001000;
            14'h0069 	:	o_val <= 16'b0000000101001011;
            14'h006a 	:	o_val <= 16'b0000000101001110;
            14'h006b 	:	o_val <= 16'b0000000101010001;
            14'h006c 	:	o_val <= 16'b0000000101010100;
            14'h006d 	:	o_val <= 16'b0000000101010111;
            14'h006e 	:	o_val <= 16'b0000000101011011;
            14'h006f 	:	o_val <= 16'b0000000101011110;
            14'h0070 	:	o_val <= 16'b0000000101100001;
            14'h0071 	:	o_val <= 16'b0000000101100100;
            14'h0072 	:	o_val <= 16'b0000000101100111;
            14'h0073 	:	o_val <= 16'b0000000101101010;
            14'h0074 	:	o_val <= 16'b0000000101101101;
            14'h0075 	:	o_val <= 16'b0000000101110001;
            14'h0076 	:	o_val <= 16'b0000000101110100;
            14'h0077 	:	o_val <= 16'b0000000101110111;
            14'h0078 	:	o_val <= 16'b0000000101111010;
            14'h0079 	:	o_val <= 16'b0000000101111101;
            14'h007a 	:	o_val <= 16'b0000000110000000;
            14'h007b 	:	o_val <= 16'b0000000110000011;
            14'h007c 	:	o_val <= 16'b0000000110000111;
            14'h007d 	:	o_val <= 16'b0000000110001010;
            14'h007e 	:	o_val <= 16'b0000000110001101;
            14'h007f 	:	o_val <= 16'b0000000110010000;
            14'h0080 	:	o_val <= 16'b0000000110010011;
            14'h0081 	:	o_val <= 16'b0000000110010110;
            14'h0082 	:	o_val <= 16'b0000000110011001;
            14'h0083 	:	o_val <= 16'b0000000110011101;
            14'h0084 	:	o_val <= 16'b0000000110100000;
            14'h0085 	:	o_val <= 16'b0000000110100011;
            14'h0086 	:	o_val <= 16'b0000000110100110;
            14'h0087 	:	o_val <= 16'b0000000110101001;
            14'h0088 	:	o_val <= 16'b0000000110101100;
            14'h0089 	:	o_val <= 16'b0000000110101111;
            14'h008a 	:	o_val <= 16'b0000000110110011;
            14'h008b 	:	o_val <= 16'b0000000110110110;
            14'h008c 	:	o_val <= 16'b0000000110111001;
            14'h008d 	:	o_val <= 16'b0000000110111100;
            14'h008e 	:	o_val <= 16'b0000000110111111;
            14'h008f 	:	o_val <= 16'b0000000111000010;
            14'h0090 	:	o_val <= 16'b0000000111000101;
            14'h0091 	:	o_val <= 16'b0000000111001001;
            14'h0092 	:	o_val <= 16'b0000000111001100;
            14'h0093 	:	o_val <= 16'b0000000111001111;
            14'h0094 	:	o_val <= 16'b0000000111010010;
            14'h0095 	:	o_val <= 16'b0000000111010101;
            14'h0096 	:	o_val <= 16'b0000000111011000;
            14'h0097 	:	o_val <= 16'b0000000111011011;
            14'h0098 	:	o_val <= 16'b0000000111011111;
            14'h0099 	:	o_val <= 16'b0000000111100010;
            14'h009a 	:	o_val <= 16'b0000000111100101;
            14'h009b 	:	o_val <= 16'b0000000111101000;
            14'h009c 	:	o_val <= 16'b0000000111101011;
            14'h009d 	:	o_val <= 16'b0000000111101110;
            14'h009e 	:	o_val <= 16'b0000000111110001;
            14'h009f 	:	o_val <= 16'b0000000111110101;
            14'h00a0 	:	o_val <= 16'b0000000111111000;
            14'h00a1 	:	o_val <= 16'b0000000111111011;
            14'h00a2 	:	o_val <= 16'b0000000111111110;
            14'h00a3 	:	o_val <= 16'b0000001000000001;
            14'h00a4 	:	o_val <= 16'b0000001000000100;
            14'h00a5 	:	o_val <= 16'b0000001000000111;
            14'h00a6 	:	o_val <= 16'b0000001000001011;
            14'h00a7 	:	o_val <= 16'b0000001000001110;
            14'h00a8 	:	o_val <= 16'b0000001000010001;
            14'h00a9 	:	o_val <= 16'b0000001000010100;
            14'h00aa 	:	o_val <= 16'b0000001000010111;
            14'h00ab 	:	o_val <= 16'b0000001000011010;
            14'h00ac 	:	o_val <= 16'b0000001000011101;
            14'h00ad 	:	o_val <= 16'b0000001000100001;
            14'h00ae 	:	o_val <= 16'b0000001000100100;
            14'h00af 	:	o_val <= 16'b0000001000100111;
            14'h00b0 	:	o_val <= 16'b0000001000101010;
            14'h00b1 	:	o_val <= 16'b0000001000101101;
            14'h00b2 	:	o_val <= 16'b0000001000110000;
            14'h00b3 	:	o_val <= 16'b0000001000110011;
            14'h00b4 	:	o_val <= 16'b0000001000110111;
            14'h00b5 	:	o_val <= 16'b0000001000111010;
            14'h00b6 	:	o_val <= 16'b0000001000111101;
            14'h00b7 	:	o_val <= 16'b0000001001000000;
            14'h00b8 	:	o_val <= 16'b0000001001000011;
            14'h00b9 	:	o_val <= 16'b0000001001000110;
            14'h00ba 	:	o_val <= 16'b0000001001001001;
            14'h00bb 	:	o_val <= 16'b0000001001001101;
            14'h00bc 	:	o_val <= 16'b0000001001010000;
            14'h00bd 	:	o_val <= 16'b0000001001010011;
            14'h00be 	:	o_val <= 16'b0000001001010110;
            14'h00bf 	:	o_val <= 16'b0000001001011001;
            14'h00c0 	:	o_val <= 16'b0000001001011100;
            14'h00c1 	:	o_val <= 16'b0000001001011111;
            14'h00c2 	:	o_val <= 16'b0000001001100011;
            14'h00c3 	:	o_val <= 16'b0000001001100110;
            14'h00c4 	:	o_val <= 16'b0000001001101001;
            14'h00c5 	:	o_val <= 16'b0000001001101100;
            14'h00c6 	:	o_val <= 16'b0000001001101111;
            14'h00c7 	:	o_val <= 16'b0000001001110010;
            14'h00c8 	:	o_val <= 16'b0000001001110101;
            14'h00c9 	:	o_val <= 16'b0000001001111000;
            14'h00ca 	:	o_val <= 16'b0000001001111100;
            14'h00cb 	:	o_val <= 16'b0000001001111111;
            14'h00cc 	:	o_val <= 16'b0000001010000010;
            14'h00cd 	:	o_val <= 16'b0000001010000101;
            14'h00ce 	:	o_val <= 16'b0000001010001000;
            14'h00cf 	:	o_val <= 16'b0000001010001011;
            14'h00d0 	:	o_val <= 16'b0000001010001110;
            14'h00d1 	:	o_val <= 16'b0000001010010010;
            14'h00d2 	:	o_val <= 16'b0000001010010101;
            14'h00d3 	:	o_val <= 16'b0000001010011000;
            14'h00d4 	:	o_val <= 16'b0000001010011011;
            14'h00d5 	:	o_val <= 16'b0000001010011110;
            14'h00d6 	:	o_val <= 16'b0000001010100001;
            14'h00d7 	:	o_val <= 16'b0000001010100100;
            14'h00d8 	:	o_val <= 16'b0000001010101000;
            14'h00d9 	:	o_val <= 16'b0000001010101011;
            14'h00da 	:	o_val <= 16'b0000001010101110;
            14'h00db 	:	o_val <= 16'b0000001010110001;
            14'h00dc 	:	o_val <= 16'b0000001010110100;
            14'h00dd 	:	o_val <= 16'b0000001010110111;
            14'h00de 	:	o_val <= 16'b0000001010111010;
            14'h00df 	:	o_val <= 16'b0000001010111110;
            14'h00e0 	:	o_val <= 16'b0000001011000001;
            14'h00e1 	:	o_val <= 16'b0000001011000100;
            14'h00e2 	:	o_val <= 16'b0000001011000111;
            14'h00e3 	:	o_val <= 16'b0000001011001010;
            14'h00e4 	:	o_val <= 16'b0000001011001101;
            14'h00e5 	:	o_val <= 16'b0000001011010000;
            14'h00e6 	:	o_val <= 16'b0000001011010100;
            14'h00e7 	:	o_val <= 16'b0000001011010111;
            14'h00e8 	:	o_val <= 16'b0000001011011010;
            14'h00e9 	:	o_val <= 16'b0000001011011101;
            14'h00ea 	:	o_val <= 16'b0000001011100000;
            14'h00eb 	:	o_val <= 16'b0000001011100011;
            14'h00ec 	:	o_val <= 16'b0000001011100110;
            14'h00ed 	:	o_val <= 16'b0000001011101010;
            14'h00ee 	:	o_val <= 16'b0000001011101101;
            14'h00ef 	:	o_val <= 16'b0000001011110000;
            14'h00f0 	:	o_val <= 16'b0000001011110011;
            14'h00f1 	:	o_val <= 16'b0000001011110110;
            14'h00f2 	:	o_val <= 16'b0000001011111001;
            14'h00f3 	:	o_val <= 16'b0000001011111100;
            14'h00f4 	:	o_val <= 16'b0000001100000000;
            14'h00f5 	:	o_val <= 16'b0000001100000011;
            14'h00f6 	:	o_val <= 16'b0000001100000110;
            14'h00f7 	:	o_val <= 16'b0000001100001001;
            14'h00f8 	:	o_val <= 16'b0000001100001100;
            14'h00f9 	:	o_val <= 16'b0000001100001111;
            14'h00fa 	:	o_val <= 16'b0000001100010010;
            14'h00fb 	:	o_val <= 16'b0000001100010110;
            14'h00fc 	:	o_val <= 16'b0000001100011001;
            14'h00fd 	:	o_val <= 16'b0000001100011100;
            14'h00fe 	:	o_val <= 16'b0000001100011111;
            14'h00ff 	:	o_val <= 16'b0000001100100010;
            14'h0100 	:	o_val <= 16'b0000001100100101;
            14'h0101 	:	o_val <= 16'b0000001100101000;
            14'h0102 	:	o_val <= 16'b0000001100101100;
            14'h0103 	:	o_val <= 16'b0000001100101111;
            14'h0104 	:	o_val <= 16'b0000001100110010;
            14'h0105 	:	o_val <= 16'b0000001100110101;
            14'h0106 	:	o_val <= 16'b0000001100111000;
            14'h0107 	:	o_val <= 16'b0000001100111011;
            14'h0108 	:	o_val <= 16'b0000001100111110;
            14'h0109 	:	o_val <= 16'b0000001101000010;
            14'h010a 	:	o_val <= 16'b0000001101000101;
            14'h010b 	:	o_val <= 16'b0000001101001000;
            14'h010c 	:	o_val <= 16'b0000001101001011;
            14'h010d 	:	o_val <= 16'b0000001101001110;
            14'h010e 	:	o_val <= 16'b0000001101010001;
            14'h010f 	:	o_val <= 16'b0000001101010100;
            14'h0110 	:	o_val <= 16'b0000001101010111;
            14'h0111 	:	o_val <= 16'b0000001101011011;
            14'h0112 	:	o_val <= 16'b0000001101011110;
            14'h0113 	:	o_val <= 16'b0000001101100001;
            14'h0114 	:	o_val <= 16'b0000001101100100;
            14'h0115 	:	o_val <= 16'b0000001101100111;
            14'h0116 	:	o_val <= 16'b0000001101101010;
            14'h0117 	:	o_val <= 16'b0000001101101101;
            14'h0118 	:	o_val <= 16'b0000001101110001;
            14'h0119 	:	o_val <= 16'b0000001101110100;
            14'h011a 	:	o_val <= 16'b0000001101110111;
            14'h011b 	:	o_val <= 16'b0000001101111010;
            14'h011c 	:	o_val <= 16'b0000001101111101;
            14'h011d 	:	o_val <= 16'b0000001110000000;
            14'h011e 	:	o_val <= 16'b0000001110000011;
            14'h011f 	:	o_val <= 16'b0000001110000111;
            14'h0120 	:	o_val <= 16'b0000001110001010;
            14'h0121 	:	o_val <= 16'b0000001110001101;
            14'h0122 	:	o_val <= 16'b0000001110010000;
            14'h0123 	:	o_val <= 16'b0000001110010011;
            14'h0124 	:	o_val <= 16'b0000001110010110;
            14'h0125 	:	o_val <= 16'b0000001110011001;
            14'h0126 	:	o_val <= 16'b0000001110011101;
            14'h0127 	:	o_val <= 16'b0000001110100000;
            14'h0128 	:	o_val <= 16'b0000001110100011;
            14'h0129 	:	o_val <= 16'b0000001110100110;
            14'h012a 	:	o_val <= 16'b0000001110101001;
            14'h012b 	:	o_val <= 16'b0000001110101100;
            14'h012c 	:	o_val <= 16'b0000001110101111;
            14'h012d 	:	o_val <= 16'b0000001110110011;
            14'h012e 	:	o_val <= 16'b0000001110110110;
            14'h012f 	:	o_val <= 16'b0000001110111001;
            14'h0130 	:	o_val <= 16'b0000001110111100;
            14'h0131 	:	o_val <= 16'b0000001110111111;
            14'h0132 	:	o_val <= 16'b0000001111000010;
            14'h0133 	:	o_val <= 16'b0000001111000101;
            14'h0134 	:	o_val <= 16'b0000001111001001;
            14'h0135 	:	o_val <= 16'b0000001111001100;
            14'h0136 	:	o_val <= 16'b0000001111001111;
            14'h0137 	:	o_val <= 16'b0000001111010010;
            14'h0138 	:	o_val <= 16'b0000001111010101;
            14'h0139 	:	o_val <= 16'b0000001111011000;
            14'h013a 	:	o_val <= 16'b0000001111011011;
            14'h013b 	:	o_val <= 16'b0000001111011111;
            14'h013c 	:	o_val <= 16'b0000001111100010;
            14'h013d 	:	o_val <= 16'b0000001111100101;
            14'h013e 	:	o_val <= 16'b0000001111101000;
            14'h013f 	:	o_val <= 16'b0000001111101011;
            14'h0140 	:	o_val <= 16'b0000001111101110;
            14'h0141 	:	o_val <= 16'b0000001111110001;
            14'h0142 	:	o_val <= 16'b0000001111110101;
            14'h0143 	:	o_val <= 16'b0000001111111000;
            14'h0144 	:	o_val <= 16'b0000001111111011;
            14'h0145 	:	o_val <= 16'b0000001111111110;
            14'h0146 	:	o_val <= 16'b0000010000000001;
            14'h0147 	:	o_val <= 16'b0000010000000100;
            14'h0148 	:	o_val <= 16'b0000010000000111;
            14'h0149 	:	o_val <= 16'b0000010000001010;
            14'h014a 	:	o_val <= 16'b0000010000001110;
            14'h014b 	:	o_val <= 16'b0000010000010001;
            14'h014c 	:	o_val <= 16'b0000010000010100;
            14'h014d 	:	o_val <= 16'b0000010000010111;
            14'h014e 	:	o_val <= 16'b0000010000011010;
            14'h014f 	:	o_val <= 16'b0000010000011101;
            14'h0150 	:	o_val <= 16'b0000010000100000;
            14'h0151 	:	o_val <= 16'b0000010000100100;
            14'h0152 	:	o_val <= 16'b0000010000100111;
            14'h0153 	:	o_val <= 16'b0000010000101010;
            14'h0154 	:	o_val <= 16'b0000010000101101;
            14'h0155 	:	o_val <= 16'b0000010000110000;
            14'h0156 	:	o_val <= 16'b0000010000110011;
            14'h0157 	:	o_val <= 16'b0000010000110110;
            14'h0158 	:	o_val <= 16'b0000010000111010;
            14'h0159 	:	o_val <= 16'b0000010000111101;
            14'h015a 	:	o_val <= 16'b0000010001000000;
            14'h015b 	:	o_val <= 16'b0000010001000011;
            14'h015c 	:	o_val <= 16'b0000010001000110;
            14'h015d 	:	o_val <= 16'b0000010001001001;
            14'h015e 	:	o_val <= 16'b0000010001001100;
            14'h015f 	:	o_val <= 16'b0000010001010000;
            14'h0160 	:	o_val <= 16'b0000010001010011;
            14'h0161 	:	o_val <= 16'b0000010001010110;
            14'h0162 	:	o_val <= 16'b0000010001011001;
            14'h0163 	:	o_val <= 16'b0000010001011100;
            14'h0164 	:	o_val <= 16'b0000010001011111;
            14'h0165 	:	o_val <= 16'b0000010001100010;
            14'h0166 	:	o_val <= 16'b0000010001100110;
            14'h0167 	:	o_val <= 16'b0000010001101001;
            14'h0168 	:	o_val <= 16'b0000010001101100;
            14'h0169 	:	o_val <= 16'b0000010001101111;
            14'h016a 	:	o_val <= 16'b0000010001110010;
            14'h016b 	:	o_val <= 16'b0000010001110101;
            14'h016c 	:	o_val <= 16'b0000010001111000;
            14'h016d 	:	o_val <= 16'b0000010001111100;
            14'h016e 	:	o_val <= 16'b0000010001111111;
            14'h016f 	:	o_val <= 16'b0000010010000010;
            14'h0170 	:	o_val <= 16'b0000010010000101;
            14'h0171 	:	o_val <= 16'b0000010010001000;
            14'h0172 	:	o_val <= 16'b0000010010001011;
            14'h0173 	:	o_val <= 16'b0000010010001110;
            14'h0174 	:	o_val <= 16'b0000010010010001;
            14'h0175 	:	o_val <= 16'b0000010010010101;
            14'h0176 	:	o_val <= 16'b0000010010011000;
            14'h0177 	:	o_val <= 16'b0000010010011011;
            14'h0178 	:	o_val <= 16'b0000010010011110;
            14'h0179 	:	o_val <= 16'b0000010010100001;
            14'h017a 	:	o_val <= 16'b0000010010100100;
            14'h017b 	:	o_val <= 16'b0000010010100111;
            14'h017c 	:	o_val <= 16'b0000010010101011;
            14'h017d 	:	o_val <= 16'b0000010010101110;
            14'h017e 	:	o_val <= 16'b0000010010110001;
            14'h017f 	:	o_val <= 16'b0000010010110100;
            14'h0180 	:	o_val <= 16'b0000010010110111;
            14'h0181 	:	o_val <= 16'b0000010010111010;
            14'h0182 	:	o_val <= 16'b0000010010111101;
            14'h0183 	:	o_val <= 16'b0000010011000001;
            14'h0184 	:	o_val <= 16'b0000010011000100;
            14'h0185 	:	o_val <= 16'b0000010011000111;
            14'h0186 	:	o_val <= 16'b0000010011001010;
            14'h0187 	:	o_val <= 16'b0000010011001101;
            14'h0188 	:	o_val <= 16'b0000010011010000;
            14'h0189 	:	o_val <= 16'b0000010011010011;
            14'h018a 	:	o_val <= 16'b0000010011010111;
            14'h018b 	:	o_val <= 16'b0000010011011010;
            14'h018c 	:	o_val <= 16'b0000010011011101;
            14'h018d 	:	o_val <= 16'b0000010011100000;
            14'h018e 	:	o_val <= 16'b0000010011100011;
            14'h018f 	:	o_val <= 16'b0000010011100110;
            14'h0190 	:	o_val <= 16'b0000010011101001;
            14'h0191 	:	o_val <= 16'b0000010011101101;
            14'h0192 	:	o_val <= 16'b0000010011110000;
            14'h0193 	:	o_val <= 16'b0000010011110011;
            14'h0194 	:	o_val <= 16'b0000010011110110;
            14'h0195 	:	o_val <= 16'b0000010011111001;
            14'h0196 	:	o_val <= 16'b0000010011111100;
            14'h0197 	:	o_val <= 16'b0000010011111111;
            14'h0198 	:	o_val <= 16'b0000010100000011;
            14'h0199 	:	o_val <= 16'b0000010100000110;
            14'h019a 	:	o_val <= 16'b0000010100001001;
            14'h019b 	:	o_val <= 16'b0000010100001100;
            14'h019c 	:	o_val <= 16'b0000010100001111;
            14'h019d 	:	o_val <= 16'b0000010100010010;
            14'h019e 	:	o_val <= 16'b0000010100010101;
            14'h019f 	:	o_val <= 16'b0000010100011000;
            14'h01a0 	:	o_val <= 16'b0000010100011100;
            14'h01a1 	:	o_val <= 16'b0000010100011111;
            14'h01a2 	:	o_val <= 16'b0000010100100010;
            14'h01a3 	:	o_val <= 16'b0000010100100101;
            14'h01a4 	:	o_val <= 16'b0000010100101000;
            14'h01a5 	:	o_val <= 16'b0000010100101011;
            14'h01a6 	:	o_val <= 16'b0000010100101110;
            14'h01a7 	:	o_val <= 16'b0000010100110010;
            14'h01a8 	:	o_val <= 16'b0000010100110101;
            14'h01a9 	:	o_val <= 16'b0000010100111000;
            14'h01aa 	:	o_val <= 16'b0000010100111011;
            14'h01ab 	:	o_val <= 16'b0000010100111110;
            14'h01ac 	:	o_val <= 16'b0000010101000001;
            14'h01ad 	:	o_val <= 16'b0000010101000100;
            14'h01ae 	:	o_val <= 16'b0000010101001000;
            14'h01af 	:	o_val <= 16'b0000010101001011;
            14'h01b0 	:	o_val <= 16'b0000010101001110;
            14'h01b1 	:	o_val <= 16'b0000010101010001;
            14'h01b2 	:	o_val <= 16'b0000010101010100;
            14'h01b3 	:	o_val <= 16'b0000010101010111;
            14'h01b4 	:	o_val <= 16'b0000010101011010;
            14'h01b5 	:	o_val <= 16'b0000010101011110;
            14'h01b6 	:	o_val <= 16'b0000010101100001;
            14'h01b7 	:	o_val <= 16'b0000010101100100;
            14'h01b8 	:	o_val <= 16'b0000010101100111;
            14'h01b9 	:	o_val <= 16'b0000010101101010;
            14'h01ba 	:	o_val <= 16'b0000010101101101;
            14'h01bb 	:	o_val <= 16'b0000010101110000;
            14'h01bc 	:	o_val <= 16'b0000010101110100;
            14'h01bd 	:	o_val <= 16'b0000010101110111;
            14'h01be 	:	o_val <= 16'b0000010101111010;
            14'h01bf 	:	o_val <= 16'b0000010101111101;
            14'h01c0 	:	o_val <= 16'b0000010110000000;
            14'h01c1 	:	o_val <= 16'b0000010110000011;
            14'h01c2 	:	o_val <= 16'b0000010110000110;
            14'h01c3 	:	o_val <= 16'b0000010110001001;
            14'h01c4 	:	o_val <= 16'b0000010110001101;
            14'h01c5 	:	o_val <= 16'b0000010110010000;
            14'h01c6 	:	o_val <= 16'b0000010110010011;
            14'h01c7 	:	o_val <= 16'b0000010110010110;
            14'h01c8 	:	o_val <= 16'b0000010110011001;
            14'h01c9 	:	o_val <= 16'b0000010110011100;
            14'h01ca 	:	o_val <= 16'b0000010110011111;
            14'h01cb 	:	o_val <= 16'b0000010110100011;
            14'h01cc 	:	o_val <= 16'b0000010110100110;
            14'h01cd 	:	o_val <= 16'b0000010110101001;
            14'h01ce 	:	o_val <= 16'b0000010110101100;
            14'h01cf 	:	o_val <= 16'b0000010110101111;
            14'h01d0 	:	o_val <= 16'b0000010110110010;
            14'h01d1 	:	o_val <= 16'b0000010110110101;
            14'h01d2 	:	o_val <= 16'b0000010110111001;
            14'h01d3 	:	o_val <= 16'b0000010110111100;
            14'h01d4 	:	o_val <= 16'b0000010110111111;
            14'h01d5 	:	o_val <= 16'b0000010111000010;
            14'h01d6 	:	o_val <= 16'b0000010111000101;
            14'h01d7 	:	o_val <= 16'b0000010111001000;
            14'h01d8 	:	o_val <= 16'b0000010111001011;
            14'h01d9 	:	o_val <= 16'b0000010111001111;
            14'h01da 	:	o_val <= 16'b0000010111010010;
            14'h01db 	:	o_val <= 16'b0000010111010101;
            14'h01dc 	:	o_val <= 16'b0000010111011000;
            14'h01dd 	:	o_val <= 16'b0000010111011011;
            14'h01de 	:	o_val <= 16'b0000010111011110;
            14'h01df 	:	o_val <= 16'b0000010111100001;
            14'h01e0 	:	o_val <= 16'b0000010111100101;
            14'h01e1 	:	o_val <= 16'b0000010111101000;
            14'h01e2 	:	o_val <= 16'b0000010111101011;
            14'h01e3 	:	o_val <= 16'b0000010111101110;
            14'h01e4 	:	o_val <= 16'b0000010111110001;
            14'h01e5 	:	o_val <= 16'b0000010111110100;
            14'h01e6 	:	o_val <= 16'b0000010111110111;
            14'h01e7 	:	o_val <= 16'b0000010111111010;
            14'h01e8 	:	o_val <= 16'b0000010111111110;
            14'h01e9 	:	o_val <= 16'b0000011000000001;
            14'h01ea 	:	o_val <= 16'b0000011000000100;
            14'h01eb 	:	o_val <= 16'b0000011000000111;
            14'h01ec 	:	o_val <= 16'b0000011000001010;
            14'h01ed 	:	o_val <= 16'b0000011000001101;
            14'h01ee 	:	o_val <= 16'b0000011000010000;
            14'h01ef 	:	o_val <= 16'b0000011000010100;
            14'h01f0 	:	o_val <= 16'b0000011000010111;
            14'h01f1 	:	o_val <= 16'b0000011000011010;
            14'h01f2 	:	o_val <= 16'b0000011000011101;
            14'h01f3 	:	o_val <= 16'b0000011000100000;
            14'h01f4 	:	o_val <= 16'b0000011000100011;
            14'h01f5 	:	o_val <= 16'b0000011000100110;
            14'h01f6 	:	o_val <= 16'b0000011000101010;
            14'h01f7 	:	o_val <= 16'b0000011000101101;
            14'h01f8 	:	o_val <= 16'b0000011000110000;
            14'h01f9 	:	o_val <= 16'b0000011000110011;
            14'h01fa 	:	o_val <= 16'b0000011000110110;
            14'h01fb 	:	o_val <= 16'b0000011000111001;
            14'h01fc 	:	o_val <= 16'b0000011000111100;
            14'h01fd 	:	o_val <= 16'b0000011001000000;
            14'h01fe 	:	o_val <= 16'b0000011001000011;
            14'h01ff 	:	o_val <= 16'b0000011001000110;
            14'h0200 	:	o_val <= 16'b0000011001001001;
            14'h0201 	:	o_val <= 16'b0000011001001100;
            14'h0202 	:	o_val <= 16'b0000011001001111;
            14'h0203 	:	o_val <= 16'b0000011001010010;
            14'h0204 	:	o_val <= 16'b0000011001010101;
            14'h0205 	:	o_val <= 16'b0000011001011001;
            14'h0206 	:	o_val <= 16'b0000011001011100;
            14'h0207 	:	o_val <= 16'b0000011001011111;
            14'h0208 	:	o_val <= 16'b0000011001100010;
            14'h0209 	:	o_val <= 16'b0000011001100101;
            14'h020a 	:	o_val <= 16'b0000011001101000;
            14'h020b 	:	o_val <= 16'b0000011001101011;
            14'h020c 	:	o_val <= 16'b0000011001101111;
            14'h020d 	:	o_val <= 16'b0000011001110010;
            14'h020e 	:	o_val <= 16'b0000011001110101;
            14'h020f 	:	o_val <= 16'b0000011001111000;
            14'h0210 	:	o_val <= 16'b0000011001111011;
            14'h0211 	:	o_val <= 16'b0000011001111110;
            14'h0212 	:	o_val <= 16'b0000011010000001;
            14'h0213 	:	o_val <= 16'b0000011010000101;
            14'h0214 	:	o_val <= 16'b0000011010001000;
            14'h0215 	:	o_val <= 16'b0000011010001011;
            14'h0216 	:	o_val <= 16'b0000011010001110;
            14'h0217 	:	o_val <= 16'b0000011010010001;
            14'h0218 	:	o_val <= 16'b0000011010010100;
            14'h0219 	:	o_val <= 16'b0000011010010111;
            14'h021a 	:	o_val <= 16'b0000011010011010;
            14'h021b 	:	o_val <= 16'b0000011010011110;
            14'h021c 	:	o_val <= 16'b0000011010100001;
            14'h021d 	:	o_val <= 16'b0000011010100100;
            14'h021e 	:	o_val <= 16'b0000011010100111;
            14'h021f 	:	o_val <= 16'b0000011010101010;
            14'h0220 	:	o_val <= 16'b0000011010101101;
            14'h0221 	:	o_val <= 16'b0000011010110000;
            14'h0222 	:	o_val <= 16'b0000011010110100;
            14'h0223 	:	o_val <= 16'b0000011010110111;
            14'h0224 	:	o_val <= 16'b0000011010111010;
            14'h0225 	:	o_val <= 16'b0000011010111101;
            14'h0226 	:	o_val <= 16'b0000011011000000;
            14'h0227 	:	o_val <= 16'b0000011011000011;
            14'h0228 	:	o_val <= 16'b0000011011000110;
            14'h0229 	:	o_val <= 16'b0000011011001010;
            14'h022a 	:	o_val <= 16'b0000011011001101;
            14'h022b 	:	o_val <= 16'b0000011011010000;
            14'h022c 	:	o_val <= 16'b0000011011010011;
            14'h022d 	:	o_val <= 16'b0000011011010110;
            14'h022e 	:	o_val <= 16'b0000011011011001;
            14'h022f 	:	o_val <= 16'b0000011011011100;
            14'h0230 	:	o_val <= 16'b0000011011100000;
            14'h0231 	:	o_val <= 16'b0000011011100011;
            14'h0232 	:	o_val <= 16'b0000011011100110;
            14'h0233 	:	o_val <= 16'b0000011011101001;
            14'h0234 	:	o_val <= 16'b0000011011101100;
            14'h0235 	:	o_val <= 16'b0000011011101111;
            14'h0236 	:	o_val <= 16'b0000011011110010;
            14'h0237 	:	o_val <= 16'b0000011011110101;
            14'h0238 	:	o_val <= 16'b0000011011111001;
            14'h0239 	:	o_val <= 16'b0000011011111100;
            14'h023a 	:	o_val <= 16'b0000011011111111;
            14'h023b 	:	o_val <= 16'b0000011100000010;
            14'h023c 	:	o_val <= 16'b0000011100000101;
            14'h023d 	:	o_val <= 16'b0000011100001000;
            14'h023e 	:	o_val <= 16'b0000011100001011;
            14'h023f 	:	o_val <= 16'b0000011100001111;
            14'h0240 	:	o_val <= 16'b0000011100010010;
            14'h0241 	:	o_val <= 16'b0000011100010101;
            14'h0242 	:	o_val <= 16'b0000011100011000;
            14'h0243 	:	o_val <= 16'b0000011100011011;
            14'h0244 	:	o_val <= 16'b0000011100011110;
            14'h0245 	:	o_val <= 16'b0000011100100001;
            14'h0246 	:	o_val <= 16'b0000011100100101;
            14'h0247 	:	o_val <= 16'b0000011100101000;
            14'h0248 	:	o_val <= 16'b0000011100101011;
            14'h0249 	:	o_val <= 16'b0000011100101110;
            14'h024a 	:	o_val <= 16'b0000011100110001;
            14'h024b 	:	o_val <= 16'b0000011100110100;
            14'h024c 	:	o_val <= 16'b0000011100110111;
            14'h024d 	:	o_val <= 16'b0000011100111010;
            14'h024e 	:	o_val <= 16'b0000011100111110;
            14'h024f 	:	o_val <= 16'b0000011101000001;
            14'h0250 	:	o_val <= 16'b0000011101000100;
            14'h0251 	:	o_val <= 16'b0000011101000111;
            14'h0252 	:	o_val <= 16'b0000011101001010;
            14'h0253 	:	o_val <= 16'b0000011101001101;
            14'h0254 	:	o_val <= 16'b0000011101010000;
            14'h0255 	:	o_val <= 16'b0000011101010100;
            14'h0256 	:	o_val <= 16'b0000011101010111;
            14'h0257 	:	o_val <= 16'b0000011101011010;
            14'h0258 	:	o_val <= 16'b0000011101011101;
            14'h0259 	:	o_val <= 16'b0000011101100000;
            14'h025a 	:	o_val <= 16'b0000011101100011;
            14'h025b 	:	o_val <= 16'b0000011101100110;
            14'h025c 	:	o_val <= 16'b0000011101101010;
            14'h025d 	:	o_val <= 16'b0000011101101101;
            14'h025e 	:	o_val <= 16'b0000011101110000;
            14'h025f 	:	o_val <= 16'b0000011101110011;
            14'h0260 	:	o_val <= 16'b0000011101110110;
            14'h0261 	:	o_val <= 16'b0000011101111001;
            14'h0262 	:	o_val <= 16'b0000011101111100;
            14'h0263 	:	o_val <= 16'b0000011101111111;
            14'h0264 	:	o_val <= 16'b0000011110000011;
            14'h0265 	:	o_val <= 16'b0000011110000110;
            14'h0266 	:	o_val <= 16'b0000011110001001;
            14'h0267 	:	o_val <= 16'b0000011110001100;
            14'h0268 	:	o_val <= 16'b0000011110001111;
            14'h0269 	:	o_val <= 16'b0000011110010010;
            14'h026a 	:	o_val <= 16'b0000011110010101;
            14'h026b 	:	o_val <= 16'b0000011110011001;
            14'h026c 	:	o_val <= 16'b0000011110011100;
            14'h026d 	:	o_val <= 16'b0000011110011111;
            14'h026e 	:	o_val <= 16'b0000011110100010;
            14'h026f 	:	o_val <= 16'b0000011110100101;
            14'h0270 	:	o_val <= 16'b0000011110101000;
            14'h0271 	:	o_val <= 16'b0000011110101011;
            14'h0272 	:	o_val <= 16'b0000011110101111;
            14'h0273 	:	o_val <= 16'b0000011110110010;
            14'h0274 	:	o_val <= 16'b0000011110110101;
            14'h0275 	:	o_val <= 16'b0000011110111000;
            14'h0276 	:	o_val <= 16'b0000011110111011;
            14'h0277 	:	o_val <= 16'b0000011110111110;
            14'h0278 	:	o_val <= 16'b0000011111000001;
            14'h0279 	:	o_val <= 16'b0000011111000100;
            14'h027a 	:	o_val <= 16'b0000011111001000;
            14'h027b 	:	o_val <= 16'b0000011111001011;
            14'h027c 	:	o_val <= 16'b0000011111001110;
            14'h027d 	:	o_val <= 16'b0000011111010001;
            14'h027e 	:	o_val <= 16'b0000011111010100;
            14'h027f 	:	o_val <= 16'b0000011111010111;
            14'h0280 	:	o_val <= 16'b0000011111011010;
            14'h0281 	:	o_val <= 16'b0000011111011110;
            14'h0282 	:	o_val <= 16'b0000011111100001;
            14'h0283 	:	o_val <= 16'b0000011111100100;
            14'h0284 	:	o_val <= 16'b0000011111100111;
            14'h0285 	:	o_val <= 16'b0000011111101010;
            14'h0286 	:	o_val <= 16'b0000011111101101;
            14'h0287 	:	o_val <= 16'b0000011111110000;
            14'h0288 	:	o_val <= 16'b0000011111110100;
            14'h0289 	:	o_val <= 16'b0000011111110111;
            14'h028a 	:	o_val <= 16'b0000011111111010;
            14'h028b 	:	o_val <= 16'b0000011111111101;
            14'h028c 	:	o_val <= 16'b0000100000000000;
            14'h028d 	:	o_val <= 16'b0000100000000011;
            14'h028e 	:	o_val <= 16'b0000100000000110;
            14'h028f 	:	o_val <= 16'b0000100000001001;
            14'h0290 	:	o_val <= 16'b0000100000001101;
            14'h0291 	:	o_val <= 16'b0000100000010000;
            14'h0292 	:	o_val <= 16'b0000100000010011;
            14'h0293 	:	o_val <= 16'b0000100000010110;
            14'h0294 	:	o_val <= 16'b0000100000011001;
            14'h0295 	:	o_val <= 16'b0000100000011100;
            14'h0296 	:	o_val <= 16'b0000100000011111;
            14'h0297 	:	o_val <= 16'b0000100000100011;
            14'h0298 	:	o_val <= 16'b0000100000100110;
            14'h0299 	:	o_val <= 16'b0000100000101001;
            14'h029a 	:	o_val <= 16'b0000100000101100;
            14'h029b 	:	o_val <= 16'b0000100000101111;
            14'h029c 	:	o_val <= 16'b0000100000110010;
            14'h029d 	:	o_val <= 16'b0000100000110101;
            14'h029e 	:	o_val <= 16'b0000100000111000;
            14'h029f 	:	o_val <= 16'b0000100000111100;
            14'h02a0 	:	o_val <= 16'b0000100000111111;
            14'h02a1 	:	o_val <= 16'b0000100001000010;
            14'h02a2 	:	o_val <= 16'b0000100001000101;
            14'h02a3 	:	o_val <= 16'b0000100001001000;
            14'h02a4 	:	o_val <= 16'b0000100001001011;
            14'h02a5 	:	o_val <= 16'b0000100001001110;
            14'h02a6 	:	o_val <= 16'b0000100001010010;
            14'h02a7 	:	o_val <= 16'b0000100001010101;
            14'h02a8 	:	o_val <= 16'b0000100001011000;
            14'h02a9 	:	o_val <= 16'b0000100001011011;
            14'h02aa 	:	o_val <= 16'b0000100001011110;
            14'h02ab 	:	o_val <= 16'b0000100001100001;
            14'h02ac 	:	o_val <= 16'b0000100001100100;
            14'h02ad 	:	o_val <= 16'b0000100001101000;
            14'h02ae 	:	o_val <= 16'b0000100001101011;
            14'h02af 	:	o_val <= 16'b0000100001101110;
            14'h02b0 	:	o_val <= 16'b0000100001110001;
            14'h02b1 	:	o_val <= 16'b0000100001110100;
            14'h02b2 	:	o_val <= 16'b0000100001110111;
            14'h02b3 	:	o_val <= 16'b0000100001111010;
            14'h02b4 	:	o_val <= 16'b0000100001111101;
            14'h02b5 	:	o_val <= 16'b0000100010000001;
            14'h02b6 	:	o_val <= 16'b0000100010000100;
            14'h02b7 	:	o_val <= 16'b0000100010000111;
            14'h02b8 	:	o_val <= 16'b0000100010001010;
            14'h02b9 	:	o_val <= 16'b0000100010001101;
            14'h02ba 	:	o_val <= 16'b0000100010010000;
            14'h02bb 	:	o_val <= 16'b0000100010010011;
            14'h02bc 	:	o_val <= 16'b0000100010010111;
            14'h02bd 	:	o_val <= 16'b0000100010011010;
            14'h02be 	:	o_val <= 16'b0000100010011101;
            14'h02bf 	:	o_val <= 16'b0000100010100000;
            14'h02c0 	:	o_val <= 16'b0000100010100011;
            14'h02c1 	:	o_val <= 16'b0000100010100110;
            14'h02c2 	:	o_val <= 16'b0000100010101001;
            14'h02c3 	:	o_val <= 16'b0000100010101100;
            14'h02c4 	:	o_val <= 16'b0000100010110000;
            14'h02c5 	:	o_val <= 16'b0000100010110011;
            14'h02c6 	:	o_val <= 16'b0000100010110110;
            14'h02c7 	:	o_val <= 16'b0000100010111001;
            14'h02c8 	:	o_val <= 16'b0000100010111100;
            14'h02c9 	:	o_val <= 16'b0000100010111111;
            14'h02ca 	:	o_val <= 16'b0000100011000010;
            14'h02cb 	:	o_val <= 16'b0000100011000110;
            14'h02cc 	:	o_val <= 16'b0000100011001001;
            14'h02cd 	:	o_val <= 16'b0000100011001100;
            14'h02ce 	:	o_val <= 16'b0000100011001111;
            14'h02cf 	:	o_val <= 16'b0000100011010010;
            14'h02d0 	:	o_val <= 16'b0000100011010101;
            14'h02d1 	:	o_val <= 16'b0000100011011000;
            14'h02d2 	:	o_val <= 16'b0000100011011011;
            14'h02d3 	:	o_val <= 16'b0000100011011111;
            14'h02d4 	:	o_val <= 16'b0000100011100010;
            14'h02d5 	:	o_val <= 16'b0000100011100101;
            14'h02d6 	:	o_val <= 16'b0000100011101000;
            14'h02d7 	:	o_val <= 16'b0000100011101011;
            14'h02d8 	:	o_val <= 16'b0000100011101110;
            14'h02d9 	:	o_val <= 16'b0000100011110001;
            14'h02da 	:	o_val <= 16'b0000100011110101;
            14'h02db 	:	o_val <= 16'b0000100011111000;
            14'h02dc 	:	o_val <= 16'b0000100011111011;
            14'h02dd 	:	o_val <= 16'b0000100011111110;
            14'h02de 	:	o_val <= 16'b0000100100000001;
            14'h02df 	:	o_val <= 16'b0000100100000100;
            14'h02e0 	:	o_val <= 16'b0000100100000111;
            14'h02e1 	:	o_val <= 16'b0000100100001010;
            14'h02e2 	:	o_val <= 16'b0000100100001110;
            14'h02e3 	:	o_val <= 16'b0000100100010001;
            14'h02e4 	:	o_val <= 16'b0000100100010100;
            14'h02e5 	:	o_val <= 16'b0000100100010111;
            14'h02e6 	:	o_val <= 16'b0000100100011010;
            14'h02e7 	:	o_val <= 16'b0000100100011101;
            14'h02e8 	:	o_val <= 16'b0000100100100000;
            14'h02e9 	:	o_val <= 16'b0000100100100100;
            14'h02ea 	:	o_val <= 16'b0000100100100111;
            14'h02eb 	:	o_val <= 16'b0000100100101010;
            14'h02ec 	:	o_val <= 16'b0000100100101101;
            14'h02ed 	:	o_val <= 16'b0000100100110000;
            14'h02ee 	:	o_val <= 16'b0000100100110011;
            14'h02ef 	:	o_val <= 16'b0000100100110110;
            14'h02f0 	:	o_val <= 16'b0000100100111001;
            14'h02f1 	:	o_val <= 16'b0000100100111101;
            14'h02f2 	:	o_val <= 16'b0000100101000000;
            14'h02f3 	:	o_val <= 16'b0000100101000011;
            14'h02f4 	:	o_val <= 16'b0000100101000110;
            14'h02f5 	:	o_val <= 16'b0000100101001001;
            14'h02f6 	:	o_val <= 16'b0000100101001100;
            14'h02f7 	:	o_val <= 16'b0000100101001111;
            14'h02f8 	:	o_val <= 16'b0000100101010011;
            14'h02f9 	:	o_val <= 16'b0000100101010110;
            14'h02fa 	:	o_val <= 16'b0000100101011001;
            14'h02fb 	:	o_val <= 16'b0000100101011100;
            14'h02fc 	:	o_val <= 16'b0000100101011111;
            14'h02fd 	:	o_val <= 16'b0000100101100010;
            14'h02fe 	:	o_val <= 16'b0000100101100101;
            14'h02ff 	:	o_val <= 16'b0000100101101000;
            14'h0300 	:	o_val <= 16'b0000100101101100;
            14'h0301 	:	o_val <= 16'b0000100101101111;
            14'h0302 	:	o_val <= 16'b0000100101110010;
            14'h0303 	:	o_val <= 16'b0000100101110101;
            14'h0304 	:	o_val <= 16'b0000100101111000;
            14'h0305 	:	o_val <= 16'b0000100101111011;
            14'h0306 	:	o_val <= 16'b0000100101111110;
            14'h0307 	:	o_val <= 16'b0000100110000010;
            14'h0308 	:	o_val <= 16'b0000100110000101;
            14'h0309 	:	o_val <= 16'b0000100110001000;
            14'h030a 	:	o_val <= 16'b0000100110001011;
            14'h030b 	:	o_val <= 16'b0000100110001110;
            14'h030c 	:	o_val <= 16'b0000100110010001;
            14'h030d 	:	o_val <= 16'b0000100110010100;
            14'h030e 	:	o_val <= 16'b0000100110010111;
            14'h030f 	:	o_val <= 16'b0000100110011011;
            14'h0310 	:	o_val <= 16'b0000100110011110;
            14'h0311 	:	o_val <= 16'b0000100110100001;
            14'h0312 	:	o_val <= 16'b0000100110100100;
            14'h0313 	:	o_val <= 16'b0000100110100111;
            14'h0314 	:	o_val <= 16'b0000100110101010;
            14'h0315 	:	o_val <= 16'b0000100110101101;
            14'h0316 	:	o_val <= 16'b0000100110110001;
            14'h0317 	:	o_val <= 16'b0000100110110100;
            14'h0318 	:	o_val <= 16'b0000100110110111;
            14'h0319 	:	o_val <= 16'b0000100110111010;
            14'h031a 	:	o_val <= 16'b0000100110111101;
            14'h031b 	:	o_val <= 16'b0000100111000000;
            14'h031c 	:	o_val <= 16'b0000100111000011;
            14'h031d 	:	o_val <= 16'b0000100111000110;
            14'h031e 	:	o_val <= 16'b0000100111001010;
            14'h031f 	:	o_val <= 16'b0000100111001101;
            14'h0320 	:	o_val <= 16'b0000100111010000;
            14'h0321 	:	o_val <= 16'b0000100111010011;
            14'h0322 	:	o_val <= 16'b0000100111010110;
            14'h0323 	:	o_val <= 16'b0000100111011001;
            14'h0324 	:	o_val <= 16'b0000100111011100;
            14'h0325 	:	o_val <= 16'b0000100111100000;
            14'h0326 	:	o_val <= 16'b0000100111100011;
            14'h0327 	:	o_val <= 16'b0000100111100110;
            14'h0328 	:	o_val <= 16'b0000100111101001;
            14'h0329 	:	o_val <= 16'b0000100111101100;
            14'h032a 	:	o_val <= 16'b0000100111101111;
            14'h032b 	:	o_val <= 16'b0000100111110010;
            14'h032c 	:	o_val <= 16'b0000100111110101;
            14'h032d 	:	o_val <= 16'b0000100111111001;
            14'h032e 	:	o_val <= 16'b0000100111111100;
            14'h032f 	:	o_val <= 16'b0000100111111111;
            14'h0330 	:	o_val <= 16'b0000101000000010;
            14'h0331 	:	o_val <= 16'b0000101000000101;
            14'h0332 	:	o_val <= 16'b0000101000001000;
            14'h0333 	:	o_val <= 16'b0000101000001011;
            14'h0334 	:	o_val <= 16'b0000101000001111;
            14'h0335 	:	o_val <= 16'b0000101000010010;
            14'h0336 	:	o_val <= 16'b0000101000010101;
            14'h0337 	:	o_val <= 16'b0000101000011000;
            14'h0338 	:	o_val <= 16'b0000101000011011;
            14'h0339 	:	o_val <= 16'b0000101000011110;
            14'h033a 	:	o_val <= 16'b0000101000100001;
            14'h033b 	:	o_val <= 16'b0000101000100100;
            14'h033c 	:	o_val <= 16'b0000101000101000;
            14'h033d 	:	o_val <= 16'b0000101000101011;
            14'h033e 	:	o_val <= 16'b0000101000101110;
            14'h033f 	:	o_val <= 16'b0000101000110001;
            14'h0340 	:	o_val <= 16'b0000101000110100;
            14'h0341 	:	o_val <= 16'b0000101000110111;
            14'h0342 	:	o_val <= 16'b0000101000111010;
            14'h0343 	:	o_val <= 16'b0000101000111101;
            14'h0344 	:	o_val <= 16'b0000101001000001;
            14'h0345 	:	o_val <= 16'b0000101001000100;
            14'h0346 	:	o_val <= 16'b0000101001000111;
            14'h0347 	:	o_val <= 16'b0000101001001010;
            14'h0348 	:	o_val <= 16'b0000101001001101;
            14'h0349 	:	o_val <= 16'b0000101001010000;
            14'h034a 	:	o_val <= 16'b0000101001010011;
            14'h034b 	:	o_val <= 16'b0000101001010111;
            14'h034c 	:	o_val <= 16'b0000101001011010;
            14'h034d 	:	o_val <= 16'b0000101001011101;
            14'h034e 	:	o_val <= 16'b0000101001100000;
            14'h034f 	:	o_val <= 16'b0000101001100011;
            14'h0350 	:	o_val <= 16'b0000101001100110;
            14'h0351 	:	o_val <= 16'b0000101001101001;
            14'h0352 	:	o_val <= 16'b0000101001101100;
            14'h0353 	:	o_val <= 16'b0000101001110000;
            14'h0354 	:	o_val <= 16'b0000101001110011;
            14'h0355 	:	o_val <= 16'b0000101001110110;
            14'h0356 	:	o_val <= 16'b0000101001111001;
            14'h0357 	:	o_val <= 16'b0000101001111100;
            14'h0358 	:	o_val <= 16'b0000101001111111;
            14'h0359 	:	o_val <= 16'b0000101010000010;
            14'h035a 	:	o_val <= 16'b0000101010000110;
            14'h035b 	:	o_val <= 16'b0000101010001001;
            14'h035c 	:	o_val <= 16'b0000101010001100;
            14'h035d 	:	o_val <= 16'b0000101010001111;
            14'h035e 	:	o_val <= 16'b0000101010010010;
            14'h035f 	:	o_val <= 16'b0000101010010101;
            14'h0360 	:	o_val <= 16'b0000101010011000;
            14'h0361 	:	o_val <= 16'b0000101010011011;
            14'h0362 	:	o_val <= 16'b0000101010011111;
            14'h0363 	:	o_val <= 16'b0000101010100010;
            14'h0364 	:	o_val <= 16'b0000101010100101;
            14'h0365 	:	o_val <= 16'b0000101010101000;
            14'h0366 	:	o_val <= 16'b0000101010101011;
            14'h0367 	:	o_val <= 16'b0000101010101110;
            14'h0368 	:	o_val <= 16'b0000101010110001;
            14'h0369 	:	o_val <= 16'b0000101010110100;
            14'h036a 	:	o_val <= 16'b0000101010111000;
            14'h036b 	:	o_val <= 16'b0000101010111011;
            14'h036c 	:	o_val <= 16'b0000101010111110;
            14'h036d 	:	o_val <= 16'b0000101011000001;
            14'h036e 	:	o_val <= 16'b0000101011000100;
            14'h036f 	:	o_val <= 16'b0000101011000111;
            14'h0370 	:	o_val <= 16'b0000101011001010;
            14'h0371 	:	o_val <= 16'b0000101011001110;
            14'h0372 	:	o_val <= 16'b0000101011010001;
            14'h0373 	:	o_val <= 16'b0000101011010100;
            14'h0374 	:	o_val <= 16'b0000101011010111;
            14'h0375 	:	o_val <= 16'b0000101011011010;
            14'h0376 	:	o_val <= 16'b0000101011011101;
            14'h0377 	:	o_val <= 16'b0000101011100000;
            14'h0378 	:	o_val <= 16'b0000101011100011;
            14'h0379 	:	o_val <= 16'b0000101011100111;
            14'h037a 	:	o_val <= 16'b0000101011101010;
            14'h037b 	:	o_val <= 16'b0000101011101101;
            14'h037c 	:	o_val <= 16'b0000101011110000;
            14'h037d 	:	o_val <= 16'b0000101011110011;
            14'h037e 	:	o_val <= 16'b0000101011110110;
            14'h037f 	:	o_val <= 16'b0000101011111001;
            14'h0380 	:	o_val <= 16'b0000101011111100;
            14'h0381 	:	o_val <= 16'b0000101100000000;
            14'h0382 	:	o_val <= 16'b0000101100000011;
            14'h0383 	:	o_val <= 16'b0000101100000110;
            14'h0384 	:	o_val <= 16'b0000101100001001;
            14'h0385 	:	o_val <= 16'b0000101100001100;
            14'h0386 	:	o_val <= 16'b0000101100001111;
            14'h0387 	:	o_val <= 16'b0000101100010010;
            14'h0388 	:	o_val <= 16'b0000101100010110;
            14'h0389 	:	o_val <= 16'b0000101100011001;
            14'h038a 	:	o_val <= 16'b0000101100011100;
            14'h038b 	:	o_val <= 16'b0000101100011111;
            14'h038c 	:	o_val <= 16'b0000101100100010;
            14'h038d 	:	o_val <= 16'b0000101100100101;
            14'h038e 	:	o_val <= 16'b0000101100101000;
            14'h038f 	:	o_val <= 16'b0000101100101011;
            14'h0390 	:	o_val <= 16'b0000101100101111;
            14'h0391 	:	o_val <= 16'b0000101100110010;
            14'h0392 	:	o_val <= 16'b0000101100110101;
            14'h0393 	:	o_val <= 16'b0000101100111000;
            14'h0394 	:	o_val <= 16'b0000101100111011;
            14'h0395 	:	o_val <= 16'b0000101100111110;
            14'h0396 	:	o_val <= 16'b0000101101000001;
            14'h0397 	:	o_val <= 16'b0000101101000100;
            14'h0398 	:	o_val <= 16'b0000101101001000;
            14'h0399 	:	o_val <= 16'b0000101101001011;
            14'h039a 	:	o_val <= 16'b0000101101001110;
            14'h039b 	:	o_val <= 16'b0000101101010001;
            14'h039c 	:	o_val <= 16'b0000101101010100;
            14'h039d 	:	o_val <= 16'b0000101101010111;
            14'h039e 	:	o_val <= 16'b0000101101011010;
            14'h039f 	:	o_val <= 16'b0000101101011101;
            14'h03a0 	:	o_val <= 16'b0000101101100001;
            14'h03a1 	:	o_val <= 16'b0000101101100100;
            14'h03a2 	:	o_val <= 16'b0000101101100111;
            14'h03a3 	:	o_val <= 16'b0000101101101010;
            14'h03a4 	:	o_val <= 16'b0000101101101101;
            14'h03a5 	:	o_val <= 16'b0000101101110000;
            14'h03a6 	:	o_val <= 16'b0000101101110011;
            14'h03a7 	:	o_val <= 16'b0000101101110111;
            14'h03a8 	:	o_val <= 16'b0000101101111010;
            14'h03a9 	:	o_val <= 16'b0000101101111101;
            14'h03aa 	:	o_val <= 16'b0000101110000000;
            14'h03ab 	:	o_val <= 16'b0000101110000011;
            14'h03ac 	:	o_val <= 16'b0000101110000110;
            14'h03ad 	:	o_val <= 16'b0000101110001001;
            14'h03ae 	:	o_val <= 16'b0000101110001100;
            14'h03af 	:	o_val <= 16'b0000101110010000;
            14'h03b0 	:	o_val <= 16'b0000101110010011;
            14'h03b1 	:	o_val <= 16'b0000101110010110;
            14'h03b2 	:	o_val <= 16'b0000101110011001;
            14'h03b3 	:	o_val <= 16'b0000101110011100;
            14'h03b4 	:	o_val <= 16'b0000101110011111;
            14'h03b5 	:	o_val <= 16'b0000101110100010;
            14'h03b6 	:	o_val <= 16'b0000101110100101;
            14'h03b7 	:	o_val <= 16'b0000101110101001;
            14'h03b8 	:	o_val <= 16'b0000101110101100;
            14'h03b9 	:	o_val <= 16'b0000101110101111;
            14'h03ba 	:	o_val <= 16'b0000101110110010;
            14'h03bb 	:	o_val <= 16'b0000101110110101;
            14'h03bc 	:	o_val <= 16'b0000101110111000;
            14'h03bd 	:	o_val <= 16'b0000101110111011;
            14'h03be 	:	o_val <= 16'b0000101110111110;
            14'h03bf 	:	o_val <= 16'b0000101111000010;
            14'h03c0 	:	o_val <= 16'b0000101111000101;
            14'h03c1 	:	o_val <= 16'b0000101111001000;
            14'h03c2 	:	o_val <= 16'b0000101111001011;
            14'h03c3 	:	o_val <= 16'b0000101111001110;
            14'h03c4 	:	o_val <= 16'b0000101111010001;
            14'h03c5 	:	o_val <= 16'b0000101111010100;
            14'h03c6 	:	o_val <= 16'b0000101111011000;
            14'h03c7 	:	o_val <= 16'b0000101111011011;
            14'h03c8 	:	o_val <= 16'b0000101111011110;
            14'h03c9 	:	o_val <= 16'b0000101111100001;
            14'h03ca 	:	o_val <= 16'b0000101111100100;
            14'h03cb 	:	o_val <= 16'b0000101111100111;
            14'h03cc 	:	o_val <= 16'b0000101111101010;
            14'h03cd 	:	o_val <= 16'b0000101111101101;
            14'h03ce 	:	o_val <= 16'b0000101111110001;
            14'h03cf 	:	o_val <= 16'b0000101111110100;
            14'h03d0 	:	o_val <= 16'b0000101111110111;
            14'h03d1 	:	o_val <= 16'b0000101111111010;
            14'h03d2 	:	o_val <= 16'b0000101111111101;
            14'h03d3 	:	o_val <= 16'b0000110000000000;
            14'h03d4 	:	o_val <= 16'b0000110000000011;
            14'h03d5 	:	o_val <= 16'b0000110000000110;
            14'h03d6 	:	o_val <= 16'b0000110000001010;
            14'h03d7 	:	o_val <= 16'b0000110000001101;
            14'h03d8 	:	o_val <= 16'b0000110000010000;
            14'h03d9 	:	o_val <= 16'b0000110000010011;
            14'h03da 	:	o_val <= 16'b0000110000010110;
            14'h03db 	:	o_val <= 16'b0000110000011001;
            14'h03dc 	:	o_val <= 16'b0000110000011100;
            14'h03dd 	:	o_val <= 16'b0000110000011111;
            14'h03de 	:	o_val <= 16'b0000110000100011;
            14'h03df 	:	o_val <= 16'b0000110000100110;
            14'h03e0 	:	o_val <= 16'b0000110000101001;
            14'h03e1 	:	o_val <= 16'b0000110000101100;
            14'h03e2 	:	o_val <= 16'b0000110000101111;
            14'h03e3 	:	o_val <= 16'b0000110000110010;
            14'h03e4 	:	o_val <= 16'b0000110000110101;
            14'h03e5 	:	o_val <= 16'b0000110000111000;
            14'h03e6 	:	o_val <= 16'b0000110000111100;
            14'h03e7 	:	o_val <= 16'b0000110000111111;
            14'h03e8 	:	o_val <= 16'b0000110001000010;
            14'h03e9 	:	o_val <= 16'b0000110001000101;
            14'h03ea 	:	o_val <= 16'b0000110001001000;
            14'h03eb 	:	o_val <= 16'b0000110001001011;
            14'h03ec 	:	o_val <= 16'b0000110001001110;
            14'h03ed 	:	o_val <= 16'b0000110001010001;
            14'h03ee 	:	o_val <= 16'b0000110001010101;
            14'h03ef 	:	o_val <= 16'b0000110001011000;
            14'h03f0 	:	o_val <= 16'b0000110001011011;
            14'h03f1 	:	o_val <= 16'b0000110001011110;
            14'h03f2 	:	o_val <= 16'b0000110001100001;
            14'h03f3 	:	o_val <= 16'b0000110001100100;
            14'h03f4 	:	o_val <= 16'b0000110001100111;
            14'h03f5 	:	o_val <= 16'b0000110001101010;
            14'h03f6 	:	o_val <= 16'b0000110001101110;
            14'h03f7 	:	o_val <= 16'b0000110001110001;
            14'h03f8 	:	o_val <= 16'b0000110001110100;
            14'h03f9 	:	o_val <= 16'b0000110001110111;
            14'h03fa 	:	o_val <= 16'b0000110001111010;
            14'h03fb 	:	o_val <= 16'b0000110001111101;
            14'h03fc 	:	o_val <= 16'b0000110010000000;
            14'h03fd 	:	o_val <= 16'b0000110010000100;
            14'h03fe 	:	o_val <= 16'b0000110010000111;
            14'h03ff 	:	o_val <= 16'b0000110010001010;
            14'h0400 	:	o_val <= 16'b0000110010001101;
            14'h0401 	:	o_val <= 16'b0000110010010000;
            14'h0402 	:	o_val <= 16'b0000110010010011;
            14'h0403 	:	o_val <= 16'b0000110010010110;
            14'h0404 	:	o_val <= 16'b0000110010011001;
            14'h0405 	:	o_val <= 16'b0000110010011101;
            14'h0406 	:	o_val <= 16'b0000110010100000;
            14'h0407 	:	o_val <= 16'b0000110010100011;
            14'h0408 	:	o_val <= 16'b0000110010100110;
            14'h0409 	:	o_val <= 16'b0000110010101001;
            14'h040a 	:	o_val <= 16'b0000110010101100;
            14'h040b 	:	o_val <= 16'b0000110010101111;
            14'h040c 	:	o_val <= 16'b0000110010110010;
            14'h040d 	:	o_val <= 16'b0000110010110110;
            14'h040e 	:	o_val <= 16'b0000110010111001;
            14'h040f 	:	o_val <= 16'b0000110010111100;
            14'h0410 	:	o_val <= 16'b0000110010111111;
            14'h0411 	:	o_val <= 16'b0000110011000010;
            14'h0412 	:	o_val <= 16'b0000110011000101;
            14'h0413 	:	o_val <= 16'b0000110011001000;
            14'h0414 	:	o_val <= 16'b0000110011001011;
            14'h0415 	:	o_val <= 16'b0000110011001111;
            14'h0416 	:	o_val <= 16'b0000110011010010;
            14'h0417 	:	o_val <= 16'b0000110011010101;
            14'h0418 	:	o_val <= 16'b0000110011011000;
            14'h0419 	:	o_val <= 16'b0000110011011011;
            14'h041a 	:	o_val <= 16'b0000110011011110;
            14'h041b 	:	o_val <= 16'b0000110011100001;
            14'h041c 	:	o_val <= 16'b0000110011100100;
            14'h041d 	:	o_val <= 16'b0000110011101000;
            14'h041e 	:	o_val <= 16'b0000110011101011;
            14'h041f 	:	o_val <= 16'b0000110011101110;
            14'h0420 	:	o_val <= 16'b0000110011110001;
            14'h0421 	:	o_val <= 16'b0000110011110100;
            14'h0422 	:	o_val <= 16'b0000110011110111;
            14'h0423 	:	o_val <= 16'b0000110011111010;
            14'h0424 	:	o_val <= 16'b0000110011111101;
            14'h0425 	:	o_val <= 16'b0000110100000001;
            14'h0426 	:	o_val <= 16'b0000110100000100;
            14'h0427 	:	o_val <= 16'b0000110100000111;
            14'h0428 	:	o_val <= 16'b0000110100001010;
            14'h0429 	:	o_val <= 16'b0000110100001101;
            14'h042a 	:	o_val <= 16'b0000110100010000;
            14'h042b 	:	o_val <= 16'b0000110100010011;
            14'h042c 	:	o_val <= 16'b0000110100010110;
            14'h042d 	:	o_val <= 16'b0000110100011010;
            14'h042e 	:	o_val <= 16'b0000110100011101;
            14'h042f 	:	o_val <= 16'b0000110100100000;
            14'h0430 	:	o_val <= 16'b0000110100100011;
            14'h0431 	:	o_val <= 16'b0000110100100110;
            14'h0432 	:	o_val <= 16'b0000110100101001;
            14'h0433 	:	o_val <= 16'b0000110100101100;
            14'h0434 	:	o_val <= 16'b0000110100101111;
            14'h0435 	:	o_val <= 16'b0000110100110011;
            14'h0436 	:	o_val <= 16'b0000110100110110;
            14'h0437 	:	o_val <= 16'b0000110100111001;
            14'h0438 	:	o_val <= 16'b0000110100111100;
            14'h0439 	:	o_val <= 16'b0000110100111111;
            14'h043a 	:	o_val <= 16'b0000110101000010;
            14'h043b 	:	o_val <= 16'b0000110101000101;
            14'h043c 	:	o_val <= 16'b0000110101001000;
            14'h043d 	:	o_val <= 16'b0000110101001100;
            14'h043e 	:	o_val <= 16'b0000110101001111;
            14'h043f 	:	o_val <= 16'b0000110101010010;
            14'h0440 	:	o_val <= 16'b0000110101010101;
            14'h0441 	:	o_val <= 16'b0000110101011000;
            14'h0442 	:	o_val <= 16'b0000110101011011;
            14'h0443 	:	o_val <= 16'b0000110101011110;
            14'h0444 	:	o_val <= 16'b0000110101100001;
            14'h0445 	:	o_val <= 16'b0000110101100101;
            14'h0446 	:	o_val <= 16'b0000110101101000;
            14'h0447 	:	o_val <= 16'b0000110101101011;
            14'h0448 	:	o_val <= 16'b0000110101101110;
            14'h0449 	:	o_val <= 16'b0000110101110001;
            14'h044a 	:	o_val <= 16'b0000110101110100;
            14'h044b 	:	o_val <= 16'b0000110101110111;
            14'h044c 	:	o_val <= 16'b0000110101111010;
            14'h044d 	:	o_val <= 16'b0000110101111110;
            14'h044e 	:	o_val <= 16'b0000110110000001;
            14'h044f 	:	o_val <= 16'b0000110110000100;
            14'h0450 	:	o_val <= 16'b0000110110000111;
            14'h0451 	:	o_val <= 16'b0000110110001010;
            14'h0452 	:	o_val <= 16'b0000110110001101;
            14'h0453 	:	o_val <= 16'b0000110110010000;
            14'h0454 	:	o_val <= 16'b0000110110010011;
            14'h0455 	:	o_val <= 16'b0000110110010111;
            14'h0456 	:	o_val <= 16'b0000110110011010;
            14'h0457 	:	o_val <= 16'b0000110110011101;
            14'h0458 	:	o_val <= 16'b0000110110100000;
            14'h0459 	:	o_val <= 16'b0000110110100011;
            14'h045a 	:	o_val <= 16'b0000110110100110;
            14'h045b 	:	o_val <= 16'b0000110110101001;
            14'h045c 	:	o_val <= 16'b0000110110101100;
            14'h045d 	:	o_val <= 16'b0000110110110000;
            14'h045e 	:	o_val <= 16'b0000110110110011;
            14'h045f 	:	o_val <= 16'b0000110110110110;
            14'h0460 	:	o_val <= 16'b0000110110111001;
            14'h0461 	:	o_val <= 16'b0000110110111100;
            14'h0462 	:	o_val <= 16'b0000110110111111;
            14'h0463 	:	o_val <= 16'b0000110111000010;
            14'h0464 	:	o_val <= 16'b0000110111000101;
            14'h0465 	:	o_val <= 16'b0000110111001001;
            14'h0466 	:	o_val <= 16'b0000110111001100;
            14'h0467 	:	o_val <= 16'b0000110111001111;
            14'h0468 	:	o_val <= 16'b0000110111010010;
            14'h0469 	:	o_val <= 16'b0000110111010101;
            14'h046a 	:	o_val <= 16'b0000110111011000;
            14'h046b 	:	o_val <= 16'b0000110111011011;
            14'h046c 	:	o_val <= 16'b0000110111011110;
            14'h046d 	:	o_val <= 16'b0000110111100001;
            14'h046e 	:	o_val <= 16'b0000110111100101;
            14'h046f 	:	o_val <= 16'b0000110111101000;
            14'h0470 	:	o_val <= 16'b0000110111101011;
            14'h0471 	:	o_val <= 16'b0000110111101110;
            14'h0472 	:	o_val <= 16'b0000110111110001;
            14'h0473 	:	o_val <= 16'b0000110111110100;
            14'h0474 	:	o_val <= 16'b0000110111110111;
            14'h0475 	:	o_val <= 16'b0000110111111010;
            14'h0476 	:	o_val <= 16'b0000110111111110;
            14'h0477 	:	o_val <= 16'b0000111000000001;
            14'h0478 	:	o_val <= 16'b0000111000000100;
            14'h0479 	:	o_val <= 16'b0000111000000111;
            14'h047a 	:	o_val <= 16'b0000111000001010;
            14'h047b 	:	o_val <= 16'b0000111000001101;
            14'h047c 	:	o_val <= 16'b0000111000010000;
            14'h047d 	:	o_val <= 16'b0000111000010011;
            14'h047e 	:	o_val <= 16'b0000111000010111;
            14'h047f 	:	o_val <= 16'b0000111000011010;
            14'h0480 	:	o_val <= 16'b0000111000011101;
            14'h0481 	:	o_val <= 16'b0000111000100000;
            14'h0482 	:	o_val <= 16'b0000111000100011;
            14'h0483 	:	o_val <= 16'b0000111000100110;
            14'h0484 	:	o_val <= 16'b0000111000101001;
            14'h0485 	:	o_val <= 16'b0000111000101100;
            14'h0486 	:	o_val <= 16'b0000111000110000;
            14'h0487 	:	o_val <= 16'b0000111000110011;
            14'h0488 	:	o_val <= 16'b0000111000110110;
            14'h0489 	:	o_val <= 16'b0000111000111001;
            14'h048a 	:	o_val <= 16'b0000111000111100;
            14'h048b 	:	o_val <= 16'b0000111000111111;
            14'h048c 	:	o_val <= 16'b0000111001000010;
            14'h048d 	:	o_val <= 16'b0000111001000101;
            14'h048e 	:	o_val <= 16'b0000111001001001;
            14'h048f 	:	o_val <= 16'b0000111001001100;
            14'h0490 	:	o_val <= 16'b0000111001001111;
            14'h0491 	:	o_val <= 16'b0000111001010010;
            14'h0492 	:	o_val <= 16'b0000111001010101;
            14'h0493 	:	o_val <= 16'b0000111001011000;
            14'h0494 	:	o_val <= 16'b0000111001011011;
            14'h0495 	:	o_val <= 16'b0000111001011110;
            14'h0496 	:	o_val <= 16'b0000111001100010;
            14'h0497 	:	o_val <= 16'b0000111001100101;
            14'h0498 	:	o_val <= 16'b0000111001101000;
            14'h0499 	:	o_val <= 16'b0000111001101011;
            14'h049a 	:	o_val <= 16'b0000111001101110;
            14'h049b 	:	o_val <= 16'b0000111001110001;
            14'h049c 	:	o_val <= 16'b0000111001110100;
            14'h049d 	:	o_val <= 16'b0000111001110111;
            14'h049e 	:	o_val <= 16'b0000111001111010;
            14'h049f 	:	o_val <= 16'b0000111001111110;
            14'h04a0 	:	o_val <= 16'b0000111010000001;
            14'h04a1 	:	o_val <= 16'b0000111010000100;
            14'h04a2 	:	o_val <= 16'b0000111010000111;
            14'h04a3 	:	o_val <= 16'b0000111010001010;
            14'h04a4 	:	o_val <= 16'b0000111010001101;
            14'h04a5 	:	o_val <= 16'b0000111010010000;
            14'h04a6 	:	o_val <= 16'b0000111010010011;
            14'h04a7 	:	o_val <= 16'b0000111010010111;
            14'h04a8 	:	o_val <= 16'b0000111010011010;
            14'h04a9 	:	o_val <= 16'b0000111010011101;
            14'h04aa 	:	o_val <= 16'b0000111010100000;
            14'h04ab 	:	o_val <= 16'b0000111010100011;
            14'h04ac 	:	o_val <= 16'b0000111010100110;
            14'h04ad 	:	o_val <= 16'b0000111010101001;
            14'h04ae 	:	o_val <= 16'b0000111010101100;
            14'h04af 	:	o_val <= 16'b0000111010110000;
            14'h04b0 	:	o_val <= 16'b0000111010110011;
            14'h04b1 	:	o_val <= 16'b0000111010110110;
            14'h04b2 	:	o_val <= 16'b0000111010111001;
            14'h04b3 	:	o_val <= 16'b0000111010111100;
            14'h04b4 	:	o_val <= 16'b0000111010111111;
            14'h04b5 	:	o_val <= 16'b0000111011000010;
            14'h04b6 	:	o_val <= 16'b0000111011000101;
            14'h04b7 	:	o_val <= 16'b0000111011001001;
            14'h04b8 	:	o_val <= 16'b0000111011001100;
            14'h04b9 	:	o_val <= 16'b0000111011001111;
            14'h04ba 	:	o_val <= 16'b0000111011010010;
            14'h04bb 	:	o_val <= 16'b0000111011010101;
            14'h04bc 	:	o_val <= 16'b0000111011011000;
            14'h04bd 	:	o_val <= 16'b0000111011011011;
            14'h04be 	:	o_val <= 16'b0000111011011110;
            14'h04bf 	:	o_val <= 16'b0000111011100001;
            14'h04c0 	:	o_val <= 16'b0000111011100101;
            14'h04c1 	:	o_val <= 16'b0000111011101000;
            14'h04c2 	:	o_val <= 16'b0000111011101011;
            14'h04c3 	:	o_val <= 16'b0000111011101110;
            14'h04c4 	:	o_val <= 16'b0000111011110001;
            14'h04c5 	:	o_val <= 16'b0000111011110100;
            14'h04c6 	:	o_val <= 16'b0000111011110111;
            14'h04c7 	:	o_val <= 16'b0000111011111010;
            14'h04c8 	:	o_val <= 16'b0000111011111110;
            14'h04c9 	:	o_val <= 16'b0000111100000001;
            14'h04ca 	:	o_val <= 16'b0000111100000100;
            14'h04cb 	:	o_val <= 16'b0000111100000111;
            14'h04cc 	:	o_val <= 16'b0000111100001010;
            14'h04cd 	:	o_val <= 16'b0000111100001101;
            14'h04ce 	:	o_val <= 16'b0000111100010000;
            14'h04cf 	:	o_val <= 16'b0000111100010011;
            14'h04d0 	:	o_val <= 16'b0000111100010111;
            14'h04d1 	:	o_val <= 16'b0000111100011010;
            14'h04d2 	:	o_val <= 16'b0000111100011101;
            14'h04d3 	:	o_val <= 16'b0000111100100000;
            14'h04d4 	:	o_val <= 16'b0000111100100011;
            14'h04d5 	:	o_val <= 16'b0000111100100110;
            14'h04d6 	:	o_val <= 16'b0000111100101001;
            14'h04d7 	:	o_val <= 16'b0000111100101100;
            14'h04d8 	:	o_val <= 16'b0000111100101111;
            14'h04d9 	:	o_val <= 16'b0000111100110011;
            14'h04da 	:	o_val <= 16'b0000111100110110;
            14'h04db 	:	o_val <= 16'b0000111100111001;
            14'h04dc 	:	o_val <= 16'b0000111100111100;
            14'h04dd 	:	o_val <= 16'b0000111100111111;
            14'h04de 	:	o_val <= 16'b0000111101000010;
            14'h04df 	:	o_val <= 16'b0000111101000101;
            14'h04e0 	:	o_val <= 16'b0000111101001000;
            14'h04e1 	:	o_val <= 16'b0000111101001100;
            14'h04e2 	:	o_val <= 16'b0000111101001111;
            14'h04e3 	:	o_val <= 16'b0000111101010010;
            14'h04e4 	:	o_val <= 16'b0000111101010101;
            14'h04e5 	:	o_val <= 16'b0000111101011000;
            14'h04e6 	:	o_val <= 16'b0000111101011011;
            14'h04e7 	:	o_val <= 16'b0000111101011110;
            14'h04e8 	:	o_val <= 16'b0000111101100001;
            14'h04e9 	:	o_val <= 16'b0000111101100100;
            14'h04ea 	:	o_val <= 16'b0000111101101000;
            14'h04eb 	:	o_val <= 16'b0000111101101011;
            14'h04ec 	:	o_val <= 16'b0000111101101110;
            14'h04ed 	:	o_val <= 16'b0000111101110001;
            14'h04ee 	:	o_val <= 16'b0000111101110100;
            14'h04ef 	:	o_val <= 16'b0000111101110111;
            14'h04f0 	:	o_val <= 16'b0000111101111010;
            14'h04f1 	:	o_val <= 16'b0000111101111101;
            14'h04f2 	:	o_val <= 16'b0000111110000001;
            14'h04f3 	:	o_val <= 16'b0000111110000100;
            14'h04f4 	:	o_val <= 16'b0000111110000111;
            14'h04f5 	:	o_val <= 16'b0000111110001010;
            14'h04f6 	:	o_val <= 16'b0000111110001101;
            14'h04f7 	:	o_val <= 16'b0000111110010000;
            14'h04f8 	:	o_val <= 16'b0000111110010011;
            14'h04f9 	:	o_val <= 16'b0000111110010110;
            14'h04fa 	:	o_val <= 16'b0000111110011010;
            14'h04fb 	:	o_val <= 16'b0000111110011101;
            14'h04fc 	:	o_val <= 16'b0000111110100000;
            14'h04fd 	:	o_val <= 16'b0000111110100011;
            14'h04fe 	:	o_val <= 16'b0000111110100110;
            14'h04ff 	:	o_val <= 16'b0000111110101001;
            14'h0500 	:	o_val <= 16'b0000111110101100;
            14'h0501 	:	o_val <= 16'b0000111110101111;
            14'h0502 	:	o_val <= 16'b0000111110110010;
            14'h0503 	:	o_val <= 16'b0000111110110110;
            14'h0504 	:	o_val <= 16'b0000111110111001;
            14'h0505 	:	o_val <= 16'b0000111110111100;
            14'h0506 	:	o_val <= 16'b0000111110111111;
            14'h0507 	:	o_val <= 16'b0000111111000010;
            14'h0508 	:	o_val <= 16'b0000111111000101;
            14'h0509 	:	o_val <= 16'b0000111111001000;
            14'h050a 	:	o_val <= 16'b0000111111001011;
            14'h050b 	:	o_val <= 16'b0000111111001111;
            14'h050c 	:	o_val <= 16'b0000111111010010;
            14'h050d 	:	o_val <= 16'b0000111111010101;
            14'h050e 	:	o_val <= 16'b0000111111011000;
            14'h050f 	:	o_val <= 16'b0000111111011011;
            14'h0510 	:	o_val <= 16'b0000111111011110;
            14'h0511 	:	o_val <= 16'b0000111111100001;
            14'h0512 	:	o_val <= 16'b0000111111100100;
            14'h0513 	:	o_val <= 16'b0000111111100111;
            14'h0514 	:	o_val <= 16'b0000111111101011;
            14'h0515 	:	o_val <= 16'b0000111111101110;
            14'h0516 	:	o_val <= 16'b0000111111110001;
            14'h0517 	:	o_val <= 16'b0000111111110100;
            14'h0518 	:	o_val <= 16'b0000111111110111;
            14'h0519 	:	o_val <= 16'b0000111111111010;
            14'h051a 	:	o_val <= 16'b0000111111111101;
            14'h051b 	:	o_val <= 16'b0001000000000000;
            14'h051c 	:	o_val <= 16'b0001000000000011;
            14'h051d 	:	o_val <= 16'b0001000000000111;
            14'h051e 	:	o_val <= 16'b0001000000001010;
            14'h051f 	:	o_val <= 16'b0001000000001101;
            14'h0520 	:	o_val <= 16'b0001000000010000;
            14'h0521 	:	o_val <= 16'b0001000000010011;
            14'h0522 	:	o_val <= 16'b0001000000010110;
            14'h0523 	:	o_val <= 16'b0001000000011001;
            14'h0524 	:	o_val <= 16'b0001000000011100;
            14'h0525 	:	o_val <= 16'b0001000000100000;
            14'h0526 	:	o_val <= 16'b0001000000100011;
            14'h0527 	:	o_val <= 16'b0001000000100110;
            14'h0528 	:	o_val <= 16'b0001000000101001;
            14'h0529 	:	o_val <= 16'b0001000000101100;
            14'h052a 	:	o_val <= 16'b0001000000101111;
            14'h052b 	:	o_val <= 16'b0001000000110010;
            14'h052c 	:	o_val <= 16'b0001000000110101;
            14'h052d 	:	o_val <= 16'b0001000000111000;
            14'h052e 	:	o_val <= 16'b0001000000111100;
            14'h052f 	:	o_val <= 16'b0001000000111111;
            14'h0530 	:	o_val <= 16'b0001000001000010;
            14'h0531 	:	o_val <= 16'b0001000001000101;
            14'h0532 	:	o_val <= 16'b0001000001001000;
            14'h0533 	:	o_val <= 16'b0001000001001011;
            14'h0534 	:	o_val <= 16'b0001000001001110;
            14'h0535 	:	o_val <= 16'b0001000001010001;
            14'h0536 	:	o_val <= 16'b0001000001010101;
            14'h0537 	:	o_val <= 16'b0001000001011000;
            14'h0538 	:	o_val <= 16'b0001000001011011;
            14'h0539 	:	o_val <= 16'b0001000001011110;
            14'h053a 	:	o_val <= 16'b0001000001100001;
            14'h053b 	:	o_val <= 16'b0001000001100100;
            14'h053c 	:	o_val <= 16'b0001000001100111;
            14'h053d 	:	o_val <= 16'b0001000001101010;
            14'h053e 	:	o_val <= 16'b0001000001101101;
            14'h053f 	:	o_val <= 16'b0001000001110001;
            14'h0540 	:	o_val <= 16'b0001000001110100;
            14'h0541 	:	o_val <= 16'b0001000001110111;
            14'h0542 	:	o_val <= 16'b0001000001111010;
            14'h0543 	:	o_val <= 16'b0001000001111101;
            14'h0544 	:	o_val <= 16'b0001000010000000;
            14'h0545 	:	o_val <= 16'b0001000010000011;
            14'h0546 	:	o_val <= 16'b0001000010000110;
            14'h0547 	:	o_val <= 16'b0001000010001001;
            14'h0548 	:	o_val <= 16'b0001000010001101;
            14'h0549 	:	o_val <= 16'b0001000010010000;
            14'h054a 	:	o_val <= 16'b0001000010010011;
            14'h054b 	:	o_val <= 16'b0001000010010110;
            14'h054c 	:	o_val <= 16'b0001000010011001;
            14'h054d 	:	o_val <= 16'b0001000010011100;
            14'h054e 	:	o_val <= 16'b0001000010011111;
            14'h054f 	:	o_val <= 16'b0001000010100010;
            14'h0550 	:	o_val <= 16'b0001000010100110;
            14'h0551 	:	o_val <= 16'b0001000010101001;
            14'h0552 	:	o_val <= 16'b0001000010101100;
            14'h0553 	:	o_val <= 16'b0001000010101111;
            14'h0554 	:	o_val <= 16'b0001000010110010;
            14'h0555 	:	o_val <= 16'b0001000010110101;
            14'h0556 	:	o_val <= 16'b0001000010111000;
            14'h0557 	:	o_val <= 16'b0001000010111011;
            14'h0558 	:	o_val <= 16'b0001000010111110;
            14'h0559 	:	o_val <= 16'b0001000011000010;
            14'h055a 	:	o_val <= 16'b0001000011000101;
            14'h055b 	:	o_val <= 16'b0001000011001000;
            14'h055c 	:	o_val <= 16'b0001000011001011;
            14'h055d 	:	o_val <= 16'b0001000011001110;
            14'h055e 	:	o_val <= 16'b0001000011010001;
            14'h055f 	:	o_val <= 16'b0001000011010100;
            14'h0560 	:	o_val <= 16'b0001000011010111;
            14'h0561 	:	o_val <= 16'b0001000011011010;
            14'h0562 	:	o_val <= 16'b0001000011011110;
            14'h0563 	:	o_val <= 16'b0001000011100001;
            14'h0564 	:	o_val <= 16'b0001000011100100;
            14'h0565 	:	o_val <= 16'b0001000011100111;
            14'h0566 	:	o_val <= 16'b0001000011101010;
            14'h0567 	:	o_val <= 16'b0001000011101101;
            14'h0568 	:	o_val <= 16'b0001000011110000;
            14'h0569 	:	o_val <= 16'b0001000011110011;
            14'h056a 	:	o_val <= 16'b0001000011110111;
            14'h056b 	:	o_val <= 16'b0001000011111010;
            14'h056c 	:	o_val <= 16'b0001000011111101;
            14'h056d 	:	o_val <= 16'b0001000100000000;
            14'h056e 	:	o_val <= 16'b0001000100000011;
            14'h056f 	:	o_val <= 16'b0001000100000110;
            14'h0570 	:	o_val <= 16'b0001000100001001;
            14'h0571 	:	o_val <= 16'b0001000100001100;
            14'h0572 	:	o_val <= 16'b0001000100001111;
            14'h0573 	:	o_val <= 16'b0001000100010011;
            14'h0574 	:	o_val <= 16'b0001000100010110;
            14'h0575 	:	o_val <= 16'b0001000100011001;
            14'h0576 	:	o_val <= 16'b0001000100011100;
            14'h0577 	:	o_val <= 16'b0001000100011111;
            14'h0578 	:	o_val <= 16'b0001000100100010;
            14'h0579 	:	o_val <= 16'b0001000100100101;
            14'h057a 	:	o_val <= 16'b0001000100101000;
            14'h057b 	:	o_val <= 16'b0001000100101011;
            14'h057c 	:	o_val <= 16'b0001000100101111;
            14'h057d 	:	o_val <= 16'b0001000100110010;
            14'h057e 	:	o_val <= 16'b0001000100110101;
            14'h057f 	:	o_val <= 16'b0001000100111000;
            14'h0580 	:	o_val <= 16'b0001000100111011;
            14'h0581 	:	o_val <= 16'b0001000100111110;
            14'h0582 	:	o_val <= 16'b0001000101000001;
            14'h0583 	:	o_val <= 16'b0001000101000100;
            14'h0584 	:	o_val <= 16'b0001000101000111;
            14'h0585 	:	o_val <= 16'b0001000101001011;
            14'h0586 	:	o_val <= 16'b0001000101001110;
            14'h0587 	:	o_val <= 16'b0001000101010001;
            14'h0588 	:	o_val <= 16'b0001000101010100;
            14'h0589 	:	o_val <= 16'b0001000101010111;
            14'h058a 	:	o_val <= 16'b0001000101011010;
            14'h058b 	:	o_val <= 16'b0001000101011101;
            14'h058c 	:	o_val <= 16'b0001000101100000;
            14'h058d 	:	o_val <= 16'b0001000101100011;
            14'h058e 	:	o_val <= 16'b0001000101100111;
            14'h058f 	:	o_val <= 16'b0001000101101010;
            14'h0590 	:	o_val <= 16'b0001000101101101;
            14'h0591 	:	o_val <= 16'b0001000101110000;
            14'h0592 	:	o_val <= 16'b0001000101110011;
            14'h0593 	:	o_val <= 16'b0001000101110110;
            14'h0594 	:	o_val <= 16'b0001000101111001;
            14'h0595 	:	o_val <= 16'b0001000101111100;
            14'h0596 	:	o_val <= 16'b0001000101111111;
            14'h0597 	:	o_val <= 16'b0001000110000011;
            14'h0598 	:	o_val <= 16'b0001000110000110;
            14'h0599 	:	o_val <= 16'b0001000110001001;
            14'h059a 	:	o_val <= 16'b0001000110001100;
            14'h059b 	:	o_val <= 16'b0001000110001111;
            14'h059c 	:	o_val <= 16'b0001000110010010;
            14'h059d 	:	o_val <= 16'b0001000110010101;
            14'h059e 	:	o_val <= 16'b0001000110011000;
            14'h059f 	:	o_val <= 16'b0001000110011011;
            14'h05a0 	:	o_val <= 16'b0001000110011111;
            14'h05a1 	:	o_val <= 16'b0001000110100010;
            14'h05a2 	:	o_val <= 16'b0001000110100101;
            14'h05a3 	:	o_val <= 16'b0001000110101000;
            14'h05a4 	:	o_val <= 16'b0001000110101011;
            14'h05a5 	:	o_val <= 16'b0001000110101110;
            14'h05a6 	:	o_val <= 16'b0001000110110001;
            14'h05a7 	:	o_val <= 16'b0001000110110100;
            14'h05a8 	:	o_val <= 16'b0001000110110111;
            14'h05a9 	:	o_val <= 16'b0001000110111011;
            14'h05aa 	:	o_val <= 16'b0001000110111110;
            14'h05ab 	:	o_val <= 16'b0001000111000001;
            14'h05ac 	:	o_val <= 16'b0001000111000100;
            14'h05ad 	:	o_val <= 16'b0001000111000111;
            14'h05ae 	:	o_val <= 16'b0001000111001010;
            14'h05af 	:	o_val <= 16'b0001000111001101;
            14'h05b0 	:	o_val <= 16'b0001000111010000;
            14'h05b1 	:	o_val <= 16'b0001000111010011;
            14'h05b2 	:	o_val <= 16'b0001000111010111;
            14'h05b3 	:	o_val <= 16'b0001000111011010;
            14'h05b4 	:	o_val <= 16'b0001000111011101;
            14'h05b5 	:	o_val <= 16'b0001000111100000;
            14'h05b6 	:	o_val <= 16'b0001000111100011;
            14'h05b7 	:	o_val <= 16'b0001000111100110;
            14'h05b8 	:	o_val <= 16'b0001000111101001;
            14'h05b9 	:	o_val <= 16'b0001000111101100;
            14'h05ba 	:	o_val <= 16'b0001000111101111;
            14'h05bb 	:	o_val <= 16'b0001000111110011;
            14'h05bc 	:	o_val <= 16'b0001000111110110;
            14'h05bd 	:	o_val <= 16'b0001000111111001;
            14'h05be 	:	o_val <= 16'b0001000111111100;
            14'h05bf 	:	o_val <= 16'b0001000111111111;
            14'h05c0 	:	o_val <= 16'b0001001000000010;
            14'h05c1 	:	o_val <= 16'b0001001000000101;
            14'h05c2 	:	o_val <= 16'b0001001000001000;
            14'h05c3 	:	o_val <= 16'b0001001000001011;
            14'h05c4 	:	o_val <= 16'b0001001000001111;
            14'h05c5 	:	o_val <= 16'b0001001000010010;
            14'h05c6 	:	o_val <= 16'b0001001000010101;
            14'h05c7 	:	o_val <= 16'b0001001000011000;
            14'h05c8 	:	o_val <= 16'b0001001000011011;
            14'h05c9 	:	o_val <= 16'b0001001000011110;
            14'h05ca 	:	o_val <= 16'b0001001000100001;
            14'h05cb 	:	o_val <= 16'b0001001000100100;
            14'h05cc 	:	o_val <= 16'b0001001000100111;
            14'h05cd 	:	o_val <= 16'b0001001000101011;
            14'h05ce 	:	o_val <= 16'b0001001000101110;
            14'h05cf 	:	o_val <= 16'b0001001000110001;
            14'h05d0 	:	o_val <= 16'b0001001000110100;
            14'h05d1 	:	o_val <= 16'b0001001000110111;
            14'h05d2 	:	o_val <= 16'b0001001000111010;
            14'h05d3 	:	o_val <= 16'b0001001000111101;
            14'h05d4 	:	o_val <= 16'b0001001001000000;
            14'h05d5 	:	o_val <= 16'b0001001001000011;
            14'h05d6 	:	o_val <= 16'b0001001001000111;
            14'h05d7 	:	o_val <= 16'b0001001001001010;
            14'h05d8 	:	o_val <= 16'b0001001001001101;
            14'h05d9 	:	o_val <= 16'b0001001001010000;
            14'h05da 	:	o_val <= 16'b0001001001010011;
            14'h05db 	:	o_val <= 16'b0001001001010110;
            14'h05dc 	:	o_val <= 16'b0001001001011001;
            14'h05dd 	:	o_val <= 16'b0001001001011100;
            14'h05de 	:	o_val <= 16'b0001001001011111;
            14'h05df 	:	o_val <= 16'b0001001001100011;
            14'h05e0 	:	o_val <= 16'b0001001001100110;
            14'h05e1 	:	o_val <= 16'b0001001001101001;
            14'h05e2 	:	o_val <= 16'b0001001001101100;
            14'h05e3 	:	o_val <= 16'b0001001001101111;
            14'h05e4 	:	o_val <= 16'b0001001001110010;
            14'h05e5 	:	o_val <= 16'b0001001001110101;
            14'h05e6 	:	o_val <= 16'b0001001001111000;
            14'h05e7 	:	o_val <= 16'b0001001001111011;
            14'h05e8 	:	o_val <= 16'b0001001001111111;
            14'h05e9 	:	o_val <= 16'b0001001010000010;
            14'h05ea 	:	o_val <= 16'b0001001010000101;
            14'h05eb 	:	o_val <= 16'b0001001010001000;
            14'h05ec 	:	o_val <= 16'b0001001010001011;
            14'h05ed 	:	o_val <= 16'b0001001010001110;
            14'h05ee 	:	o_val <= 16'b0001001010010001;
            14'h05ef 	:	o_val <= 16'b0001001010010100;
            14'h05f0 	:	o_val <= 16'b0001001010010111;
            14'h05f1 	:	o_val <= 16'b0001001010011010;
            14'h05f2 	:	o_val <= 16'b0001001010011110;
            14'h05f3 	:	o_val <= 16'b0001001010100001;
            14'h05f4 	:	o_val <= 16'b0001001010100100;
            14'h05f5 	:	o_val <= 16'b0001001010100111;
            14'h05f6 	:	o_val <= 16'b0001001010101010;
            14'h05f7 	:	o_val <= 16'b0001001010101101;
            14'h05f8 	:	o_val <= 16'b0001001010110000;
            14'h05f9 	:	o_val <= 16'b0001001010110011;
            14'h05fa 	:	o_val <= 16'b0001001010110110;
            14'h05fb 	:	o_val <= 16'b0001001010111010;
            14'h05fc 	:	o_val <= 16'b0001001010111101;
            14'h05fd 	:	o_val <= 16'b0001001011000000;
            14'h05fe 	:	o_val <= 16'b0001001011000011;
            14'h05ff 	:	o_val <= 16'b0001001011000110;
            14'h0600 	:	o_val <= 16'b0001001011001001;
            14'h0601 	:	o_val <= 16'b0001001011001100;
            14'h0602 	:	o_val <= 16'b0001001011001111;
            14'h0603 	:	o_val <= 16'b0001001011010010;
            14'h0604 	:	o_val <= 16'b0001001011010110;
            14'h0605 	:	o_val <= 16'b0001001011011001;
            14'h0606 	:	o_val <= 16'b0001001011011100;
            14'h0607 	:	o_val <= 16'b0001001011011111;
            14'h0608 	:	o_val <= 16'b0001001011100010;
            14'h0609 	:	o_val <= 16'b0001001011100101;
            14'h060a 	:	o_val <= 16'b0001001011101000;
            14'h060b 	:	o_val <= 16'b0001001011101011;
            14'h060c 	:	o_val <= 16'b0001001011101110;
            14'h060d 	:	o_val <= 16'b0001001011110010;
            14'h060e 	:	o_val <= 16'b0001001011110101;
            14'h060f 	:	o_val <= 16'b0001001011111000;
            14'h0610 	:	o_val <= 16'b0001001011111011;
            14'h0611 	:	o_val <= 16'b0001001011111110;
            14'h0612 	:	o_val <= 16'b0001001100000001;
            14'h0613 	:	o_val <= 16'b0001001100000100;
            14'h0614 	:	o_val <= 16'b0001001100000111;
            14'h0615 	:	o_val <= 16'b0001001100001010;
            14'h0616 	:	o_val <= 16'b0001001100001101;
            14'h0617 	:	o_val <= 16'b0001001100010001;
            14'h0618 	:	o_val <= 16'b0001001100010100;
            14'h0619 	:	o_val <= 16'b0001001100010111;
            14'h061a 	:	o_val <= 16'b0001001100011010;
            14'h061b 	:	o_val <= 16'b0001001100011101;
            14'h061c 	:	o_val <= 16'b0001001100100000;
            14'h061d 	:	o_val <= 16'b0001001100100011;
            14'h061e 	:	o_val <= 16'b0001001100100110;
            14'h061f 	:	o_val <= 16'b0001001100101001;
            14'h0620 	:	o_val <= 16'b0001001100101101;
            14'h0621 	:	o_val <= 16'b0001001100110000;
            14'h0622 	:	o_val <= 16'b0001001100110011;
            14'h0623 	:	o_val <= 16'b0001001100110110;
            14'h0624 	:	o_val <= 16'b0001001100111001;
            14'h0625 	:	o_val <= 16'b0001001100111100;
            14'h0626 	:	o_val <= 16'b0001001100111111;
            14'h0627 	:	o_val <= 16'b0001001101000010;
            14'h0628 	:	o_val <= 16'b0001001101000101;
            14'h0629 	:	o_val <= 16'b0001001101001000;
            14'h062a 	:	o_val <= 16'b0001001101001100;
            14'h062b 	:	o_val <= 16'b0001001101001111;
            14'h062c 	:	o_val <= 16'b0001001101010010;
            14'h062d 	:	o_val <= 16'b0001001101010101;
            14'h062e 	:	o_val <= 16'b0001001101011000;
            14'h062f 	:	o_val <= 16'b0001001101011011;
            14'h0630 	:	o_val <= 16'b0001001101011110;
            14'h0631 	:	o_val <= 16'b0001001101100001;
            14'h0632 	:	o_val <= 16'b0001001101100100;
            14'h0633 	:	o_val <= 16'b0001001101101000;
            14'h0634 	:	o_val <= 16'b0001001101101011;
            14'h0635 	:	o_val <= 16'b0001001101101110;
            14'h0636 	:	o_val <= 16'b0001001101110001;
            14'h0637 	:	o_val <= 16'b0001001101110100;
            14'h0638 	:	o_val <= 16'b0001001101110111;
            14'h0639 	:	o_val <= 16'b0001001101111010;
            14'h063a 	:	o_val <= 16'b0001001101111101;
            14'h063b 	:	o_val <= 16'b0001001110000000;
            14'h063c 	:	o_val <= 16'b0001001110000011;
            14'h063d 	:	o_val <= 16'b0001001110000111;
            14'h063e 	:	o_val <= 16'b0001001110001010;
            14'h063f 	:	o_val <= 16'b0001001110001101;
            14'h0640 	:	o_val <= 16'b0001001110010000;
            14'h0641 	:	o_val <= 16'b0001001110010011;
            14'h0642 	:	o_val <= 16'b0001001110010110;
            14'h0643 	:	o_val <= 16'b0001001110011001;
            14'h0644 	:	o_val <= 16'b0001001110011100;
            14'h0645 	:	o_val <= 16'b0001001110011111;
            14'h0646 	:	o_val <= 16'b0001001110100011;
            14'h0647 	:	o_val <= 16'b0001001110100110;
            14'h0648 	:	o_val <= 16'b0001001110101001;
            14'h0649 	:	o_val <= 16'b0001001110101100;
            14'h064a 	:	o_val <= 16'b0001001110101111;
            14'h064b 	:	o_val <= 16'b0001001110110010;
            14'h064c 	:	o_val <= 16'b0001001110110101;
            14'h064d 	:	o_val <= 16'b0001001110111000;
            14'h064e 	:	o_val <= 16'b0001001110111011;
            14'h064f 	:	o_val <= 16'b0001001110111110;
            14'h0650 	:	o_val <= 16'b0001001111000010;
            14'h0651 	:	o_val <= 16'b0001001111000101;
            14'h0652 	:	o_val <= 16'b0001001111001000;
            14'h0653 	:	o_val <= 16'b0001001111001011;
            14'h0654 	:	o_val <= 16'b0001001111001110;
            14'h0655 	:	o_val <= 16'b0001001111010001;
            14'h0656 	:	o_val <= 16'b0001001111010100;
            14'h0657 	:	o_val <= 16'b0001001111010111;
            14'h0658 	:	o_val <= 16'b0001001111011010;
            14'h0659 	:	o_val <= 16'b0001001111011110;
            14'h065a 	:	o_val <= 16'b0001001111100001;
            14'h065b 	:	o_val <= 16'b0001001111100100;
            14'h065c 	:	o_val <= 16'b0001001111100111;
            14'h065d 	:	o_val <= 16'b0001001111101010;
            14'h065e 	:	o_val <= 16'b0001001111101101;
            14'h065f 	:	o_val <= 16'b0001001111110000;
            14'h0660 	:	o_val <= 16'b0001001111110011;
            14'h0661 	:	o_val <= 16'b0001001111110110;
            14'h0662 	:	o_val <= 16'b0001001111111001;
            14'h0663 	:	o_val <= 16'b0001001111111101;
            14'h0664 	:	o_val <= 16'b0001010000000000;
            14'h0665 	:	o_val <= 16'b0001010000000011;
            14'h0666 	:	o_val <= 16'b0001010000000110;
            14'h0667 	:	o_val <= 16'b0001010000001001;
            14'h0668 	:	o_val <= 16'b0001010000001100;
            14'h0669 	:	o_val <= 16'b0001010000001111;
            14'h066a 	:	o_val <= 16'b0001010000010010;
            14'h066b 	:	o_val <= 16'b0001010000010101;
            14'h066c 	:	o_val <= 16'b0001010000011000;
            14'h066d 	:	o_val <= 16'b0001010000011100;
            14'h066e 	:	o_val <= 16'b0001010000011111;
            14'h066f 	:	o_val <= 16'b0001010000100010;
            14'h0670 	:	o_val <= 16'b0001010000100101;
            14'h0671 	:	o_val <= 16'b0001010000101000;
            14'h0672 	:	o_val <= 16'b0001010000101011;
            14'h0673 	:	o_val <= 16'b0001010000101110;
            14'h0674 	:	o_val <= 16'b0001010000110001;
            14'h0675 	:	o_val <= 16'b0001010000110100;
            14'h0676 	:	o_val <= 16'b0001010000110111;
            14'h0677 	:	o_val <= 16'b0001010000111011;
            14'h0678 	:	o_val <= 16'b0001010000111110;
            14'h0679 	:	o_val <= 16'b0001010001000001;
            14'h067a 	:	o_val <= 16'b0001010001000100;
            14'h067b 	:	o_val <= 16'b0001010001000111;
            14'h067c 	:	o_val <= 16'b0001010001001010;
            14'h067d 	:	o_val <= 16'b0001010001001101;
            14'h067e 	:	o_val <= 16'b0001010001010000;
            14'h067f 	:	o_val <= 16'b0001010001010011;
            14'h0680 	:	o_val <= 16'b0001010001010111;
            14'h0681 	:	o_val <= 16'b0001010001011010;
            14'h0682 	:	o_val <= 16'b0001010001011101;
            14'h0683 	:	o_val <= 16'b0001010001100000;
            14'h0684 	:	o_val <= 16'b0001010001100011;
            14'h0685 	:	o_val <= 16'b0001010001100110;
            14'h0686 	:	o_val <= 16'b0001010001101001;
            14'h0687 	:	o_val <= 16'b0001010001101100;
            14'h0688 	:	o_val <= 16'b0001010001101111;
            14'h0689 	:	o_val <= 16'b0001010001110010;
            14'h068a 	:	o_val <= 16'b0001010001110110;
            14'h068b 	:	o_val <= 16'b0001010001111001;
            14'h068c 	:	o_val <= 16'b0001010001111100;
            14'h068d 	:	o_val <= 16'b0001010001111111;
            14'h068e 	:	o_val <= 16'b0001010010000010;
            14'h068f 	:	o_val <= 16'b0001010010000101;
            14'h0690 	:	o_val <= 16'b0001010010001000;
            14'h0691 	:	o_val <= 16'b0001010010001011;
            14'h0692 	:	o_val <= 16'b0001010010001110;
            14'h0693 	:	o_val <= 16'b0001010010010001;
            14'h0694 	:	o_val <= 16'b0001010010010101;
            14'h0695 	:	o_val <= 16'b0001010010011000;
            14'h0696 	:	o_val <= 16'b0001010010011011;
            14'h0697 	:	o_val <= 16'b0001010010011110;
            14'h0698 	:	o_val <= 16'b0001010010100001;
            14'h0699 	:	o_val <= 16'b0001010010100100;
            14'h069a 	:	o_val <= 16'b0001010010100111;
            14'h069b 	:	o_val <= 16'b0001010010101010;
            14'h069c 	:	o_val <= 16'b0001010010101101;
            14'h069d 	:	o_val <= 16'b0001010010110000;
            14'h069e 	:	o_val <= 16'b0001010010110100;
            14'h069f 	:	o_val <= 16'b0001010010110111;
            14'h06a0 	:	o_val <= 16'b0001010010111010;
            14'h06a1 	:	o_val <= 16'b0001010010111101;
            14'h06a2 	:	o_val <= 16'b0001010011000000;
            14'h06a3 	:	o_val <= 16'b0001010011000011;
            14'h06a4 	:	o_val <= 16'b0001010011000110;
            14'h06a5 	:	o_val <= 16'b0001010011001001;
            14'h06a6 	:	o_val <= 16'b0001010011001100;
            14'h06a7 	:	o_val <= 16'b0001010011001111;
            14'h06a8 	:	o_val <= 16'b0001010011010011;
            14'h06a9 	:	o_val <= 16'b0001010011010110;
            14'h06aa 	:	o_val <= 16'b0001010011011001;
            14'h06ab 	:	o_val <= 16'b0001010011011100;
            14'h06ac 	:	o_val <= 16'b0001010011011111;
            14'h06ad 	:	o_val <= 16'b0001010011100010;
            14'h06ae 	:	o_val <= 16'b0001010011100101;
            14'h06af 	:	o_val <= 16'b0001010011101000;
            14'h06b0 	:	o_val <= 16'b0001010011101011;
            14'h06b1 	:	o_val <= 16'b0001010011101110;
            14'h06b2 	:	o_val <= 16'b0001010011110010;
            14'h06b3 	:	o_val <= 16'b0001010011110101;
            14'h06b4 	:	o_val <= 16'b0001010011111000;
            14'h06b5 	:	o_val <= 16'b0001010011111011;
            14'h06b6 	:	o_val <= 16'b0001010011111110;
            14'h06b7 	:	o_val <= 16'b0001010100000001;
            14'h06b8 	:	o_val <= 16'b0001010100000100;
            14'h06b9 	:	o_val <= 16'b0001010100000111;
            14'h06ba 	:	o_val <= 16'b0001010100001010;
            14'h06bb 	:	o_val <= 16'b0001010100001101;
            14'h06bc 	:	o_val <= 16'b0001010100010001;
            14'h06bd 	:	o_val <= 16'b0001010100010100;
            14'h06be 	:	o_val <= 16'b0001010100010111;
            14'h06bf 	:	o_val <= 16'b0001010100011010;
            14'h06c0 	:	o_val <= 16'b0001010100011101;
            14'h06c1 	:	o_val <= 16'b0001010100100000;
            14'h06c2 	:	o_val <= 16'b0001010100100011;
            14'h06c3 	:	o_val <= 16'b0001010100100110;
            14'h06c4 	:	o_val <= 16'b0001010100101001;
            14'h06c5 	:	o_val <= 16'b0001010100101100;
            14'h06c6 	:	o_val <= 16'b0001010100110000;
            14'h06c7 	:	o_val <= 16'b0001010100110011;
            14'h06c8 	:	o_val <= 16'b0001010100110110;
            14'h06c9 	:	o_val <= 16'b0001010100111001;
            14'h06ca 	:	o_val <= 16'b0001010100111100;
            14'h06cb 	:	o_val <= 16'b0001010100111111;
            14'h06cc 	:	o_val <= 16'b0001010101000010;
            14'h06cd 	:	o_val <= 16'b0001010101000101;
            14'h06ce 	:	o_val <= 16'b0001010101001000;
            14'h06cf 	:	o_val <= 16'b0001010101001011;
            14'h06d0 	:	o_val <= 16'b0001010101001110;
            14'h06d1 	:	o_val <= 16'b0001010101010010;
            14'h06d2 	:	o_val <= 16'b0001010101010101;
            14'h06d3 	:	o_val <= 16'b0001010101011000;
            14'h06d4 	:	o_val <= 16'b0001010101011011;
            14'h06d5 	:	o_val <= 16'b0001010101011110;
            14'h06d6 	:	o_val <= 16'b0001010101100001;
            14'h06d7 	:	o_val <= 16'b0001010101100100;
            14'h06d8 	:	o_val <= 16'b0001010101100111;
            14'h06d9 	:	o_val <= 16'b0001010101101010;
            14'h06da 	:	o_val <= 16'b0001010101101101;
            14'h06db 	:	o_val <= 16'b0001010101110001;
            14'h06dc 	:	o_val <= 16'b0001010101110100;
            14'h06dd 	:	o_val <= 16'b0001010101110111;
            14'h06de 	:	o_val <= 16'b0001010101111010;
            14'h06df 	:	o_val <= 16'b0001010101111101;
            14'h06e0 	:	o_val <= 16'b0001010110000000;
            14'h06e1 	:	o_val <= 16'b0001010110000011;
            14'h06e2 	:	o_val <= 16'b0001010110000110;
            14'h06e3 	:	o_val <= 16'b0001010110001001;
            14'h06e4 	:	o_val <= 16'b0001010110001100;
            14'h06e5 	:	o_val <= 16'b0001010110010000;
            14'h06e6 	:	o_val <= 16'b0001010110010011;
            14'h06e7 	:	o_val <= 16'b0001010110010110;
            14'h06e8 	:	o_val <= 16'b0001010110011001;
            14'h06e9 	:	o_val <= 16'b0001010110011100;
            14'h06ea 	:	o_val <= 16'b0001010110011111;
            14'h06eb 	:	o_val <= 16'b0001010110100010;
            14'h06ec 	:	o_val <= 16'b0001010110100101;
            14'h06ed 	:	o_val <= 16'b0001010110101000;
            14'h06ee 	:	o_val <= 16'b0001010110101011;
            14'h06ef 	:	o_val <= 16'b0001010110101110;
            14'h06f0 	:	o_val <= 16'b0001010110110010;
            14'h06f1 	:	o_val <= 16'b0001010110110101;
            14'h06f2 	:	o_val <= 16'b0001010110111000;
            14'h06f3 	:	o_val <= 16'b0001010110111011;
            14'h06f4 	:	o_val <= 16'b0001010110111110;
            14'h06f5 	:	o_val <= 16'b0001010111000001;
            14'h06f6 	:	o_val <= 16'b0001010111000100;
            14'h06f7 	:	o_val <= 16'b0001010111000111;
            14'h06f8 	:	o_val <= 16'b0001010111001010;
            14'h06f9 	:	o_val <= 16'b0001010111001101;
            14'h06fa 	:	o_val <= 16'b0001010111010001;
            14'h06fb 	:	o_val <= 16'b0001010111010100;
            14'h06fc 	:	o_val <= 16'b0001010111010111;
            14'h06fd 	:	o_val <= 16'b0001010111011010;
            14'h06fe 	:	o_val <= 16'b0001010111011101;
            14'h06ff 	:	o_val <= 16'b0001010111100000;
            14'h0700 	:	o_val <= 16'b0001010111100011;
            14'h0701 	:	o_val <= 16'b0001010111100110;
            14'h0702 	:	o_val <= 16'b0001010111101001;
            14'h0703 	:	o_val <= 16'b0001010111101100;
            14'h0704 	:	o_val <= 16'b0001010111110000;
            14'h0705 	:	o_val <= 16'b0001010111110011;
            14'h0706 	:	o_val <= 16'b0001010111110110;
            14'h0707 	:	o_val <= 16'b0001010111111001;
            14'h0708 	:	o_val <= 16'b0001010111111100;
            14'h0709 	:	o_val <= 16'b0001010111111111;
            14'h070a 	:	o_val <= 16'b0001011000000010;
            14'h070b 	:	o_val <= 16'b0001011000000101;
            14'h070c 	:	o_val <= 16'b0001011000001000;
            14'h070d 	:	o_val <= 16'b0001011000001011;
            14'h070e 	:	o_val <= 16'b0001011000001110;
            14'h070f 	:	o_val <= 16'b0001011000010010;
            14'h0710 	:	o_val <= 16'b0001011000010101;
            14'h0711 	:	o_val <= 16'b0001011000011000;
            14'h0712 	:	o_val <= 16'b0001011000011011;
            14'h0713 	:	o_val <= 16'b0001011000011110;
            14'h0714 	:	o_val <= 16'b0001011000100001;
            14'h0715 	:	o_val <= 16'b0001011000100100;
            14'h0716 	:	o_val <= 16'b0001011000100111;
            14'h0717 	:	o_val <= 16'b0001011000101010;
            14'h0718 	:	o_val <= 16'b0001011000101101;
            14'h0719 	:	o_val <= 16'b0001011000110000;
            14'h071a 	:	o_val <= 16'b0001011000110100;
            14'h071b 	:	o_val <= 16'b0001011000110111;
            14'h071c 	:	o_val <= 16'b0001011000111010;
            14'h071d 	:	o_val <= 16'b0001011000111101;
            14'h071e 	:	o_val <= 16'b0001011001000000;
            14'h071f 	:	o_val <= 16'b0001011001000011;
            14'h0720 	:	o_val <= 16'b0001011001000110;
            14'h0721 	:	o_val <= 16'b0001011001001001;
            14'h0722 	:	o_val <= 16'b0001011001001100;
            14'h0723 	:	o_val <= 16'b0001011001001111;
            14'h0724 	:	o_val <= 16'b0001011001010011;
            14'h0725 	:	o_val <= 16'b0001011001010110;
            14'h0726 	:	o_val <= 16'b0001011001011001;
            14'h0727 	:	o_val <= 16'b0001011001011100;
            14'h0728 	:	o_val <= 16'b0001011001011111;
            14'h0729 	:	o_val <= 16'b0001011001100010;
            14'h072a 	:	o_val <= 16'b0001011001100101;
            14'h072b 	:	o_val <= 16'b0001011001101000;
            14'h072c 	:	o_val <= 16'b0001011001101011;
            14'h072d 	:	o_val <= 16'b0001011001101110;
            14'h072e 	:	o_val <= 16'b0001011001110001;
            14'h072f 	:	o_val <= 16'b0001011001110101;
            14'h0730 	:	o_val <= 16'b0001011001111000;
            14'h0731 	:	o_val <= 16'b0001011001111011;
            14'h0732 	:	o_val <= 16'b0001011001111110;
            14'h0733 	:	o_val <= 16'b0001011010000001;
            14'h0734 	:	o_val <= 16'b0001011010000100;
            14'h0735 	:	o_val <= 16'b0001011010000111;
            14'h0736 	:	o_val <= 16'b0001011010001010;
            14'h0737 	:	o_val <= 16'b0001011010001101;
            14'h0738 	:	o_val <= 16'b0001011010010000;
            14'h0739 	:	o_val <= 16'b0001011010010011;
            14'h073a 	:	o_val <= 16'b0001011010010111;
            14'h073b 	:	o_val <= 16'b0001011010011010;
            14'h073c 	:	o_val <= 16'b0001011010011101;
            14'h073d 	:	o_val <= 16'b0001011010100000;
            14'h073e 	:	o_val <= 16'b0001011010100011;
            14'h073f 	:	o_val <= 16'b0001011010100110;
            14'h0740 	:	o_val <= 16'b0001011010101001;
            14'h0741 	:	o_val <= 16'b0001011010101100;
            14'h0742 	:	o_val <= 16'b0001011010101111;
            14'h0743 	:	o_val <= 16'b0001011010110010;
            14'h0744 	:	o_val <= 16'b0001011010110101;
            14'h0745 	:	o_val <= 16'b0001011010111001;
            14'h0746 	:	o_val <= 16'b0001011010111100;
            14'h0747 	:	o_val <= 16'b0001011010111111;
            14'h0748 	:	o_val <= 16'b0001011011000010;
            14'h0749 	:	o_val <= 16'b0001011011000101;
            14'h074a 	:	o_val <= 16'b0001011011001000;
            14'h074b 	:	o_val <= 16'b0001011011001011;
            14'h074c 	:	o_val <= 16'b0001011011001110;
            14'h074d 	:	o_val <= 16'b0001011011010001;
            14'h074e 	:	o_val <= 16'b0001011011010100;
            14'h074f 	:	o_val <= 16'b0001011011010111;
            14'h0750 	:	o_val <= 16'b0001011011011011;
            14'h0751 	:	o_val <= 16'b0001011011011110;
            14'h0752 	:	o_val <= 16'b0001011011100001;
            14'h0753 	:	o_val <= 16'b0001011011100100;
            14'h0754 	:	o_val <= 16'b0001011011100111;
            14'h0755 	:	o_val <= 16'b0001011011101010;
            14'h0756 	:	o_val <= 16'b0001011011101101;
            14'h0757 	:	o_val <= 16'b0001011011110000;
            14'h0758 	:	o_val <= 16'b0001011011110011;
            14'h0759 	:	o_val <= 16'b0001011011110110;
            14'h075a 	:	o_val <= 16'b0001011011111001;
            14'h075b 	:	o_val <= 16'b0001011011111101;
            14'h075c 	:	o_val <= 16'b0001011100000000;
            14'h075d 	:	o_val <= 16'b0001011100000011;
            14'h075e 	:	o_val <= 16'b0001011100000110;
            14'h075f 	:	o_val <= 16'b0001011100001001;
            14'h0760 	:	o_val <= 16'b0001011100001100;
            14'h0761 	:	o_val <= 16'b0001011100001111;
            14'h0762 	:	o_val <= 16'b0001011100010010;
            14'h0763 	:	o_val <= 16'b0001011100010101;
            14'h0764 	:	o_val <= 16'b0001011100011000;
            14'h0765 	:	o_val <= 16'b0001011100011011;
            14'h0766 	:	o_val <= 16'b0001011100011111;
            14'h0767 	:	o_val <= 16'b0001011100100010;
            14'h0768 	:	o_val <= 16'b0001011100100101;
            14'h0769 	:	o_val <= 16'b0001011100101000;
            14'h076a 	:	o_val <= 16'b0001011100101011;
            14'h076b 	:	o_val <= 16'b0001011100101110;
            14'h076c 	:	o_val <= 16'b0001011100110001;
            14'h076d 	:	o_val <= 16'b0001011100110100;
            14'h076e 	:	o_val <= 16'b0001011100110111;
            14'h076f 	:	o_val <= 16'b0001011100111010;
            14'h0770 	:	o_val <= 16'b0001011100111101;
            14'h0771 	:	o_val <= 16'b0001011101000001;
            14'h0772 	:	o_val <= 16'b0001011101000100;
            14'h0773 	:	o_val <= 16'b0001011101000111;
            14'h0774 	:	o_val <= 16'b0001011101001010;
            14'h0775 	:	o_val <= 16'b0001011101001101;
            14'h0776 	:	o_val <= 16'b0001011101010000;
            14'h0777 	:	o_val <= 16'b0001011101010011;
            14'h0778 	:	o_val <= 16'b0001011101010110;
            14'h0779 	:	o_val <= 16'b0001011101011001;
            14'h077a 	:	o_val <= 16'b0001011101011100;
            14'h077b 	:	o_val <= 16'b0001011101011111;
            14'h077c 	:	o_val <= 16'b0001011101100011;
            14'h077d 	:	o_val <= 16'b0001011101100110;
            14'h077e 	:	o_val <= 16'b0001011101101001;
            14'h077f 	:	o_val <= 16'b0001011101101100;
            14'h0780 	:	o_val <= 16'b0001011101101111;
            14'h0781 	:	o_val <= 16'b0001011101110010;
            14'h0782 	:	o_val <= 16'b0001011101110101;
            14'h0783 	:	o_val <= 16'b0001011101111000;
            14'h0784 	:	o_val <= 16'b0001011101111011;
            14'h0785 	:	o_val <= 16'b0001011101111110;
            14'h0786 	:	o_val <= 16'b0001011110000001;
            14'h0787 	:	o_val <= 16'b0001011110000101;
            14'h0788 	:	o_val <= 16'b0001011110001000;
            14'h0789 	:	o_val <= 16'b0001011110001011;
            14'h078a 	:	o_val <= 16'b0001011110001110;
            14'h078b 	:	o_val <= 16'b0001011110010001;
            14'h078c 	:	o_val <= 16'b0001011110010100;
            14'h078d 	:	o_val <= 16'b0001011110010111;
            14'h078e 	:	o_val <= 16'b0001011110011010;
            14'h078f 	:	o_val <= 16'b0001011110011101;
            14'h0790 	:	o_val <= 16'b0001011110100000;
            14'h0791 	:	o_val <= 16'b0001011110100011;
            14'h0792 	:	o_val <= 16'b0001011110100110;
            14'h0793 	:	o_val <= 16'b0001011110101010;
            14'h0794 	:	o_val <= 16'b0001011110101101;
            14'h0795 	:	o_val <= 16'b0001011110110000;
            14'h0796 	:	o_val <= 16'b0001011110110011;
            14'h0797 	:	o_val <= 16'b0001011110110110;
            14'h0798 	:	o_val <= 16'b0001011110111001;
            14'h0799 	:	o_val <= 16'b0001011110111100;
            14'h079a 	:	o_val <= 16'b0001011110111111;
            14'h079b 	:	o_val <= 16'b0001011111000010;
            14'h079c 	:	o_val <= 16'b0001011111000101;
            14'h079d 	:	o_val <= 16'b0001011111001000;
            14'h079e 	:	o_val <= 16'b0001011111001100;
            14'h079f 	:	o_val <= 16'b0001011111001111;
            14'h07a0 	:	o_val <= 16'b0001011111010010;
            14'h07a1 	:	o_val <= 16'b0001011111010101;
            14'h07a2 	:	o_val <= 16'b0001011111011000;
            14'h07a3 	:	o_val <= 16'b0001011111011011;
            14'h07a4 	:	o_val <= 16'b0001011111011110;
            14'h07a5 	:	o_val <= 16'b0001011111100001;
            14'h07a6 	:	o_val <= 16'b0001011111100100;
            14'h07a7 	:	o_val <= 16'b0001011111100111;
            14'h07a8 	:	o_val <= 16'b0001011111101010;
            14'h07a9 	:	o_val <= 16'b0001011111101101;
            14'h07aa 	:	o_val <= 16'b0001011111110001;
            14'h07ab 	:	o_val <= 16'b0001011111110100;
            14'h07ac 	:	o_val <= 16'b0001011111110111;
            14'h07ad 	:	o_val <= 16'b0001011111111010;
            14'h07ae 	:	o_val <= 16'b0001011111111101;
            14'h07af 	:	o_val <= 16'b0001100000000000;
            14'h07b0 	:	o_val <= 16'b0001100000000011;
            14'h07b1 	:	o_val <= 16'b0001100000000110;
            14'h07b2 	:	o_val <= 16'b0001100000001001;
            14'h07b3 	:	o_val <= 16'b0001100000001100;
            14'h07b4 	:	o_val <= 16'b0001100000001111;
            14'h07b5 	:	o_val <= 16'b0001100000010011;
            14'h07b6 	:	o_val <= 16'b0001100000010110;
            14'h07b7 	:	o_val <= 16'b0001100000011001;
            14'h07b8 	:	o_val <= 16'b0001100000011100;
            14'h07b9 	:	o_val <= 16'b0001100000011111;
            14'h07ba 	:	o_val <= 16'b0001100000100010;
            14'h07bb 	:	o_val <= 16'b0001100000100101;
            14'h07bc 	:	o_val <= 16'b0001100000101000;
            14'h07bd 	:	o_val <= 16'b0001100000101011;
            14'h07be 	:	o_val <= 16'b0001100000101110;
            14'h07bf 	:	o_val <= 16'b0001100000110001;
            14'h07c0 	:	o_val <= 16'b0001100000110100;
            14'h07c1 	:	o_val <= 16'b0001100000111000;
            14'h07c2 	:	o_val <= 16'b0001100000111011;
            14'h07c3 	:	o_val <= 16'b0001100000111110;
            14'h07c4 	:	o_val <= 16'b0001100001000001;
            14'h07c5 	:	o_val <= 16'b0001100001000100;
            14'h07c6 	:	o_val <= 16'b0001100001000111;
            14'h07c7 	:	o_val <= 16'b0001100001001010;
            14'h07c8 	:	o_val <= 16'b0001100001001101;
            14'h07c9 	:	o_val <= 16'b0001100001010000;
            14'h07ca 	:	o_val <= 16'b0001100001010011;
            14'h07cb 	:	o_val <= 16'b0001100001010110;
            14'h07cc 	:	o_val <= 16'b0001100001011001;
            14'h07cd 	:	o_val <= 16'b0001100001011101;
            14'h07ce 	:	o_val <= 16'b0001100001100000;
            14'h07cf 	:	o_val <= 16'b0001100001100011;
            14'h07d0 	:	o_val <= 16'b0001100001100110;
            14'h07d1 	:	o_val <= 16'b0001100001101001;
            14'h07d2 	:	o_val <= 16'b0001100001101100;
            14'h07d3 	:	o_val <= 16'b0001100001101111;
            14'h07d4 	:	o_val <= 16'b0001100001110010;
            14'h07d5 	:	o_val <= 16'b0001100001110101;
            14'h07d6 	:	o_val <= 16'b0001100001111000;
            14'h07d7 	:	o_val <= 16'b0001100001111011;
            14'h07d8 	:	o_val <= 16'b0001100001111110;
            14'h07d9 	:	o_val <= 16'b0001100010000010;
            14'h07da 	:	o_val <= 16'b0001100010000101;
            14'h07db 	:	o_val <= 16'b0001100010001000;
            14'h07dc 	:	o_val <= 16'b0001100010001011;
            14'h07dd 	:	o_val <= 16'b0001100010001110;
            14'h07de 	:	o_val <= 16'b0001100010010001;
            14'h07df 	:	o_val <= 16'b0001100010010100;
            14'h07e0 	:	o_val <= 16'b0001100010010111;
            14'h07e1 	:	o_val <= 16'b0001100010011010;
            14'h07e2 	:	o_val <= 16'b0001100010011101;
            14'h07e3 	:	o_val <= 16'b0001100010100000;
            14'h07e4 	:	o_val <= 16'b0001100010100011;
            14'h07e5 	:	o_val <= 16'b0001100010100111;
            14'h07e6 	:	o_val <= 16'b0001100010101010;
            14'h07e7 	:	o_val <= 16'b0001100010101101;
            14'h07e8 	:	o_val <= 16'b0001100010110000;
            14'h07e9 	:	o_val <= 16'b0001100010110011;
            14'h07ea 	:	o_val <= 16'b0001100010110110;
            14'h07eb 	:	o_val <= 16'b0001100010111001;
            14'h07ec 	:	o_val <= 16'b0001100010111100;
            14'h07ed 	:	o_val <= 16'b0001100010111111;
            14'h07ee 	:	o_val <= 16'b0001100011000010;
            14'h07ef 	:	o_val <= 16'b0001100011000101;
            14'h07f0 	:	o_val <= 16'b0001100011001000;
            14'h07f1 	:	o_val <= 16'b0001100011001100;
            14'h07f2 	:	o_val <= 16'b0001100011001111;
            14'h07f3 	:	o_val <= 16'b0001100011010010;
            14'h07f4 	:	o_val <= 16'b0001100011010101;
            14'h07f5 	:	o_val <= 16'b0001100011011000;
            14'h07f6 	:	o_val <= 16'b0001100011011011;
            14'h07f7 	:	o_val <= 16'b0001100011011110;
            14'h07f8 	:	o_val <= 16'b0001100011100001;
            14'h07f9 	:	o_val <= 16'b0001100011100100;
            14'h07fa 	:	o_val <= 16'b0001100011100111;
            14'h07fb 	:	o_val <= 16'b0001100011101010;
            14'h07fc 	:	o_val <= 16'b0001100011101101;
            14'h07fd 	:	o_val <= 16'b0001100011110001;
            14'h07fe 	:	o_val <= 16'b0001100011110100;
            14'h07ff 	:	o_val <= 16'b0001100011110111;
            14'h0800 	:	o_val <= 16'b0001100011111010;
            14'h0801 	:	o_val <= 16'b0001100011111101;
            14'h0802 	:	o_val <= 16'b0001100100000000;
            14'h0803 	:	o_val <= 16'b0001100100000011;
            14'h0804 	:	o_val <= 16'b0001100100000110;
            14'h0805 	:	o_val <= 16'b0001100100001001;
            14'h0806 	:	o_val <= 16'b0001100100001100;
            14'h0807 	:	o_val <= 16'b0001100100001111;
            14'h0808 	:	o_val <= 16'b0001100100010010;
            14'h0809 	:	o_val <= 16'b0001100100010101;
            14'h080a 	:	o_val <= 16'b0001100100011001;
            14'h080b 	:	o_val <= 16'b0001100100011100;
            14'h080c 	:	o_val <= 16'b0001100100011111;
            14'h080d 	:	o_val <= 16'b0001100100100010;
            14'h080e 	:	o_val <= 16'b0001100100100101;
            14'h080f 	:	o_val <= 16'b0001100100101000;
            14'h0810 	:	o_val <= 16'b0001100100101011;
            14'h0811 	:	o_val <= 16'b0001100100101110;
            14'h0812 	:	o_val <= 16'b0001100100110001;
            14'h0813 	:	o_val <= 16'b0001100100110100;
            14'h0814 	:	o_val <= 16'b0001100100110111;
            14'h0815 	:	o_val <= 16'b0001100100111010;
            14'h0816 	:	o_val <= 16'b0001100100111110;
            14'h0817 	:	o_val <= 16'b0001100101000001;
            14'h0818 	:	o_val <= 16'b0001100101000100;
            14'h0819 	:	o_val <= 16'b0001100101000111;
            14'h081a 	:	o_val <= 16'b0001100101001010;
            14'h081b 	:	o_val <= 16'b0001100101001101;
            14'h081c 	:	o_val <= 16'b0001100101010000;
            14'h081d 	:	o_val <= 16'b0001100101010011;
            14'h081e 	:	o_val <= 16'b0001100101010110;
            14'h081f 	:	o_val <= 16'b0001100101011001;
            14'h0820 	:	o_val <= 16'b0001100101011100;
            14'h0821 	:	o_val <= 16'b0001100101011111;
            14'h0822 	:	o_val <= 16'b0001100101100010;
            14'h0823 	:	o_val <= 16'b0001100101100110;
            14'h0824 	:	o_val <= 16'b0001100101101001;
            14'h0825 	:	o_val <= 16'b0001100101101100;
            14'h0826 	:	o_val <= 16'b0001100101101111;
            14'h0827 	:	o_val <= 16'b0001100101110010;
            14'h0828 	:	o_val <= 16'b0001100101110101;
            14'h0829 	:	o_val <= 16'b0001100101111000;
            14'h082a 	:	o_val <= 16'b0001100101111011;
            14'h082b 	:	o_val <= 16'b0001100101111110;
            14'h082c 	:	o_val <= 16'b0001100110000001;
            14'h082d 	:	o_val <= 16'b0001100110000100;
            14'h082e 	:	o_val <= 16'b0001100110000111;
            14'h082f 	:	o_val <= 16'b0001100110001011;
            14'h0830 	:	o_val <= 16'b0001100110001110;
            14'h0831 	:	o_val <= 16'b0001100110010001;
            14'h0832 	:	o_val <= 16'b0001100110010100;
            14'h0833 	:	o_val <= 16'b0001100110010111;
            14'h0834 	:	o_val <= 16'b0001100110011010;
            14'h0835 	:	o_val <= 16'b0001100110011101;
            14'h0836 	:	o_val <= 16'b0001100110100000;
            14'h0837 	:	o_val <= 16'b0001100110100011;
            14'h0838 	:	o_val <= 16'b0001100110100110;
            14'h0839 	:	o_val <= 16'b0001100110101001;
            14'h083a 	:	o_val <= 16'b0001100110101100;
            14'h083b 	:	o_val <= 16'b0001100110101111;
            14'h083c 	:	o_val <= 16'b0001100110110011;
            14'h083d 	:	o_val <= 16'b0001100110110110;
            14'h083e 	:	o_val <= 16'b0001100110111001;
            14'h083f 	:	o_val <= 16'b0001100110111100;
            14'h0840 	:	o_val <= 16'b0001100110111111;
            14'h0841 	:	o_val <= 16'b0001100111000010;
            14'h0842 	:	o_val <= 16'b0001100111000101;
            14'h0843 	:	o_val <= 16'b0001100111001000;
            14'h0844 	:	o_val <= 16'b0001100111001011;
            14'h0845 	:	o_val <= 16'b0001100111001110;
            14'h0846 	:	o_val <= 16'b0001100111010001;
            14'h0847 	:	o_val <= 16'b0001100111010100;
            14'h0848 	:	o_val <= 16'b0001100111010111;
            14'h0849 	:	o_val <= 16'b0001100111011011;
            14'h084a 	:	o_val <= 16'b0001100111011110;
            14'h084b 	:	o_val <= 16'b0001100111100001;
            14'h084c 	:	o_val <= 16'b0001100111100100;
            14'h084d 	:	o_val <= 16'b0001100111100111;
            14'h084e 	:	o_val <= 16'b0001100111101010;
            14'h084f 	:	o_val <= 16'b0001100111101101;
            14'h0850 	:	o_val <= 16'b0001100111110000;
            14'h0851 	:	o_val <= 16'b0001100111110011;
            14'h0852 	:	o_val <= 16'b0001100111110110;
            14'h0853 	:	o_val <= 16'b0001100111111001;
            14'h0854 	:	o_val <= 16'b0001100111111100;
            14'h0855 	:	o_val <= 16'b0001100111111111;
            14'h0856 	:	o_val <= 16'b0001101000000011;
            14'h0857 	:	o_val <= 16'b0001101000000110;
            14'h0858 	:	o_val <= 16'b0001101000001001;
            14'h0859 	:	o_val <= 16'b0001101000001100;
            14'h085a 	:	o_val <= 16'b0001101000001111;
            14'h085b 	:	o_val <= 16'b0001101000010010;
            14'h085c 	:	o_val <= 16'b0001101000010101;
            14'h085d 	:	o_val <= 16'b0001101000011000;
            14'h085e 	:	o_val <= 16'b0001101000011011;
            14'h085f 	:	o_val <= 16'b0001101000011110;
            14'h0860 	:	o_val <= 16'b0001101000100001;
            14'h0861 	:	o_val <= 16'b0001101000100100;
            14'h0862 	:	o_val <= 16'b0001101000100111;
            14'h0863 	:	o_val <= 16'b0001101000101011;
            14'h0864 	:	o_val <= 16'b0001101000101110;
            14'h0865 	:	o_val <= 16'b0001101000110001;
            14'h0866 	:	o_val <= 16'b0001101000110100;
            14'h0867 	:	o_val <= 16'b0001101000110111;
            14'h0868 	:	o_val <= 16'b0001101000111010;
            14'h0869 	:	o_val <= 16'b0001101000111101;
            14'h086a 	:	o_val <= 16'b0001101001000000;
            14'h086b 	:	o_val <= 16'b0001101001000011;
            14'h086c 	:	o_val <= 16'b0001101001000110;
            14'h086d 	:	o_val <= 16'b0001101001001001;
            14'h086e 	:	o_val <= 16'b0001101001001100;
            14'h086f 	:	o_val <= 16'b0001101001001111;
            14'h0870 	:	o_val <= 16'b0001101001010010;
            14'h0871 	:	o_val <= 16'b0001101001010110;
            14'h0872 	:	o_val <= 16'b0001101001011001;
            14'h0873 	:	o_val <= 16'b0001101001011100;
            14'h0874 	:	o_val <= 16'b0001101001011111;
            14'h0875 	:	o_val <= 16'b0001101001100010;
            14'h0876 	:	o_val <= 16'b0001101001100101;
            14'h0877 	:	o_val <= 16'b0001101001101000;
            14'h0878 	:	o_val <= 16'b0001101001101011;
            14'h0879 	:	o_val <= 16'b0001101001101110;
            14'h087a 	:	o_val <= 16'b0001101001110001;
            14'h087b 	:	o_val <= 16'b0001101001110100;
            14'h087c 	:	o_val <= 16'b0001101001110111;
            14'h087d 	:	o_val <= 16'b0001101001111010;
            14'h087e 	:	o_val <= 16'b0001101001111110;
            14'h087f 	:	o_val <= 16'b0001101010000001;
            14'h0880 	:	o_val <= 16'b0001101010000100;
            14'h0881 	:	o_val <= 16'b0001101010000111;
            14'h0882 	:	o_val <= 16'b0001101010001010;
            14'h0883 	:	o_val <= 16'b0001101010001101;
            14'h0884 	:	o_val <= 16'b0001101010010000;
            14'h0885 	:	o_val <= 16'b0001101010010011;
            14'h0886 	:	o_val <= 16'b0001101010010110;
            14'h0887 	:	o_val <= 16'b0001101010011001;
            14'h0888 	:	o_val <= 16'b0001101010011100;
            14'h0889 	:	o_val <= 16'b0001101010011111;
            14'h088a 	:	o_val <= 16'b0001101010100010;
            14'h088b 	:	o_val <= 16'b0001101010100101;
            14'h088c 	:	o_val <= 16'b0001101010101001;
            14'h088d 	:	o_val <= 16'b0001101010101100;
            14'h088e 	:	o_val <= 16'b0001101010101111;
            14'h088f 	:	o_val <= 16'b0001101010110010;
            14'h0890 	:	o_val <= 16'b0001101010110101;
            14'h0891 	:	o_val <= 16'b0001101010111000;
            14'h0892 	:	o_val <= 16'b0001101010111011;
            14'h0893 	:	o_val <= 16'b0001101010111110;
            14'h0894 	:	o_val <= 16'b0001101011000001;
            14'h0895 	:	o_val <= 16'b0001101011000100;
            14'h0896 	:	o_val <= 16'b0001101011000111;
            14'h0897 	:	o_val <= 16'b0001101011001010;
            14'h0898 	:	o_val <= 16'b0001101011001101;
            14'h0899 	:	o_val <= 16'b0001101011010000;
            14'h089a 	:	o_val <= 16'b0001101011010100;
            14'h089b 	:	o_val <= 16'b0001101011010111;
            14'h089c 	:	o_val <= 16'b0001101011011010;
            14'h089d 	:	o_val <= 16'b0001101011011101;
            14'h089e 	:	o_val <= 16'b0001101011100000;
            14'h089f 	:	o_val <= 16'b0001101011100011;
            14'h08a0 	:	o_val <= 16'b0001101011100110;
            14'h08a1 	:	o_val <= 16'b0001101011101001;
            14'h08a2 	:	o_val <= 16'b0001101011101100;
            14'h08a3 	:	o_val <= 16'b0001101011101111;
            14'h08a4 	:	o_val <= 16'b0001101011110010;
            14'h08a5 	:	o_val <= 16'b0001101011110101;
            14'h08a6 	:	o_val <= 16'b0001101011111000;
            14'h08a7 	:	o_val <= 16'b0001101011111011;
            14'h08a8 	:	o_val <= 16'b0001101011111111;
            14'h08a9 	:	o_val <= 16'b0001101100000010;
            14'h08aa 	:	o_val <= 16'b0001101100000101;
            14'h08ab 	:	o_val <= 16'b0001101100001000;
            14'h08ac 	:	o_val <= 16'b0001101100001011;
            14'h08ad 	:	o_val <= 16'b0001101100001110;
            14'h08ae 	:	o_val <= 16'b0001101100010001;
            14'h08af 	:	o_val <= 16'b0001101100010100;
            14'h08b0 	:	o_val <= 16'b0001101100010111;
            14'h08b1 	:	o_val <= 16'b0001101100011010;
            14'h08b2 	:	o_val <= 16'b0001101100011101;
            14'h08b3 	:	o_val <= 16'b0001101100100000;
            14'h08b4 	:	o_val <= 16'b0001101100100011;
            14'h08b5 	:	o_val <= 16'b0001101100100110;
            14'h08b6 	:	o_val <= 16'b0001101100101010;
            14'h08b7 	:	o_val <= 16'b0001101100101101;
            14'h08b8 	:	o_val <= 16'b0001101100110000;
            14'h08b9 	:	o_val <= 16'b0001101100110011;
            14'h08ba 	:	o_val <= 16'b0001101100110110;
            14'h08bb 	:	o_val <= 16'b0001101100111001;
            14'h08bc 	:	o_val <= 16'b0001101100111100;
            14'h08bd 	:	o_val <= 16'b0001101100111111;
            14'h08be 	:	o_val <= 16'b0001101101000010;
            14'h08bf 	:	o_val <= 16'b0001101101000101;
            14'h08c0 	:	o_val <= 16'b0001101101001000;
            14'h08c1 	:	o_val <= 16'b0001101101001011;
            14'h08c2 	:	o_val <= 16'b0001101101001110;
            14'h08c3 	:	o_val <= 16'b0001101101010001;
            14'h08c4 	:	o_val <= 16'b0001101101010101;
            14'h08c5 	:	o_val <= 16'b0001101101011000;
            14'h08c6 	:	o_val <= 16'b0001101101011011;
            14'h08c7 	:	o_val <= 16'b0001101101011110;
            14'h08c8 	:	o_val <= 16'b0001101101100001;
            14'h08c9 	:	o_val <= 16'b0001101101100100;
            14'h08ca 	:	o_val <= 16'b0001101101100111;
            14'h08cb 	:	o_val <= 16'b0001101101101010;
            14'h08cc 	:	o_val <= 16'b0001101101101101;
            14'h08cd 	:	o_val <= 16'b0001101101110000;
            14'h08ce 	:	o_val <= 16'b0001101101110011;
            14'h08cf 	:	o_val <= 16'b0001101101110110;
            14'h08d0 	:	o_val <= 16'b0001101101111001;
            14'h08d1 	:	o_val <= 16'b0001101101111100;
            14'h08d2 	:	o_val <= 16'b0001101101111111;
            14'h08d3 	:	o_val <= 16'b0001101110000011;
            14'h08d4 	:	o_val <= 16'b0001101110000110;
            14'h08d5 	:	o_val <= 16'b0001101110001001;
            14'h08d6 	:	o_val <= 16'b0001101110001100;
            14'h08d7 	:	o_val <= 16'b0001101110001111;
            14'h08d8 	:	o_val <= 16'b0001101110010010;
            14'h08d9 	:	o_val <= 16'b0001101110010101;
            14'h08da 	:	o_val <= 16'b0001101110011000;
            14'h08db 	:	o_val <= 16'b0001101110011011;
            14'h08dc 	:	o_val <= 16'b0001101110011110;
            14'h08dd 	:	o_val <= 16'b0001101110100001;
            14'h08de 	:	o_val <= 16'b0001101110100100;
            14'h08df 	:	o_val <= 16'b0001101110100111;
            14'h08e0 	:	o_val <= 16'b0001101110101010;
            14'h08e1 	:	o_val <= 16'b0001101110101101;
            14'h08e2 	:	o_val <= 16'b0001101110110001;
            14'h08e3 	:	o_val <= 16'b0001101110110100;
            14'h08e4 	:	o_val <= 16'b0001101110110111;
            14'h08e5 	:	o_val <= 16'b0001101110111010;
            14'h08e6 	:	o_val <= 16'b0001101110111101;
            14'h08e7 	:	o_val <= 16'b0001101111000000;
            14'h08e8 	:	o_val <= 16'b0001101111000011;
            14'h08e9 	:	o_val <= 16'b0001101111000110;
            14'h08ea 	:	o_val <= 16'b0001101111001001;
            14'h08eb 	:	o_val <= 16'b0001101111001100;
            14'h08ec 	:	o_val <= 16'b0001101111001111;
            14'h08ed 	:	o_val <= 16'b0001101111010010;
            14'h08ee 	:	o_val <= 16'b0001101111010101;
            14'h08ef 	:	o_val <= 16'b0001101111011000;
            14'h08f0 	:	o_val <= 16'b0001101111011011;
            14'h08f1 	:	o_val <= 16'b0001101111011111;
            14'h08f2 	:	o_val <= 16'b0001101111100010;
            14'h08f3 	:	o_val <= 16'b0001101111100101;
            14'h08f4 	:	o_val <= 16'b0001101111101000;
            14'h08f5 	:	o_val <= 16'b0001101111101011;
            14'h08f6 	:	o_val <= 16'b0001101111101110;
            14'h08f7 	:	o_val <= 16'b0001101111110001;
            14'h08f8 	:	o_val <= 16'b0001101111110100;
            14'h08f9 	:	o_val <= 16'b0001101111110111;
            14'h08fa 	:	o_val <= 16'b0001101111111010;
            14'h08fb 	:	o_val <= 16'b0001101111111101;
            14'h08fc 	:	o_val <= 16'b0001110000000000;
            14'h08fd 	:	o_val <= 16'b0001110000000011;
            14'h08fe 	:	o_val <= 16'b0001110000000110;
            14'h08ff 	:	o_val <= 16'b0001110000001001;
            14'h0900 	:	o_val <= 16'b0001110000001101;
            14'h0901 	:	o_val <= 16'b0001110000010000;
            14'h0902 	:	o_val <= 16'b0001110000010011;
            14'h0903 	:	o_val <= 16'b0001110000010110;
            14'h0904 	:	o_val <= 16'b0001110000011001;
            14'h0905 	:	o_val <= 16'b0001110000011100;
            14'h0906 	:	o_val <= 16'b0001110000011111;
            14'h0907 	:	o_val <= 16'b0001110000100010;
            14'h0908 	:	o_val <= 16'b0001110000100101;
            14'h0909 	:	o_val <= 16'b0001110000101000;
            14'h090a 	:	o_val <= 16'b0001110000101011;
            14'h090b 	:	o_val <= 16'b0001110000101110;
            14'h090c 	:	o_val <= 16'b0001110000110001;
            14'h090d 	:	o_val <= 16'b0001110000110100;
            14'h090e 	:	o_val <= 16'b0001110000110111;
            14'h090f 	:	o_val <= 16'b0001110000111011;
            14'h0910 	:	o_val <= 16'b0001110000111110;
            14'h0911 	:	o_val <= 16'b0001110001000001;
            14'h0912 	:	o_val <= 16'b0001110001000100;
            14'h0913 	:	o_val <= 16'b0001110001000111;
            14'h0914 	:	o_val <= 16'b0001110001001010;
            14'h0915 	:	o_val <= 16'b0001110001001101;
            14'h0916 	:	o_val <= 16'b0001110001010000;
            14'h0917 	:	o_val <= 16'b0001110001010011;
            14'h0918 	:	o_val <= 16'b0001110001010110;
            14'h0919 	:	o_val <= 16'b0001110001011001;
            14'h091a 	:	o_val <= 16'b0001110001011100;
            14'h091b 	:	o_val <= 16'b0001110001011111;
            14'h091c 	:	o_val <= 16'b0001110001100010;
            14'h091d 	:	o_val <= 16'b0001110001100101;
            14'h091e 	:	o_val <= 16'b0001110001101000;
            14'h091f 	:	o_val <= 16'b0001110001101100;
            14'h0920 	:	o_val <= 16'b0001110001101111;
            14'h0921 	:	o_val <= 16'b0001110001110010;
            14'h0922 	:	o_val <= 16'b0001110001110101;
            14'h0923 	:	o_val <= 16'b0001110001111000;
            14'h0924 	:	o_val <= 16'b0001110001111011;
            14'h0925 	:	o_val <= 16'b0001110001111110;
            14'h0926 	:	o_val <= 16'b0001110010000001;
            14'h0927 	:	o_val <= 16'b0001110010000100;
            14'h0928 	:	o_val <= 16'b0001110010000111;
            14'h0929 	:	o_val <= 16'b0001110010001010;
            14'h092a 	:	o_val <= 16'b0001110010001101;
            14'h092b 	:	o_val <= 16'b0001110010010000;
            14'h092c 	:	o_val <= 16'b0001110010010011;
            14'h092d 	:	o_val <= 16'b0001110010010110;
            14'h092e 	:	o_val <= 16'b0001110010011001;
            14'h092f 	:	o_val <= 16'b0001110010011101;
            14'h0930 	:	o_val <= 16'b0001110010100000;
            14'h0931 	:	o_val <= 16'b0001110010100011;
            14'h0932 	:	o_val <= 16'b0001110010100110;
            14'h0933 	:	o_val <= 16'b0001110010101001;
            14'h0934 	:	o_val <= 16'b0001110010101100;
            14'h0935 	:	o_val <= 16'b0001110010101111;
            14'h0936 	:	o_val <= 16'b0001110010110010;
            14'h0937 	:	o_val <= 16'b0001110010110101;
            14'h0938 	:	o_val <= 16'b0001110010111000;
            14'h0939 	:	o_val <= 16'b0001110010111011;
            14'h093a 	:	o_val <= 16'b0001110010111110;
            14'h093b 	:	o_val <= 16'b0001110011000001;
            14'h093c 	:	o_val <= 16'b0001110011000100;
            14'h093d 	:	o_val <= 16'b0001110011000111;
            14'h093e 	:	o_val <= 16'b0001110011001010;
            14'h093f 	:	o_val <= 16'b0001110011001110;
            14'h0940 	:	o_val <= 16'b0001110011010001;
            14'h0941 	:	o_val <= 16'b0001110011010100;
            14'h0942 	:	o_val <= 16'b0001110011010111;
            14'h0943 	:	o_val <= 16'b0001110011011010;
            14'h0944 	:	o_val <= 16'b0001110011011101;
            14'h0945 	:	o_val <= 16'b0001110011100000;
            14'h0946 	:	o_val <= 16'b0001110011100011;
            14'h0947 	:	o_val <= 16'b0001110011100110;
            14'h0948 	:	o_val <= 16'b0001110011101001;
            14'h0949 	:	o_val <= 16'b0001110011101100;
            14'h094a 	:	o_val <= 16'b0001110011101111;
            14'h094b 	:	o_val <= 16'b0001110011110010;
            14'h094c 	:	o_val <= 16'b0001110011110101;
            14'h094d 	:	o_val <= 16'b0001110011111000;
            14'h094e 	:	o_val <= 16'b0001110011111011;
            14'h094f 	:	o_val <= 16'b0001110011111110;
            14'h0950 	:	o_val <= 16'b0001110100000010;
            14'h0951 	:	o_val <= 16'b0001110100000101;
            14'h0952 	:	o_val <= 16'b0001110100001000;
            14'h0953 	:	o_val <= 16'b0001110100001011;
            14'h0954 	:	o_val <= 16'b0001110100001110;
            14'h0955 	:	o_val <= 16'b0001110100010001;
            14'h0956 	:	o_val <= 16'b0001110100010100;
            14'h0957 	:	o_val <= 16'b0001110100010111;
            14'h0958 	:	o_val <= 16'b0001110100011010;
            14'h0959 	:	o_val <= 16'b0001110100011101;
            14'h095a 	:	o_val <= 16'b0001110100100000;
            14'h095b 	:	o_val <= 16'b0001110100100011;
            14'h095c 	:	o_val <= 16'b0001110100100110;
            14'h095d 	:	o_val <= 16'b0001110100101001;
            14'h095e 	:	o_val <= 16'b0001110100101100;
            14'h095f 	:	o_val <= 16'b0001110100101111;
            14'h0960 	:	o_val <= 16'b0001110100110010;
            14'h0961 	:	o_val <= 16'b0001110100110110;
            14'h0962 	:	o_val <= 16'b0001110100111001;
            14'h0963 	:	o_val <= 16'b0001110100111100;
            14'h0964 	:	o_val <= 16'b0001110100111111;
            14'h0965 	:	o_val <= 16'b0001110101000010;
            14'h0966 	:	o_val <= 16'b0001110101000101;
            14'h0967 	:	o_val <= 16'b0001110101001000;
            14'h0968 	:	o_val <= 16'b0001110101001011;
            14'h0969 	:	o_val <= 16'b0001110101001110;
            14'h096a 	:	o_val <= 16'b0001110101010001;
            14'h096b 	:	o_val <= 16'b0001110101010100;
            14'h096c 	:	o_val <= 16'b0001110101010111;
            14'h096d 	:	o_val <= 16'b0001110101011010;
            14'h096e 	:	o_val <= 16'b0001110101011101;
            14'h096f 	:	o_val <= 16'b0001110101100000;
            14'h0970 	:	o_val <= 16'b0001110101100011;
            14'h0971 	:	o_val <= 16'b0001110101100110;
            14'h0972 	:	o_val <= 16'b0001110101101010;
            14'h0973 	:	o_val <= 16'b0001110101101101;
            14'h0974 	:	o_val <= 16'b0001110101110000;
            14'h0975 	:	o_val <= 16'b0001110101110011;
            14'h0976 	:	o_val <= 16'b0001110101110110;
            14'h0977 	:	o_val <= 16'b0001110101111001;
            14'h0978 	:	o_val <= 16'b0001110101111100;
            14'h0979 	:	o_val <= 16'b0001110101111111;
            14'h097a 	:	o_val <= 16'b0001110110000010;
            14'h097b 	:	o_val <= 16'b0001110110000101;
            14'h097c 	:	o_val <= 16'b0001110110001000;
            14'h097d 	:	o_val <= 16'b0001110110001011;
            14'h097e 	:	o_val <= 16'b0001110110001110;
            14'h097f 	:	o_val <= 16'b0001110110010001;
            14'h0980 	:	o_val <= 16'b0001110110010100;
            14'h0981 	:	o_val <= 16'b0001110110010111;
            14'h0982 	:	o_val <= 16'b0001110110011010;
            14'h0983 	:	o_val <= 16'b0001110110011110;
            14'h0984 	:	o_val <= 16'b0001110110100001;
            14'h0985 	:	o_val <= 16'b0001110110100100;
            14'h0986 	:	o_val <= 16'b0001110110100111;
            14'h0987 	:	o_val <= 16'b0001110110101010;
            14'h0988 	:	o_val <= 16'b0001110110101101;
            14'h0989 	:	o_val <= 16'b0001110110110000;
            14'h098a 	:	o_val <= 16'b0001110110110011;
            14'h098b 	:	o_val <= 16'b0001110110110110;
            14'h098c 	:	o_val <= 16'b0001110110111001;
            14'h098d 	:	o_val <= 16'b0001110110111100;
            14'h098e 	:	o_val <= 16'b0001110110111111;
            14'h098f 	:	o_val <= 16'b0001110111000010;
            14'h0990 	:	o_val <= 16'b0001110111000101;
            14'h0991 	:	o_val <= 16'b0001110111001000;
            14'h0992 	:	o_val <= 16'b0001110111001011;
            14'h0993 	:	o_val <= 16'b0001110111001110;
            14'h0994 	:	o_val <= 16'b0001110111010001;
            14'h0995 	:	o_val <= 16'b0001110111010101;
            14'h0996 	:	o_val <= 16'b0001110111011000;
            14'h0997 	:	o_val <= 16'b0001110111011011;
            14'h0998 	:	o_val <= 16'b0001110111011110;
            14'h0999 	:	o_val <= 16'b0001110111100001;
            14'h099a 	:	o_val <= 16'b0001110111100100;
            14'h099b 	:	o_val <= 16'b0001110111100111;
            14'h099c 	:	o_val <= 16'b0001110111101010;
            14'h099d 	:	o_val <= 16'b0001110111101101;
            14'h099e 	:	o_val <= 16'b0001110111110000;
            14'h099f 	:	o_val <= 16'b0001110111110011;
            14'h09a0 	:	o_val <= 16'b0001110111110110;
            14'h09a1 	:	o_val <= 16'b0001110111111001;
            14'h09a2 	:	o_val <= 16'b0001110111111100;
            14'h09a3 	:	o_val <= 16'b0001110111111111;
            14'h09a4 	:	o_val <= 16'b0001111000000010;
            14'h09a5 	:	o_val <= 16'b0001111000000101;
            14'h09a6 	:	o_val <= 16'b0001111000001000;
            14'h09a7 	:	o_val <= 16'b0001111000001011;
            14'h09a8 	:	o_val <= 16'b0001111000001111;
            14'h09a9 	:	o_val <= 16'b0001111000010010;
            14'h09aa 	:	o_val <= 16'b0001111000010101;
            14'h09ab 	:	o_val <= 16'b0001111000011000;
            14'h09ac 	:	o_val <= 16'b0001111000011011;
            14'h09ad 	:	o_val <= 16'b0001111000011110;
            14'h09ae 	:	o_val <= 16'b0001111000100001;
            14'h09af 	:	o_val <= 16'b0001111000100100;
            14'h09b0 	:	o_val <= 16'b0001111000100111;
            14'h09b1 	:	o_val <= 16'b0001111000101010;
            14'h09b2 	:	o_val <= 16'b0001111000101101;
            14'h09b3 	:	o_val <= 16'b0001111000110000;
            14'h09b4 	:	o_val <= 16'b0001111000110011;
            14'h09b5 	:	o_val <= 16'b0001111000110110;
            14'h09b6 	:	o_val <= 16'b0001111000111001;
            14'h09b7 	:	o_val <= 16'b0001111000111100;
            14'h09b8 	:	o_val <= 16'b0001111000111111;
            14'h09b9 	:	o_val <= 16'b0001111001000010;
            14'h09ba 	:	o_val <= 16'b0001111001000110;
            14'h09bb 	:	o_val <= 16'b0001111001001001;
            14'h09bc 	:	o_val <= 16'b0001111001001100;
            14'h09bd 	:	o_val <= 16'b0001111001001111;
            14'h09be 	:	o_val <= 16'b0001111001010010;
            14'h09bf 	:	o_val <= 16'b0001111001010101;
            14'h09c0 	:	o_val <= 16'b0001111001011000;
            14'h09c1 	:	o_val <= 16'b0001111001011011;
            14'h09c2 	:	o_val <= 16'b0001111001011110;
            14'h09c3 	:	o_val <= 16'b0001111001100001;
            14'h09c4 	:	o_val <= 16'b0001111001100100;
            14'h09c5 	:	o_val <= 16'b0001111001100111;
            14'h09c6 	:	o_val <= 16'b0001111001101010;
            14'h09c7 	:	o_val <= 16'b0001111001101101;
            14'h09c8 	:	o_val <= 16'b0001111001110000;
            14'h09c9 	:	o_val <= 16'b0001111001110011;
            14'h09ca 	:	o_val <= 16'b0001111001110110;
            14'h09cb 	:	o_val <= 16'b0001111001111001;
            14'h09cc 	:	o_val <= 16'b0001111001111100;
            14'h09cd 	:	o_val <= 16'b0001111001111111;
            14'h09ce 	:	o_val <= 16'b0001111010000011;
            14'h09cf 	:	o_val <= 16'b0001111010000110;
            14'h09d0 	:	o_val <= 16'b0001111010001001;
            14'h09d1 	:	o_val <= 16'b0001111010001100;
            14'h09d2 	:	o_val <= 16'b0001111010001111;
            14'h09d3 	:	o_val <= 16'b0001111010010010;
            14'h09d4 	:	o_val <= 16'b0001111010010101;
            14'h09d5 	:	o_val <= 16'b0001111010011000;
            14'h09d6 	:	o_val <= 16'b0001111010011011;
            14'h09d7 	:	o_val <= 16'b0001111010011110;
            14'h09d8 	:	o_val <= 16'b0001111010100001;
            14'h09d9 	:	o_val <= 16'b0001111010100100;
            14'h09da 	:	o_val <= 16'b0001111010100111;
            14'h09db 	:	o_val <= 16'b0001111010101010;
            14'h09dc 	:	o_val <= 16'b0001111010101101;
            14'h09dd 	:	o_val <= 16'b0001111010110000;
            14'h09de 	:	o_val <= 16'b0001111010110011;
            14'h09df 	:	o_val <= 16'b0001111010110110;
            14'h09e0 	:	o_val <= 16'b0001111010111001;
            14'h09e1 	:	o_val <= 16'b0001111010111100;
            14'h09e2 	:	o_val <= 16'b0001111011000000;
            14'h09e3 	:	o_val <= 16'b0001111011000011;
            14'h09e4 	:	o_val <= 16'b0001111011000110;
            14'h09e5 	:	o_val <= 16'b0001111011001001;
            14'h09e6 	:	o_val <= 16'b0001111011001100;
            14'h09e7 	:	o_val <= 16'b0001111011001111;
            14'h09e8 	:	o_val <= 16'b0001111011010010;
            14'h09e9 	:	o_val <= 16'b0001111011010101;
            14'h09ea 	:	o_val <= 16'b0001111011011000;
            14'h09eb 	:	o_val <= 16'b0001111011011011;
            14'h09ec 	:	o_val <= 16'b0001111011011110;
            14'h09ed 	:	o_val <= 16'b0001111011100001;
            14'h09ee 	:	o_val <= 16'b0001111011100100;
            14'h09ef 	:	o_val <= 16'b0001111011100111;
            14'h09f0 	:	o_val <= 16'b0001111011101010;
            14'h09f1 	:	o_val <= 16'b0001111011101101;
            14'h09f2 	:	o_val <= 16'b0001111011110000;
            14'h09f3 	:	o_val <= 16'b0001111011110011;
            14'h09f4 	:	o_val <= 16'b0001111011110110;
            14'h09f5 	:	o_val <= 16'b0001111011111001;
            14'h09f6 	:	o_val <= 16'b0001111011111101;
            14'h09f7 	:	o_val <= 16'b0001111100000000;
            14'h09f8 	:	o_val <= 16'b0001111100000011;
            14'h09f9 	:	o_val <= 16'b0001111100000110;
            14'h09fa 	:	o_val <= 16'b0001111100001001;
            14'h09fb 	:	o_val <= 16'b0001111100001100;
            14'h09fc 	:	o_val <= 16'b0001111100001111;
            14'h09fd 	:	o_val <= 16'b0001111100010010;
            14'h09fe 	:	o_val <= 16'b0001111100010101;
            14'h09ff 	:	o_val <= 16'b0001111100011000;
            14'h0a00 	:	o_val <= 16'b0001111100011011;
            14'h0a01 	:	o_val <= 16'b0001111100011110;
            14'h0a02 	:	o_val <= 16'b0001111100100001;
            14'h0a03 	:	o_val <= 16'b0001111100100100;
            14'h0a04 	:	o_val <= 16'b0001111100100111;
            14'h0a05 	:	o_val <= 16'b0001111100101010;
            14'h0a06 	:	o_val <= 16'b0001111100101101;
            14'h0a07 	:	o_val <= 16'b0001111100110000;
            14'h0a08 	:	o_val <= 16'b0001111100110011;
            14'h0a09 	:	o_val <= 16'b0001111100110110;
            14'h0a0a 	:	o_val <= 16'b0001111100111001;
            14'h0a0b 	:	o_val <= 16'b0001111100111101;
            14'h0a0c 	:	o_val <= 16'b0001111101000000;
            14'h0a0d 	:	o_val <= 16'b0001111101000011;
            14'h0a0e 	:	o_val <= 16'b0001111101000110;
            14'h0a0f 	:	o_val <= 16'b0001111101001001;
            14'h0a10 	:	o_val <= 16'b0001111101001100;
            14'h0a11 	:	o_val <= 16'b0001111101001111;
            14'h0a12 	:	o_val <= 16'b0001111101010010;
            14'h0a13 	:	o_val <= 16'b0001111101010101;
            14'h0a14 	:	o_val <= 16'b0001111101011000;
            14'h0a15 	:	o_val <= 16'b0001111101011011;
            14'h0a16 	:	o_val <= 16'b0001111101011110;
            14'h0a17 	:	o_val <= 16'b0001111101100001;
            14'h0a18 	:	o_val <= 16'b0001111101100100;
            14'h0a19 	:	o_val <= 16'b0001111101100111;
            14'h0a1a 	:	o_val <= 16'b0001111101101010;
            14'h0a1b 	:	o_val <= 16'b0001111101101101;
            14'h0a1c 	:	o_val <= 16'b0001111101110000;
            14'h0a1d 	:	o_val <= 16'b0001111101110011;
            14'h0a1e 	:	o_val <= 16'b0001111101110110;
            14'h0a1f 	:	o_val <= 16'b0001111101111001;
            14'h0a20 	:	o_val <= 16'b0001111101111100;
            14'h0a21 	:	o_val <= 16'b0001111110000000;
            14'h0a22 	:	o_val <= 16'b0001111110000011;
            14'h0a23 	:	o_val <= 16'b0001111110000110;
            14'h0a24 	:	o_val <= 16'b0001111110001001;
            14'h0a25 	:	o_val <= 16'b0001111110001100;
            14'h0a26 	:	o_val <= 16'b0001111110001111;
            14'h0a27 	:	o_val <= 16'b0001111110010010;
            14'h0a28 	:	o_val <= 16'b0001111110010101;
            14'h0a29 	:	o_val <= 16'b0001111110011000;
            14'h0a2a 	:	o_val <= 16'b0001111110011011;
            14'h0a2b 	:	o_val <= 16'b0001111110011110;
            14'h0a2c 	:	o_val <= 16'b0001111110100001;
            14'h0a2d 	:	o_val <= 16'b0001111110100100;
            14'h0a2e 	:	o_val <= 16'b0001111110100111;
            14'h0a2f 	:	o_val <= 16'b0001111110101010;
            14'h0a30 	:	o_val <= 16'b0001111110101101;
            14'h0a31 	:	o_val <= 16'b0001111110110000;
            14'h0a32 	:	o_val <= 16'b0001111110110011;
            14'h0a33 	:	o_val <= 16'b0001111110110110;
            14'h0a34 	:	o_val <= 16'b0001111110111001;
            14'h0a35 	:	o_val <= 16'b0001111110111100;
            14'h0a36 	:	o_val <= 16'b0001111110111111;
            14'h0a37 	:	o_val <= 16'b0001111111000010;
            14'h0a38 	:	o_val <= 16'b0001111111000110;
            14'h0a39 	:	o_val <= 16'b0001111111001001;
            14'h0a3a 	:	o_val <= 16'b0001111111001100;
            14'h0a3b 	:	o_val <= 16'b0001111111001111;
            14'h0a3c 	:	o_val <= 16'b0001111111010010;
            14'h0a3d 	:	o_val <= 16'b0001111111010101;
            14'h0a3e 	:	o_val <= 16'b0001111111011000;
            14'h0a3f 	:	o_val <= 16'b0001111111011011;
            14'h0a40 	:	o_val <= 16'b0001111111011110;
            14'h0a41 	:	o_val <= 16'b0001111111100001;
            14'h0a42 	:	o_val <= 16'b0001111111100100;
            14'h0a43 	:	o_val <= 16'b0001111111100111;
            14'h0a44 	:	o_val <= 16'b0001111111101010;
            14'h0a45 	:	o_val <= 16'b0001111111101101;
            14'h0a46 	:	o_val <= 16'b0001111111110000;
            14'h0a47 	:	o_val <= 16'b0001111111110011;
            14'h0a48 	:	o_val <= 16'b0001111111110110;
            14'h0a49 	:	o_val <= 16'b0001111111111001;
            14'h0a4a 	:	o_val <= 16'b0001111111111100;
            14'h0a4b 	:	o_val <= 16'b0001111111111111;
            14'h0a4c 	:	o_val <= 16'b0010000000000010;
            14'h0a4d 	:	o_val <= 16'b0010000000000101;
            14'h0a4e 	:	o_val <= 16'b0010000000001000;
            14'h0a4f 	:	o_val <= 16'b0010000000001100;
            14'h0a50 	:	o_val <= 16'b0010000000001111;
            14'h0a51 	:	o_val <= 16'b0010000000010010;
            14'h0a52 	:	o_val <= 16'b0010000000010101;
            14'h0a53 	:	o_val <= 16'b0010000000011000;
            14'h0a54 	:	o_val <= 16'b0010000000011011;
            14'h0a55 	:	o_val <= 16'b0010000000011110;
            14'h0a56 	:	o_val <= 16'b0010000000100001;
            14'h0a57 	:	o_val <= 16'b0010000000100100;
            14'h0a58 	:	o_val <= 16'b0010000000100111;
            14'h0a59 	:	o_val <= 16'b0010000000101010;
            14'h0a5a 	:	o_val <= 16'b0010000000101101;
            14'h0a5b 	:	o_val <= 16'b0010000000110000;
            14'h0a5c 	:	o_val <= 16'b0010000000110011;
            14'h0a5d 	:	o_val <= 16'b0010000000110110;
            14'h0a5e 	:	o_val <= 16'b0010000000111001;
            14'h0a5f 	:	o_val <= 16'b0010000000111100;
            14'h0a60 	:	o_val <= 16'b0010000000111111;
            14'h0a61 	:	o_val <= 16'b0010000001000010;
            14'h0a62 	:	o_val <= 16'b0010000001000101;
            14'h0a63 	:	o_val <= 16'b0010000001001000;
            14'h0a64 	:	o_val <= 16'b0010000001001011;
            14'h0a65 	:	o_val <= 16'b0010000001001110;
            14'h0a66 	:	o_val <= 16'b0010000001010001;
            14'h0a67 	:	o_val <= 16'b0010000001010100;
            14'h0a68 	:	o_val <= 16'b0010000001011000;
            14'h0a69 	:	o_val <= 16'b0010000001011011;
            14'h0a6a 	:	o_val <= 16'b0010000001011110;
            14'h0a6b 	:	o_val <= 16'b0010000001100001;
            14'h0a6c 	:	o_val <= 16'b0010000001100100;
            14'h0a6d 	:	o_val <= 16'b0010000001100111;
            14'h0a6e 	:	o_val <= 16'b0010000001101010;
            14'h0a6f 	:	o_val <= 16'b0010000001101101;
            14'h0a70 	:	o_val <= 16'b0010000001110000;
            14'h0a71 	:	o_val <= 16'b0010000001110011;
            14'h0a72 	:	o_val <= 16'b0010000001110110;
            14'h0a73 	:	o_val <= 16'b0010000001111001;
            14'h0a74 	:	o_val <= 16'b0010000001111100;
            14'h0a75 	:	o_val <= 16'b0010000001111111;
            14'h0a76 	:	o_val <= 16'b0010000010000010;
            14'h0a77 	:	o_val <= 16'b0010000010000101;
            14'h0a78 	:	o_val <= 16'b0010000010001000;
            14'h0a79 	:	o_val <= 16'b0010000010001011;
            14'h0a7a 	:	o_val <= 16'b0010000010001110;
            14'h0a7b 	:	o_val <= 16'b0010000010010001;
            14'h0a7c 	:	o_val <= 16'b0010000010010100;
            14'h0a7d 	:	o_val <= 16'b0010000010010111;
            14'h0a7e 	:	o_val <= 16'b0010000010011010;
            14'h0a7f 	:	o_val <= 16'b0010000010011101;
            14'h0a80 	:	o_val <= 16'b0010000010100000;
            14'h0a81 	:	o_val <= 16'b0010000010100011;
            14'h0a82 	:	o_val <= 16'b0010000010100111;
            14'h0a83 	:	o_val <= 16'b0010000010101010;
            14'h0a84 	:	o_val <= 16'b0010000010101101;
            14'h0a85 	:	o_val <= 16'b0010000010110000;
            14'h0a86 	:	o_val <= 16'b0010000010110011;
            14'h0a87 	:	o_val <= 16'b0010000010110110;
            14'h0a88 	:	o_val <= 16'b0010000010111001;
            14'h0a89 	:	o_val <= 16'b0010000010111100;
            14'h0a8a 	:	o_val <= 16'b0010000010111111;
            14'h0a8b 	:	o_val <= 16'b0010000011000010;
            14'h0a8c 	:	o_val <= 16'b0010000011000101;
            14'h0a8d 	:	o_val <= 16'b0010000011001000;
            14'h0a8e 	:	o_val <= 16'b0010000011001011;
            14'h0a8f 	:	o_val <= 16'b0010000011001110;
            14'h0a90 	:	o_val <= 16'b0010000011010001;
            14'h0a91 	:	o_val <= 16'b0010000011010100;
            14'h0a92 	:	o_val <= 16'b0010000011010111;
            14'h0a93 	:	o_val <= 16'b0010000011011010;
            14'h0a94 	:	o_val <= 16'b0010000011011101;
            14'h0a95 	:	o_val <= 16'b0010000011100000;
            14'h0a96 	:	o_val <= 16'b0010000011100011;
            14'h0a97 	:	o_val <= 16'b0010000011100110;
            14'h0a98 	:	o_val <= 16'b0010000011101001;
            14'h0a99 	:	o_val <= 16'b0010000011101100;
            14'h0a9a 	:	o_val <= 16'b0010000011101111;
            14'h0a9b 	:	o_val <= 16'b0010000011110010;
            14'h0a9c 	:	o_val <= 16'b0010000011110101;
            14'h0a9d 	:	o_val <= 16'b0010000011111001;
            14'h0a9e 	:	o_val <= 16'b0010000011111100;
            14'h0a9f 	:	o_val <= 16'b0010000011111111;
            14'h0aa0 	:	o_val <= 16'b0010000100000010;
            14'h0aa1 	:	o_val <= 16'b0010000100000101;
            14'h0aa2 	:	o_val <= 16'b0010000100001000;
            14'h0aa3 	:	o_val <= 16'b0010000100001011;
            14'h0aa4 	:	o_val <= 16'b0010000100001110;
            14'h0aa5 	:	o_val <= 16'b0010000100010001;
            14'h0aa6 	:	o_val <= 16'b0010000100010100;
            14'h0aa7 	:	o_val <= 16'b0010000100010111;
            14'h0aa8 	:	o_val <= 16'b0010000100011010;
            14'h0aa9 	:	o_val <= 16'b0010000100011101;
            14'h0aaa 	:	o_val <= 16'b0010000100100000;
            14'h0aab 	:	o_val <= 16'b0010000100100011;
            14'h0aac 	:	o_val <= 16'b0010000100100110;
            14'h0aad 	:	o_val <= 16'b0010000100101001;
            14'h0aae 	:	o_val <= 16'b0010000100101100;
            14'h0aaf 	:	o_val <= 16'b0010000100101111;
            14'h0ab0 	:	o_val <= 16'b0010000100110010;
            14'h0ab1 	:	o_val <= 16'b0010000100110101;
            14'h0ab2 	:	o_val <= 16'b0010000100111000;
            14'h0ab3 	:	o_val <= 16'b0010000100111011;
            14'h0ab4 	:	o_val <= 16'b0010000100111110;
            14'h0ab5 	:	o_val <= 16'b0010000101000001;
            14'h0ab6 	:	o_val <= 16'b0010000101000100;
            14'h0ab7 	:	o_val <= 16'b0010000101000111;
            14'h0ab8 	:	o_val <= 16'b0010000101001010;
            14'h0ab9 	:	o_val <= 16'b0010000101001101;
            14'h0aba 	:	o_val <= 16'b0010000101010001;
            14'h0abb 	:	o_val <= 16'b0010000101010100;
            14'h0abc 	:	o_val <= 16'b0010000101010111;
            14'h0abd 	:	o_val <= 16'b0010000101011010;
            14'h0abe 	:	o_val <= 16'b0010000101011101;
            14'h0abf 	:	o_val <= 16'b0010000101100000;
            14'h0ac0 	:	o_val <= 16'b0010000101100011;
            14'h0ac1 	:	o_val <= 16'b0010000101100110;
            14'h0ac2 	:	o_val <= 16'b0010000101101001;
            14'h0ac3 	:	o_val <= 16'b0010000101101100;
            14'h0ac4 	:	o_val <= 16'b0010000101101111;
            14'h0ac5 	:	o_val <= 16'b0010000101110010;
            14'h0ac6 	:	o_val <= 16'b0010000101110101;
            14'h0ac7 	:	o_val <= 16'b0010000101111000;
            14'h0ac8 	:	o_val <= 16'b0010000101111011;
            14'h0ac9 	:	o_val <= 16'b0010000101111110;
            14'h0aca 	:	o_val <= 16'b0010000110000001;
            14'h0acb 	:	o_val <= 16'b0010000110000100;
            14'h0acc 	:	o_val <= 16'b0010000110000111;
            14'h0acd 	:	o_val <= 16'b0010000110001010;
            14'h0ace 	:	o_val <= 16'b0010000110001101;
            14'h0acf 	:	o_val <= 16'b0010000110010000;
            14'h0ad0 	:	o_val <= 16'b0010000110010011;
            14'h0ad1 	:	o_val <= 16'b0010000110010110;
            14'h0ad2 	:	o_val <= 16'b0010000110011001;
            14'h0ad3 	:	o_val <= 16'b0010000110011100;
            14'h0ad4 	:	o_val <= 16'b0010000110011111;
            14'h0ad5 	:	o_val <= 16'b0010000110100010;
            14'h0ad6 	:	o_val <= 16'b0010000110100101;
            14'h0ad7 	:	o_val <= 16'b0010000110101000;
            14'h0ad8 	:	o_val <= 16'b0010000110101011;
            14'h0ad9 	:	o_val <= 16'b0010000110101111;
            14'h0ada 	:	o_val <= 16'b0010000110110010;
            14'h0adb 	:	o_val <= 16'b0010000110110101;
            14'h0adc 	:	o_val <= 16'b0010000110111000;
            14'h0add 	:	o_val <= 16'b0010000110111011;
            14'h0ade 	:	o_val <= 16'b0010000110111110;
            14'h0adf 	:	o_val <= 16'b0010000111000001;
            14'h0ae0 	:	o_val <= 16'b0010000111000100;
            14'h0ae1 	:	o_val <= 16'b0010000111000111;
            14'h0ae2 	:	o_val <= 16'b0010000111001010;
            14'h0ae3 	:	o_val <= 16'b0010000111001101;
            14'h0ae4 	:	o_val <= 16'b0010000111010000;
            14'h0ae5 	:	o_val <= 16'b0010000111010011;
            14'h0ae6 	:	o_val <= 16'b0010000111010110;
            14'h0ae7 	:	o_val <= 16'b0010000111011001;
            14'h0ae8 	:	o_val <= 16'b0010000111011100;
            14'h0ae9 	:	o_val <= 16'b0010000111011111;
            14'h0aea 	:	o_val <= 16'b0010000111100010;
            14'h0aeb 	:	o_val <= 16'b0010000111100101;
            14'h0aec 	:	o_val <= 16'b0010000111101000;
            14'h0aed 	:	o_val <= 16'b0010000111101011;
            14'h0aee 	:	o_val <= 16'b0010000111101110;
            14'h0aef 	:	o_val <= 16'b0010000111110001;
            14'h0af0 	:	o_val <= 16'b0010000111110100;
            14'h0af1 	:	o_val <= 16'b0010000111110111;
            14'h0af2 	:	o_val <= 16'b0010000111111010;
            14'h0af3 	:	o_val <= 16'b0010000111111101;
            14'h0af4 	:	o_val <= 16'b0010001000000000;
            14'h0af5 	:	o_val <= 16'b0010001000000011;
            14'h0af6 	:	o_val <= 16'b0010001000000110;
            14'h0af7 	:	o_val <= 16'b0010001000001001;
            14'h0af8 	:	o_val <= 16'b0010001000001100;
            14'h0af9 	:	o_val <= 16'b0010001000001111;
            14'h0afa 	:	o_val <= 16'b0010001000010010;
            14'h0afb 	:	o_val <= 16'b0010001000010110;
            14'h0afc 	:	o_val <= 16'b0010001000011001;
            14'h0afd 	:	o_val <= 16'b0010001000011100;
            14'h0afe 	:	o_val <= 16'b0010001000011111;
            14'h0aff 	:	o_val <= 16'b0010001000100010;
            14'h0b00 	:	o_val <= 16'b0010001000100101;
            14'h0b01 	:	o_val <= 16'b0010001000101000;
            14'h0b02 	:	o_val <= 16'b0010001000101011;
            14'h0b03 	:	o_val <= 16'b0010001000101110;
            14'h0b04 	:	o_val <= 16'b0010001000110001;
            14'h0b05 	:	o_val <= 16'b0010001000110100;
            14'h0b06 	:	o_val <= 16'b0010001000110111;
            14'h0b07 	:	o_val <= 16'b0010001000111010;
            14'h0b08 	:	o_val <= 16'b0010001000111101;
            14'h0b09 	:	o_val <= 16'b0010001001000000;
            14'h0b0a 	:	o_val <= 16'b0010001001000011;
            14'h0b0b 	:	o_val <= 16'b0010001001000110;
            14'h0b0c 	:	o_val <= 16'b0010001001001001;
            14'h0b0d 	:	o_val <= 16'b0010001001001100;
            14'h0b0e 	:	o_val <= 16'b0010001001001111;
            14'h0b0f 	:	o_val <= 16'b0010001001010010;
            14'h0b10 	:	o_val <= 16'b0010001001010101;
            14'h0b11 	:	o_val <= 16'b0010001001011000;
            14'h0b12 	:	o_val <= 16'b0010001001011011;
            14'h0b13 	:	o_val <= 16'b0010001001011110;
            14'h0b14 	:	o_val <= 16'b0010001001100001;
            14'h0b15 	:	o_val <= 16'b0010001001100100;
            14'h0b16 	:	o_val <= 16'b0010001001100111;
            14'h0b17 	:	o_val <= 16'b0010001001101010;
            14'h0b18 	:	o_val <= 16'b0010001001101101;
            14'h0b19 	:	o_val <= 16'b0010001001110000;
            14'h0b1a 	:	o_val <= 16'b0010001001110011;
            14'h0b1b 	:	o_val <= 16'b0010001001110110;
            14'h0b1c 	:	o_val <= 16'b0010001001111001;
            14'h0b1d 	:	o_val <= 16'b0010001001111100;
            14'h0b1e 	:	o_val <= 16'b0010001001111111;
            14'h0b1f 	:	o_val <= 16'b0010001010000010;
            14'h0b20 	:	o_val <= 16'b0010001010000110;
            14'h0b21 	:	o_val <= 16'b0010001010001001;
            14'h0b22 	:	o_val <= 16'b0010001010001100;
            14'h0b23 	:	o_val <= 16'b0010001010001111;
            14'h0b24 	:	o_val <= 16'b0010001010010010;
            14'h0b25 	:	o_val <= 16'b0010001010010101;
            14'h0b26 	:	o_val <= 16'b0010001010011000;
            14'h0b27 	:	o_val <= 16'b0010001010011011;
            14'h0b28 	:	o_val <= 16'b0010001010011110;
            14'h0b29 	:	o_val <= 16'b0010001010100001;
            14'h0b2a 	:	o_val <= 16'b0010001010100100;
            14'h0b2b 	:	o_val <= 16'b0010001010100111;
            14'h0b2c 	:	o_val <= 16'b0010001010101010;
            14'h0b2d 	:	o_val <= 16'b0010001010101101;
            14'h0b2e 	:	o_val <= 16'b0010001010110000;
            14'h0b2f 	:	o_val <= 16'b0010001010110011;
            14'h0b30 	:	o_val <= 16'b0010001010110110;
            14'h0b31 	:	o_val <= 16'b0010001010111001;
            14'h0b32 	:	o_val <= 16'b0010001010111100;
            14'h0b33 	:	o_val <= 16'b0010001010111111;
            14'h0b34 	:	o_val <= 16'b0010001011000010;
            14'h0b35 	:	o_val <= 16'b0010001011000101;
            14'h0b36 	:	o_val <= 16'b0010001011001000;
            14'h0b37 	:	o_val <= 16'b0010001011001011;
            14'h0b38 	:	o_val <= 16'b0010001011001110;
            14'h0b39 	:	o_val <= 16'b0010001011010001;
            14'h0b3a 	:	o_val <= 16'b0010001011010100;
            14'h0b3b 	:	o_val <= 16'b0010001011010111;
            14'h0b3c 	:	o_val <= 16'b0010001011011010;
            14'h0b3d 	:	o_val <= 16'b0010001011011101;
            14'h0b3e 	:	o_val <= 16'b0010001011100000;
            14'h0b3f 	:	o_val <= 16'b0010001011100011;
            14'h0b40 	:	o_val <= 16'b0010001011100110;
            14'h0b41 	:	o_val <= 16'b0010001011101001;
            14'h0b42 	:	o_val <= 16'b0010001011101100;
            14'h0b43 	:	o_val <= 16'b0010001011101111;
            14'h0b44 	:	o_val <= 16'b0010001011110010;
            14'h0b45 	:	o_val <= 16'b0010001011110101;
            14'h0b46 	:	o_val <= 16'b0010001011111000;
            14'h0b47 	:	o_val <= 16'b0010001011111011;
            14'h0b48 	:	o_val <= 16'b0010001011111110;
            14'h0b49 	:	o_val <= 16'b0010001100000001;
            14'h0b4a 	:	o_val <= 16'b0010001100000100;
            14'h0b4b 	:	o_val <= 16'b0010001100001000;
            14'h0b4c 	:	o_val <= 16'b0010001100001011;
            14'h0b4d 	:	o_val <= 16'b0010001100001110;
            14'h0b4e 	:	o_val <= 16'b0010001100010001;
            14'h0b4f 	:	o_val <= 16'b0010001100010100;
            14'h0b50 	:	o_val <= 16'b0010001100010111;
            14'h0b51 	:	o_val <= 16'b0010001100011010;
            14'h0b52 	:	o_val <= 16'b0010001100011101;
            14'h0b53 	:	o_val <= 16'b0010001100100000;
            14'h0b54 	:	o_val <= 16'b0010001100100011;
            14'h0b55 	:	o_val <= 16'b0010001100100110;
            14'h0b56 	:	o_val <= 16'b0010001100101001;
            14'h0b57 	:	o_val <= 16'b0010001100101100;
            14'h0b58 	:	o_val <= 16'b0010001100101111;
            14'h0b59 	:	o_val <= 16'b0010001100110010;
            14'h0b5a 	:	o_val <= 16'b0010001100110101;
            14'h0b5b 	:	o_val <= 16'b0010001100111000;
            14'h0b5c 	:	o_val <= 16'b0010001100111011;
            14'h0b5d 	:	o_val <= 16'b0010001100111110;
            14'h0b5e 	:	o_val <= 16'b0010001101000001;
            14'h0b5f 	:	o_val <= 16'b0010001101000100;
            14'h0b60 	:	o_val <= 16'b0010001101000111;
            14'h0b61 	:	o_val <= 16'b0010001101001010;
            14'h0b62 	:	o_val <= 16'b0010001101001101;
            14'h0b63 	:	o_val <= 16'b0010001101010000;
            14'h0b64 	:	o_val <= 16'b0010001101010011;
            14'h0b65 	:	o_val <= 16'b0010001101010110;
            14'h0b66 	:	o_val <= 16'b0010001101011001;
            14'h0b67 	:	o_val <= 16'b0010001101011100;
            14'h0b68 	:	o_val <= 16'b0010001101011111;
            14'h0b69 	:	o_val <= 16'b0010001101100010;
            14'h0b6a 	:	o_val <= 16'b0010001101100101;
            14'h0b6b 	:	o_val <= 16'b0010001101101000;
            14'h0b6c 	:	o_val <= 16'b0010001101101011;
            14'h0b6d 	:	o_val <= 16'b0010001101101110;
            14'h0b6e 	:	o_val <= 16'b0010001101110001;
            14'h0b6f 	:	o_val <= 16'b0010001101110100;
            14'h0b70 	:	o_val <= 16'b0010001101110111;
            14'h0b71 	:	o_val <= 16'b0010001101111010;
            14'h0b72 	:	o_val <= 16'b0010001101111101;
            14'h0b73 	:	o_val <= 16'b0010001110000000;
            14'h0b74 	:	o_val <= 16'b0010001110000011;
            14'h0b75 	:	o_val <= 16'b0010001110000110;
            14'h0b76 	:	o_val <= 16'b0010001110001001;
            14'h0b77 	:	o_val <= 16'b0010001110001100;
            14'h0b78 	:	o_val <= 16'b0010001110001111;
            14'h0b79 	:	o_val <= 16'b0010001110010010;
            14'h0b7a 	:	o_val <= 16'b0010001110010101;
            14'h0b7b 	:	o_val <= 16'b0010001110011000;
            14'h0b7c 	:	o_val <= 16'b0010001110011011;
            14'h0b7d 	:	o_val <= 16'b0010001110011110;
            14'h0b7e 	:	o_val <= 16'b0010001110100010;
            14'h0b7f 	:	o_val <= 16'b0010001110100101;
            14'h0b80 	:	o_val <= 16'b0010001110101000;
            14'h0b81 	:	o_val <= 16'b0010001110101011;
            14'h0b82 	:	o_val <= 16'b0010001110101110;
            14'h0b83 	:	o_val <= 16'b0010001110110001;
            14'h0b84 	:	o_val <= 16'b0010001110110100;
            14'h0b85 	:	o_val <= 16'b0010001110110111;
            14'h0b86 	:	o_val <= 16'b0010001110111010;
            14'h0b87 	:	o_val <= 16'b0010001110111101;
            14'h0b88 	:	o_val <= 16'b0010001111000000;
            14'h0b89 	:	o_val <= 16'b0010001111000011;
            14'h0b8a 	:	o_val <= 16'b0010001111000110;
            14'h0b8b 	:	o_val <= 16'b0010001111001001;
            14'h0b8c 	:	o_val <= 16'b0010001111001100;
            14'h0b8d 	:	o_val <= 16'b0010001111001111;
            14'h0b8e 	:	o_val <= 16'b0010001111010010;
            14'h0b8f 	:	o_val <= 16'b0010001111010101;
            14'h0b90 	:	o_val <= 16'b0010001111011000;
            14'h0b91 	:	o_val <= 16'b0010001111011011;
            14'h0b92 	:	o_val <= 16'b0010001111011110;
            14'h0b93 	:	o_val <= 16'b0010001111100001;
            14'h0b94 	:	o_val <= 16'b0010001111100100;
            14'h0b95 	:	o_val <= 16'b0010001111100111;
            14'h0b96 	:	o_val <= 16'b0010001111101010;
            14'h0b97 	:	o_val <= 16'b0010001111101101;
            14'h0b98 	:	o_val <= 16'b0010001111110000;
            14'h0b99 	:	o_val <= 16'b0010001111110011;
            14'h0b9a 	:	o_val <= 16'b0010001111110110;
            14'h0b9b 	:	o_val <= 16'b0010001111111001;
            14'h0b9c 	:	o_val <= 16'b0010001111111100;
            14'h0b9d 	:	o_val <= 16'b0010001111111111;
            14'h0b9e 	:	o_val <= 16'b0010010000000010;
            14'h0b9f 	:	o_val <= 16'b0010010000000101;
            14'h0ba0 	:	o_val <= 16'b0010010000001000;
            14'h0ba1 	:	o_val <= 16'b0010010000001011;
            14'h0ba2 	:	o_val <= 16'b0010010000001110;
            14'h0ba3 	:	o_val <= 16'b0010010000010001;
            14'h0ba4 	:	o_val <= 16'b0010010000010100;
            14'h0ba5 	:	o_val <= 16'b0010010000010111;
            14'h0ba6 	:	o_val <= 16'b0010010000011010;
            14'h0ba7 	:	o_val <= 16'b0010010000011101;
            14'h0ba8 	:	o_val <= 16'b0010010000100000;
            14'h0ba9 	:	o_val <= 16'b0010010000100011;
            14'h0baa 	:	o_val <= 16'b0010010000100110;
            14'h0bab 	:	o_val <= 16'b0010010000101001;
            14'h0bac 	:	o_val <= 16'b0010010000101100;
            14'h0bad 	:	o_val <= 16'b0010010000101111;
            14'h0bae 	:	o_val <= 16'b0010010000110010;
            14'h0baf 	:	o_val <= 16'b0010010000110101;
            14'h0bb0 	:	o_val <= 16'b0010010000111000;
            14'h0bb1 	:	o_val <= 16'b0010010000111011;
            14'h0bb2 	:	o_val <= 16'b0010010000111110;
            14'h0bb3 	:	o_val <= 16'b0010010001000001;
            14'h0bb4 	:	o_val <= 16'b0010010001000100;
            14'h0bb5 	:	o_val <= 16'b0010010001000111;
            14'h0bb6 	:	o_val <= 16'b0010010001001010;
            14'h0bb7 	:	o_val <= 16'b0010010001001101;
            14'h0bb8 	:	o_val <= 16'b0010010001010000;
            14'h0bb9 	:	o_val <= 16'b0010010001010011;
            14'h0bba 	:	o_val <= 16'b0010010001010110;
            14'h0bbb 	:	o_val <= 16'b0010010001011001;
            14'h0bbc 	:	o_val <= 16'b0010010001011100;
            14'h0bbd 	:	o_val <= 16'b0010010001011111;
            14'h0bbe 	:	o_val <= 16'b0010010001100010;
            14'h0bbf 	:	o_val <= 16'b0010010001100101;
            14'h0bc0 	:	o_val <= 16'b0010010001101000;
            14'h0bc1 	:	o_val <= 16'b0010010001101011;
            14'h0bc2 	:	o_val <= 16'b0010010001101110;
            14'h0bc3 	:	o_val <= 16'b0010010001110010;
            14'h0bc4 	:	o_val <= 16'b0010010001110101;
            14'h0bc5 	:	o_val <= 16'b0010010001111000;
            14'h0bc6 	:	o_val <= 16'b0010010001111011;
            14'h0bc7 	:	o_val <= 16'b0010010001111110;
            14'h0bc8 	:	o_val <= 16'b0010010010000001;
            14'h0bc9 	:	o_val <= 16'b0010010010000100;
            14'h0bca 	:	o_val <= 16'b0010010010000111;
            14'h0bcb 	:	o_val <= 16'b0010010010001010;
            14'h0bcc 	:	o_val <= 16'b0010010010001101;
            14'h0bcd 	:	o_val <= 16'b0010010010010000;
            14'h0bce 	:	o_val <= 16'b0010010010010011;
            14'h0bcf 	:	o_val <= 16'b0010010010010110;
            14'h0bd0 	:	o_val <= 16'b0010010010011001;
            14'h0bd1 	:	o_val <= 16'b0010010010011100;
            14'h0bd2 	:	o_val <= 16'b0010010010011111;
            14'h0bd3 	:	o_val <= 16'b0010010010100010;
            14'h0bd4 	:	o_val <= 16'b0010010010100101;
            14'h0bd5 	:	o_val <= 16'b0010010010101000;
            14'h0bd6 	:	o_val <= 16'b0010010010101011;
            14'h0bd7 	:	o_val <= 16'b0010010010101110;
            14'h0bd8 	:	o_val <= 16'b0010010010110001;
            14'h0bd9 	:	o_val <= 16'b0010010010110100;
            14'h0bda 	:	o_val <= 16'b0010010010110111;
            14'h0bdb 	:	o_val <= 16'b0010010010111010;
            14'h0bdc 	:	o_val <= 16'b0010010010111101;
            14'h0bdd 	:	o_val <= 16'b0010010011000000;
            14'h0bde 	:	o_val <= 16'b0010010011000011;
            14'h0bdf 	:	o_val <= 16'b0010010011000110;
            14'h0be0 	:	o_val <= 16'b0010010011001001;
            14'h0be1 	:	o_val <= 16'b0010010011001100;
            14'h0be2 	:	o_val <= 16'b0010010011001111;
            14'h0be3 	:	o_val <= 16'b0010010011010010;
            14'h0be4 	:	o_val <= 16'b0010010011010101;
            14'h0be5 	:	o_val <= 16'b0010010011011000;
            14'h0be6 	:	o_val <= 16'b0010010011011011;
            14'h0be7 	:	o_val <= 16'b0010010011011110;
            14'h0be8 	:	o_val <= 16'b0010010011100001;
            14'h0be9 	:	o_val <= 16'b0010010011100100;
            14'h0bea 	:	o_val <= 16'b0010010011100111;
            14'h0beb 	:	o_val <= 16'b0010010011101010;
            14'h0bec 	:	o_val <= 16'b0010010011101101;
            14'h0bed 	:	o_val <= 16'b0010010011110000;
            14'h0bee 	:	o_val <= 16'b0010010011110011;
            14'h0bef 	:	o_val <= 16'b0010010011110110;
            14'h0bf0 	:	o_val <= 16'b0010010011111001;
            14'h0bf1 	:	o_val <= 16'b0010010011111100;
            14'h0bf2 	:	o_val <= 16'b0010010011111111;
            14'h0bf3 	:	o_val <= 16'b0010010100000010;
            14'h0bf4 	:	o_val <= 16'b0010010100000101;
            14'h0bf5 	:	o_val <= 16'b0010010100001000;
            14'h0bf6 	:	o_val <= 16'b0010010100001011;
            14'h0bf7 	:	o_val <= 16'b0010010100001110;
            14'h0bf8 	:	o_val <= 16'b0010010100010001;
            14'h0bf9 	:	o_val <= 16'b0010010100010100;
            14'h0bfa 	:	o_val <= 16'b0010010100010111;
            14'h0bfb 	:	o_val <= 16'b0010010100011010;
            14'h0bfc 	:	o_val <= 16'b0010010100011101;
            14'h0bfd 	:	o_val <= 16'b0010010100100000;
            14'h0bfe 	:	o_val <= 16'b0010010100100011;
            14'h0bff 	:	o_val <= 16'b0010010100100110;
            14'h0c00 	:	o_val <= 16'b0010010100101001;
            14'h0c01 	:	o_val <= 16'b0010010100101100;
            14'h0c02 	:	o_val <= 16'b0010010100101111;
            14'h0c03 	:	o_val <= 16'b0010010100110010;
            14'h0c04 	:	o_val <= 16'b0010010100110101;
            14'h0c05 	:	o_val <= 16'b0010010100111000;
            14'h0c06 	:	o_val <= 16'b0010010100111011;
            14'h0c07 	:	o_val <= 16'b0010010100111110;
            14'h0c08 	:	o_val <= 16'b0010010101000001;
            14'h0c09 	:	o_val <= 16'b0010010101000100;
            14'h0c0a 	:	o_val <= 16'b0010010101000111;
            14'h0c0b 	:	o_val <= 16'b0010010101001010;
            14'h0c0c 	:	o_val <= 16'b0010010101001101;
            14'h0c0d 	:	o_val <= 16'b0010010101010000;
            14'h0c0e 	:	o_val <= 16'b0010010101010011;
            14'h0c0f 	:	o_val <= 16'b0010010101010110;
            14'h0c10 	:	o_val <= 16'b0010010101011001;
            14'h0c11 	:	o_val <= 16'b0010010101011100;
            14'h0c12 	:	o_val <= 16'b0010010101011111;
            14'h0c13 	:	o_val <= 16'b0010010101100010;
            14'h0c14 	:	o_val <= 16'b0010010101100101;
            14'h0c15 	:	o_val <= 16'b0010010101101000;
            14'h0c16 	:	o_val <= 16'b0010010101101011;
            14'h0c17 	:	o_val <= 16'b0010010101101110;
            14'h0c18 	:	o_val <= 16'b0010010101110001;
            14'h0c19 	:	o_val <= 16'b0010010101110100;
            14'h0c1a 	:	o_val <= 16'b0010010101110111;
            14'h0c1b 	:	o_val <= 16'b0010010101111010;
            14'h0c1c 	:	o_val <= 16'b0010010101111101;
            14'h0c1d 	:	o_val <= 16'b0010010110000000;
            14'h0c1e 	:	o_val <= 16'b0010010110000011;
            14'h0c1f 	:	o_val <= 16'b0010010110000110;
            14'h0c20 	:	o_val <= 16'b0010010110001001;
            14'h0c21 	:	o_val <= 16'b0010010110001100;
            14'h0c22 	:	o_val <= 16'b0010010110001111;
            14'h0c23 	:	o_val <= 16'b0010010110010010;
            14'h0c24 	:	o_val <= 16'b0010010110010101;
            14'h0c25 	:	o_val <= 16'b0010010110011000;
            14'h0c26 	:	o_val <= 16'b0010010110011011;
            14'h0c27 	:	o_val <= 16'b0010010110011110;
            14'h0c28 	:	o_val <= 16'b0010010110100001;
            14'h0c29 	:	o_val <= 16'b0010010110100100;
            14'h0c2a 	:	o_val <= 16'b0010010110100111;
            14'h0c2b 	:	o_val <= 16'b0010010110101010;
            14'h0c2c 	:	o_val <= 16'b0010010110101101;
            14'h0c2d 	:	o_val <= 16'b0010010110110000;
            14'h0c2e 	:	o_val <= 16'b0010010110110011;
            14'h0c2f 	:	o_val <= 16'b0010010110110110;
            14'h0c30 	:	o_val <= 16'b0010010110111001;
            14'h0c31 	:	o_val <= 16'b0010010110111100;
            14'h0c32 	:	o_val <= 16'b0010010110111111;
            14'h0c33 	:	o_val <= 16'b0010010111000010;
            14'h0c34 	:	o_val <= 16'b0010010111000101;
            14'h0c35 	:	o_val <= 16'b0010010111001000;
            14'h0c36 	:	o_val <= 16'b0010010111001011;
            14'h0c37 	:	o_val <= 16'b0010010111001110;
            14'h0c38 	:	o_val <= 16'b0010010111010001;
            14'h0c39 	:	o_val <= 16'b0010010111010100;
            14'h0c3a 	:	o_val <= 16'b0010010111010111;
            14'h0c3b 	:	o_val <= 16'b0010010111011010;
            14'h0c3c 	:	o_val <= 16'b0010010111011101;
            14'h0c3d 	:	o_val <= 16'b0010010111100000;
            14'h0c3e 	:	o_val <= 16'b0010010111100011;
            14'h0c3f 	:	o_val <= 16'b0010010111100110;
            14'h0c40 	:	o_val <= 16'b0010010111101001;
            14'h0c41 	:	o_val <= 16'b0010010111101100;
            14'h0c42 	:	o_val <= 16'b0010010111101111;
            14'h0c43 	:	o_val <= 16'b0010010111110010;
            14'h0c44 	:	o_val <= 16'b0010010111110101;
            14'h0c45 	:	o_val <= 16'b0010010111111000;
            14'h0c46 	:	o_val <= 16'b0010010111111011;
            14'h0c47 	:	o_val <= 16'b0010010111111110;
            14'h0c48 	:	o_val <= 16'b0010011000000001;
            14'h0c49 	:	o_val <= 16'b0010011000000100;
            14'h0c4a 	:	o_val <= 16'b0010011000000111;
            14'h0c4b 	:	o_val <= 16'b0010011000001010;
            14'h0c4c 	:	o_val <= 16'b0010011000001101;
            14'h0c4d 	:	o_val <= 16'b0010011000010000;
            14'h0c4e 	:	o_val <= 16'b0010011000010011;
            14'h0c4f 	:	o_val <= 16'b0010011000010110;
            14'h0c50 	:	o_val <= 16'b0010011000011001;
            14'h0c51 	:	o_val <= 16'b0010011000011100;
            14'h0c52 	:	o_val <= 16'b0010011000011111;
            14'h0c53 	:	o_val <= 16'b0010011000100010;
            14'h0c54 	:	o_val <= 16'b0010011000100101;
            14'h0c55 	:	o_val <= 16'b0010011000101000;
            14'h0c56 	:	o_val <= 16'b0010011000101011;
            14'h0c57 	:	o_val <= 16'b0010011000101110;
            14'h0c58 	:	o_val <= 16'b0010011000110001;
            14'h0c59 	:	o_val <= 16'b0010011000110100;
            14'h0c5a 	:	o_val <= 16'b0010011000110111;
            14'h0c5b 	:	o_val <= 16'b0010011000111010;
            14'h0c5c 	:	o_val <= 16'b0010011000111101;
            14'h0c5d 	:	o_val <= 16'b0010011001000000;
            14'h0c5e 	:	o_val <= 16'b0010011001000011;
            14'h0c5f 	:	o_val <= 16'b0010011001000110;
            14'h0c60 	:	o_val <= 16'b0010011001001001;
            14'h0c61 	:	o_val <= 16'b0010011001001100;
            14'h0c62 	:	o_val <= 16'b0010011001001111;
            14'h0c63 	:	o_val <= 16'b0010011001010010;
            14'h0c64 	:	o_val <= 16'b0010011001010101;
            14'h0c65 	:	o_val <= 16'b0010011001011000;
            14'h0c66 	:	o_val <= 16'b0010011001011011;
            14'h0c67 	:	o_val <= 16'b0010011001011110;
            14'h0c68 	:	o_val <= 16'b0010011001100001;
            14'h0c69 	:	o_val <= 16'b0010011001100100;
            14'h0c6a 	:	o_val <= 16'b0010011001100111;
            14'h0c6b 	:	o_val <= 16'b0010011001101010;
            14'h0c6c 	:	o_val <= 16'b0010011001101101;
            14'h0c6d 	:	o_val <= 16'b0010011001110000;
            14'h0c6e 	:	o_val <= 16'b0010011001110011;
            14'h0c6f 	:	o_val <= 16'b0010011001110110;
            14'h0c70 	:	o_val <= 16'b0010011001111001;
            14'h0c71 	:	o_val <= 16'b0010011001111100;
            14'h0c72 	:	o_val <= 16'b0010011001111111;
            14'h0c73 	:	o_val <= 16'b0010011010000010;
            14'h0c74 	:	o_val <= 16'b0010011010000101;
            14'h0c75 	:	o_val <= 16'b0010011010001000;
            14'h0c76 	:	o_val <= 16'b0010011010001011;
            14'h0c77 	:	o_val <= 16'b0010011010001110;
            14'h0c78 	:	o_val <= 16'b0010011010010001;
            14'h0c79 	:	o_val <= 16'b0010011010010100;
            14'h0c7a 	:	o_val <= 16'b0010011010010111;
            14'h0c7b 	:	o_val <= 16'b0010011010011010;
            14'h0c7c 	:	o_val <= 16'b0010011010011101;
            14'h0c7d 	:	o_val <= 16'b0010011010100000;
            14'h0c7e 	:	o_val <= 16'b0010011010100011;
            14'h0c7f 	:	o_val <= 16'b0010011010100110;
            14'h0c80 	:	o_val <= 16'b0010011010101001;
            14'h0c81 	:	o_val <= 16'b0010011010101100;
            14'h0c82 	:	o_val <= 16'b0010011010101111;
            14'h0c83 	:	o_val <= 16'b0010011010110010;
            14'h0c84 	:	o_val <= 16'b0010011010110101;
            14'h0c85 	:	o_val <= 16'b0010011010111000;
            14'h0c86 	:	o_val <= 16'b0010011010111011;
            14'h0c87 	:	o_val <= 16'b0010011010111110;
            14'h0c88 	:	o_val <= 16'b0010011011000001;
            14'h0c89 	:	o_val <= 16'b0010011011000100;
            14'h0c8a 	:	o_val <= 16'b0010011011000111;
            14'h0c8b 	:	o_val <= 16'b0010011011001010;
            14'h0c8c 	:	o_val <= 16'b0010011011001101;
            14'h0c8d 	:	o_val <= 16'b0010011011010000;
            14'h0c8e 	:	o_val <= 16'b0010011011010011;
            14'h0c8f 	:	o_val <= 16'b0010011011010110;
            14'h0c90 	:	o_val <= 16'b0010011011011001;
            14'h0c91 	:	o_val <= 16'b0010011011011100;
            14'h0c92 	:	o_val <= 16'b0010011011011111;
            14'h0c93 	:	o_val <= 16'b0010011011100010;
            14'h0c94 	:	o_val <= 16'b0010011011100101;
            14'h0c95 	:	o_val <= 16'b0010011011101000;
            14'h0c96 	:	o_val <= 16'b0010011011101011;
            14'h0c97 	:	o_val <= 16'b0010011011101110;
            14'h0c98 	:	o_val <= 16'b0010011011110001;
            14'h0c99 	:	o_val <= 16'b0010011011110100;
            14'h0c9a 	:	o_val <= 16'b0010011011110111;
            14'h0c9b 	:	o_val <= 16'b0010011011111010;
            14'h0c9c 	:	o_val <= 16'b0010011011111101;
            14'h0c9d 	:	o_val <= 16'b0010011100000000;
            14'h0c9e 	:	o_val <= 16'b0010011100000011;
            14'h0c9f 	:	o_val <= 16'b0010011100000110;
            14'h0ca0 	:	o_val <= 16'b0010011100001001;
            14'h0ca1 	:	o_val <= 16'b0010011100001100;
            14'h0ca2 	:	o_val <= 16'b0010011100001111;
            14'h0ca3 	:	o_val <= 16'b0010011100010010;
            14'h0ca4 	:	o_val <= 16'b0010011100010101;
            14'h0ca5 	:	o_val <= 16'b0010011100011000;
            14'h0ca6 	:	o_val <= 16'b0010011100011011;
            14'h0ca7 	:	o_val <= 16'b0010011100011110;
            14'h0ca8 	:	o_val <= 16'b0010011100100001;
            14'h0ca9 	:	o_val <= 16'b0010011100100100;
            14'h0caa 	:	o_val <= 16'b0010011100100111;
            14'h0cab 	:	o_val <= 16'b0010011100101010;
            14'h0cac 	:	o_val <= 16'b0010011100101101;
            14'h0cad 	:	o_val <= 16'b0010011100110000;
            14'h0cae 	:	o_val <= 16'b0010011100110011;
            14'h0caf 	:	o_val <= 16'b0010011100110110;
            14'h0cb0 	:	o_val <= 16'b0010011100111001;
            14'h0cb1 	:	o_val <= 16'b0010011100111100;
            14'h0cb2 	:	o_val <= 16'b0010011100111111;
            14'h0cb3 	:	o_val <= 16'b0010011101000010;
            14'h0cb4 	:	o_val <= 16'b0010011101000101;
            14'h0cb5 	:	o_val <= 16'b0010011101001000;
            14'h0cb6 	:	o_val <= 16'b0010011101001011;
            14'h0cb7 	:	o_val <= 16'b0010011101001110;
            14'h0cb8 	:	o_val <= 16'b0010011101010001;
            14'h0cb9 	:	o_val <= 16'b0010011101010100;
            14'h0cba 	:	o_val <= 16'b0010011101010111;
            14'h0cbb 	:	o_val <= 16'b0010011101011010;
            14'h0cbc 	:	o_val <= 16'b0010011101011101;
            14'h0cbd 	:	o_val <= 16'b0010011101100000;
            14'h0cbe 	:	o_val <= 16'b0010011101100011;
            14'h0cbf 	:	o_val <= 16'b0010011101100110;
            14'h0cc0 	:	o_val <= 16'b0010011101101001;
            14'h0cc1 	:	o_val <= 16'b0010011101101100;
            14'h0cc2 	:	o_val <= 16'b0010011101101111;
            14'h0cc3 	:	o_val <= 16'b0010011101110010;
            14'h0cc4 	:	o_val <= 16'b0010011101110101;
            14'h0cc5 	:	o_val <= 16'b0010011101111000;
            14'h0cc6 	:	o_val <= 16'b0010011101111011;
            14'h0cc7 	:	o_val <= 16'b0010011101111110;
            14'h0cc8 	:	o_val <= 16'b0010011110000001;
            14'h0cc9 	:	o_val <= 16'b0010011110000100;
            14'h0cca 	:	o_val <= 16'b0010011110000110;
            14'h0ccb 	:	o_val <= 16'b0010011110001001;
            14'h0ccc 	:	o_val <= 16'b0010011110001100;
            14'h0ccd 	:	o_val <= 16'b0010011110001111;
            14'h0cce 	:	o_val <= 16'b0010011110010010;
            14'h0ccf 	:	o_val <= 16'b0010011110010101;
            14'h0cd0 	:	o_val <= 16'b0010011110011000;
            14'h0cd1 	:	o_val <= 16'b0010011110011011;
            14'h0cd2 	:	o_val <= 16'b0010011110011110;
            14'h0cd3 	:	o_val <= 16'b0010011110100001;
            14'h0cd4 	:	o_val <= 16'b0010011110100100;
            14'h0cd5 	:	o_val <= 16'b0010011110100111;
            14'h0cd6 	:	o_val <= 16'b0010011110101010;
            14'h0cd7 	:	o_val <= 16'b0010011110101101;
            14'h0cd8 	:	o_val <= 16'b0010011110110000;
            14'h0cd9 	:	o_val <= 16'b0010011110110011;
            14'h0cda 	:	o_val <= 16'b0010011110110110;
            14'h0cdb 	:	o_val <= 16'b0010011110111001;
            14'h0cdc 	:	o_val <= 16'b0010011110111100;
            14'h0cdd 	:	o_val <= 16'b0010011110111111;
            14'h0cde 	:	o_val <= 16'b0010011111000010;
            14'h0cdf 	:	o_val <= 16'b0010011111000101;
            14'h0ce0 	:	o_val <= 16'b0010011111001000;
            14'h0ce1 	:	o_val <= 16'b0010011111001011;
            14'h0ce2 	:	o_val <= 16'b0010011111001110;
            14'h0ce3 	:	o_val <= 16'b0010011111010001;
            14'h0ce4 	:	o_val <= 16'b0010011111010100;
            14'h0ce5 	:	o_val <= 16'b0010011111010111;
            14'h0ce6 	:	o_val <= 16'b0010011111011010;
            14'h0ce7 	:	o_val <= 16'b0010011111011101;
            14'h0ce8 	:	o_val <= 16'b0010011111100000;
            14'h0ce9 	:	o_val <= 16'b0010011111100011;
            14'h0cea 	:	o_val <= 16'b0010011111100110;
            14'h0ceb 	:	o_val <= 16'b0010011111101001;
            14'h0cec 	:	o_val <= 16'b0010011111101100;
            14'h0ced 	:	o_val <= 16'b0010011111101111;
            14'h0cee 	:	o_val <= 16'b0010011111110010;
            14'h0cef 	:	o_val <= 16'b0010011111110101;
            14'h0cf0 	:	o_val <= 16'b0010011111111000;
            14'h0cf1 	:	o_val <= 16'b0010011111111011;
            14'h0cf2 	:	o_val <= 16'b0010011111111110;
            14'h0cf3 	:	o_val <= 16'b0010100000000001;
            14'h0cf4 	:	o_val <= 16'b0010100000000100;
            14'h0cf5 	:	o_val <= 16'b0010100000000111;
            14'h0cf6 	:	o_val <= 16'b0010100000001010;
            14'h0cf7 	:	o_val <= 16'b0010100000001101;
            14'h0cf8 	:	o_val <= 16'b0010100000010000;
            14'h0cf9 	:	o_val <= 16'b0010100000010011;
            14'h0cfa 	:	o_val <= 16'b0010100000010110;
            14'h0cfb 	:	o_val <= 16'b0010100000011001;
            14'h0cfc 	:	o_val <= 16'b0010100000011100;
            14'h0cfd 	:	o_val <= 16'b0010100000011111;
            14'h0cfe 	:	o_val <= 16'b0010100000100010;
            14'h0cff 	:	o_val <= 16'b0010100000100101;
            14'h0d00 	:	o_val <= 16'b0010100000101000;
            14'h0d01 	:	o_val <= 16'b0010100000101011;
            14'h0d02 	:	o_val <= 16'b0010100000101110;
            14'h0d03 	:	o_val <= 16'b0010100000110001;
            14'h0d04 	:	o_val <= 16'b0010100000110100;
            14'h0d05 	:	o_val <= 16'b0010100000110111;
            14'h0d06 	:	o_val <= 16'b0010100000111010;
            14'h0d07 	:	o_val <= 16'b0010100000111101;
            14'h0d08 	:	o_val <= 16'b0010100001000000;
            14'h0d09 	:	o_val <= 16'b0010100001000011;
            14'h0d0a 	:	o_val <= 16'b0010100001000110;
            14'h0d0b 	:	o_val <= 16'b0010100001001001;
            14'h0d0c 	:	o_val <= 16'b0010100001001100;
            14'h0d0d 	:	o_val <= 16'b0010100001001110;
            14'h0d0e 	:	o_val <= 16'b0010100001010001;
            14'h0d0f 	:	o_val <= 16'b0010100001010100;
            14'h0d10 	:	o_val <= 16'b0010100001010111;
            14'h0d11 	:	o_val <= 16'b0010100001011010;
            14'h0d12 	:	o_val <= 16'b0010100001011101;
            14'h0d13 	:	o_val <= 16'b0010100001100000;
            14'h0d14 	:	o_val <= 16'b0010100001100011;
            14'h0d15 	:	o_val <= 16'b0010100001100110;
            14'h0d16 	:	o_val <= 16'b0010100001101001;
            14'h0d17 	:	o_val <= 16'b0010100001101100;
            14'h0d18 	:	o_val <= 16'b0010100001101111;
            14'h0d19 	:	o_val <= 16'b0010100001110010;
            14'h0d1a 	:	o_val <= 16'b0010100001110101;
            14'h0d1b 	:	o_val <= 16'b0010100001111000;
            14'h0d1c 	:	o_val <= 16'b0010100001111011;
            14'h0d1d 	:	o_val <= 16'b0010100001111110;
            14'h0d1e 	:	o_val <= 16'b0010100010000001;
            14'h0d1f 	:	o_val <= 16'b0010100010000100;
            14'h0d20 	:	o_val <= 16'b0010100010000111;
            14'h0d21 	:	o_val <= 16'b0010100010001010;
            14'h0d22 	:	o_val <= 16'b0010100010001101;
            14'h0d23 	:	o_val <= 16'b0010100010010000;
            14'h0d24 	:	o_val <= 16'b0010100010010011;
            14'h0d25 	:	o_val <= 16'b0010100010010110;
            14'h0d26 	:	o_val <= 16'b0010100010011001;
            14'h0d27 	:	o_val <= 16'b0010100010011100;
            14'h0d28 	:	o_val <= 16'b0010100010011111;
            14'h0d29 	:	o_val <= 16'b0010100010100010;
            14'h0d2a 	:	o_val <= 16'b0010100010100101;
            14'h0d2b 	:	o_val <= 16'b0010100010101000;
            14'h0d2c 	:	o_val <= 16'b0010100010101011;
            14'h0d2d 	:	o_val <= 16'b0010100010101110;
            14'h0d2e 	:	o_val <= 16'b0010100010110001;
            14'h0d2f 	:	o_val <= 16'b0010100010110100;
            14'h0d30 	:	o_val <= 16'b0010100010110111;
            14'h0d31 	:	o_val <= 16'b0010100010111010;
            14'h0d32 	:	o_val <= 16'b0010100010111101;
            14'h0d33 	:	o_val <= 16'b0010100011000000;
            14'h0d34 	:	o_val <= 16'b0010100011000011;
            14'h0d35 	:	o_val <= 16'b0010100011000110;
            14'h0d36 	:	o_val <= 16'b0010100011001001;
            14'h0d37 	:	o_val <= 16'b0010100011001100;
            14'h0d38 	:	o_val <= 16'b0010100011001111;
            14'h0d39 	:	o_val <= 16'b0010100011010010;
            14'h0d3a 	:	o_val <= 16'b0010100011010101;
            14'h0d3b 	:	o_val <= 16'b0010100011011000;
            14'h0d3c 	:	o_val <= 16'b0010100011011011;
            14'h0d3d 	:	o_val <= 16'b0010100011011101;
            14'h0d3e 	:	o_val <= 16'b0010100011100000;
            14'h0d3f 	:	o_val <= 16'b0010100011100011;
            14'h0d40 	:	o_val <= 16'b0010100011100110;
            14'h0d41 	:	o_val <= 16'b0010100011101001;
            14'h0d42 	:	o_val <= 16'b0010100011101100;
            14'h0d43 	:	o_val <= 16'b0010100011101111;
            14'h0d44 	:	o_val <= 16'b0010100011110010;
            14'h0d45 	:	o_val <= 16'b0010100011110101;
            14'h0d46 	:	o_val <= 16'b0010100011111000;
            14'h0d47 	:	o_val <= 16'b0010100011111011;
            14'h0d48 	:	o_val <= 16'b0010100011111110;
            14'h0d49 	:	o_val <= 16'b0010100100000001;
            14'h0d4a 	:	o_val <= 16'b0010100100000100;
            14'h0d4b 	:	o_val <= 16'b0010100100000111;
            14'h0d4c 	:	o_val <= 16'b0010100100001010;
            14'h0d4d 	:	o_val <= 16'b0010100100001101;
            14'h0d4e 	:	o_val <= 16'b0010100100010000;
            14'h0d4f 	:	o_val <= 16'b0010100100010011;
            14'h0d50 	:	o_val <= 16'b0010100100010110;
            14'h0d51 	:	o_val <= 16'b0010100100011001;
            14'h0d52 	:	o_val <= 16'b0010100100011100;
            14'h0d53 	:	o_val <= 16'b0010100100011111;
            14'h0d54 	:	o_val <= 16'b0010100100100010;
            14'h0d55 	:	o_val <= 16'b0010100100100101;
            14'h0d56 	:	o_val <= 16'b0010100100101000;
            14'h0d57 	:	o_val <= 16'b0010100100101011;
            14'h0d58 	:	o_val <= 16'b0010100100101110;
            14'h0d59 	:	o_val <= 16'b0010100100110001;
            14'h0d5a 	:	o_val <= 16'b0010100100110100;
            14'h0d5b 	:	o_val <= 16'b0010100100110111;
            14'h0d5c 	:	o_val <= 16'b0010100100111010;
            14'h0d5d 	:	o_val <= 16'b0010100100111101;
            14'h0d5e 	:	o_val <= 16'b0010100101000000;
            14'h0d5f 	:	o_val <= 16'b0010100101000011;
            14'h0d60 	:	o_val <= 16'b0010100101000110;
            14'h0d61 	:	o_val <= 16'b0010100101001001;
            14'h0d62 	:	o_val <= 16'b0010100101001100;
            14'h0d63 	:	o_val <= 16'b0010100101001111;
            14'h0d64 	:	o_val <= 16'b0010100101010010;
            14'h0d65 	:	o_val <= 16'b0010100101010101;
            14'h0d66 	:	o_val <= 16'b0010100101010111;
            14'h0d67 	:	o_val <= 16'b0010100101011010;
            14'h0d68 	:	o_val <= 16'b0010100101011101;
            14'h0d69 	:	o_val <= 16'b0010100101100000;
            14'h0d6a 	:	o_val <= 16'b0010100101100011;
            14'h0d6b 	:	o_val <= 16'b0010100101100110;
            14'h0d6c 	:	o_val <= 16'b0010100101101001;
            14'h0d6d 	:	o_val <= 16'b0010100101101100;
            14'h0d6e 	:	o_val <= 16'b0010100101101111;
            14'h0d6f 	:	o_val <= 16'b0010100101110010;
            14'h0d70 	:	o_val <= 16'b0010100101110101;
            14'h0d71 	:	o_val <= 16'b0010100101111000;
            14'h0d72 	:	o_val <= 16'b0010100101111011;
            14'h0d73 	:	o_val <= 16'b0010100101111110;
            14'h0d74 	:	o_val <= 16'b0010100110000001;
            14'h0d75 	:	o_val <= 16'b0010100110000100;
            14'h0d76 	:	o_val <= 16'b0010100110000111;
            14'h0d77 	:	o_val <= 16'b0010100110001010;
            14'h0d78 	:	o_val <= 16'b0010100110001101;
            14'h0d79 	:	o_val <= 16'b0010100110010000;
            14'h0d7a 	:	o_val <= 16'b0010100110010011;
            14'h0d7b 	:	o_val <= 16'b0010100110010110;
            14'h0d7c 	:	o_val <= 16'b0010100110011001;
            14'h0d7d 	:	o_val <= 16'b0010100110011100;
            14'h0d7e 	:	o_val <= 16'b0010100110011111;
            14'h0d7f 	:	o_val <= 16'b0010100110100010;
            14'h0d80 	:	o_val <= 16'b0010100110100101;
            14'h0d81 	:	o_val <= 16'b0010100110101000;
            14'h0d82 	:	o_val <= 16'b0010100110101011;
            14'h0d83 	:	o_val <= 16'b0010100110101110;
            14'h0d84 	:	o_val <= 16'b0010100110110001;
            14'h0d85 	:	o_val <= 16'b0010100110110100;
            14'h0d86 	:	o_val <= 16'b0010100110110111;
            14'h0d87 	:	o_val <= 16'b0010100110111010;
            14'h0d88 	:	o_val <= 16'b0010100110111101;
            14'h0d89 	:	o_val <= 16'b0010100110111111;
            14'h0d8a 	:	o_val <= 16'b0010100111000010;
            14'h0d8b 	:	o_val <= 16'b0010100111000101;
            14'h0d8c 	:	o_val <= 16'b0010100111001000;
            14'h0d8d 	:	o_val <= 16'b0010100111001011;
            14'h0d8e 	:	o_val <= 16'b0010100111001110;
            14'h0d8f 	:	o_val <= 16'b0010100111010001;
            14'h0d90 	:	o_val <= 16'b0010100111010100;
            14'h0d91 	:	o_val <= 16'b0010100111010111;
            14'h0d92 	:	o_val <= 16'b0010100111011010;
            14'h0d93 	:	o_val <= 16'b0010100111011101;
            14'h0d94 	:	o_val <= 16'b0010100111100000;
            14'h0d95 	:	o_val <= 16'b0010100111100011;
            14'h0d96 	:	o_val <= 16'b0010100111100110;
            14'h0d97 	:	o_val <= 16'b0010100111101001;
            14'h0d98 	:	o_val <= 16'b0010100111101100;
            14'h0d99 	:	o_val <= 16'b0010100111101111;
            14'h0d9a 	:	o_val <= 16'b0010100111110010;
            14'h0d9b 	:	o_val <= 16'b0010100111110101;
            14'h0d9c 	:	o_val <= 16'b0010100111111000;
            14'h0d9d 	:	o_val <= 16'b0010100111111011;
            14'h0d9e 	:	o_val <= 16'b0010100111111110;
            14'h0d9f 	:	o_val <= 16'b0010101000000001;
            14'h0da0 	:	o_val <= 16'b0010101000000100;
            14'h0da1 	:	o_val <= 16'b0010101000000111;
            14'h0da2 	:	o_val <= 16'b0010101000001010;
            14'h0da3 	:	o_val <= 16'b0010101000001101;
            14'h0da4 	:	o_val <= 16'b0010101000010000;
            14'h0da5 	:	o_val <= 16'b0010101000010011;
            14'h0da6 	:	o_val <= 16'b0010101000010110;
            14'h0da7 	:	o_val <= 16'b0010101000011001;
            14'h0da8 	:	o_val <= 16'b0010101000011100;
            14'h0da9 	:	o_val <= 16'b0010101000011110;
            14'h0daa 	:	o_val <= 16'b0010101000100001;
            14'h0dab 	:	o_val <= 16'b0010101000100100;
            14'h0dac 	:	o_val <= 16'b0010101000100111;
            14'h0dad 	:	o_val <= 16'b0010101000101010;
            14'h0dae 	:	o_val <= 16'b0010101000101101;
            14'h0daf 	:	o_val <= 16'b0010101000110000;
            14'h0db0 	:	o_val <= 16'b0010101000110011;
            14'h0db1 	:	o_val <= 16'b0010101000110110;
            14'h0db2 	:	o_val <= 16'b0010101000111001;
            14'h0db3 	:	o_val <= 16'b0010101000111100;
            14'h0db4 	:	o_val <= 16'b0010101000111111;
            14'h0db5 	:	o_val <= 16'b0010101001000010;
            14'h0db6 	:	o_val <= 16'b0010101001000101;
            14'h0db7 	:	o_val <= 16'b0010101001001000;
            14'h0db8 	:	o_val <= 16'b0010101001001011;
            14'h0db9 	:	o_val <= 16'b0010101001001110;
            14'h0dba 	:	o_val <= 16'b0010101001010001;
            14'h0dbb 	:	o_val <= 16'b0010101001010100;
            14'h0dbc 	:	o_val <= 16'b0010101001010111;
            14'h0dbd 	:	o_val <= 16'b0010101001011010;
            14'h0dbe 	:	o_val <= 16'b0010101001011101;
            14'h0dbf 	:	o_val <= 16'b0010101001100000;
            14'h0dc0 	:	o_val <= 16'b0010101001100011;
            14'h0dc1 	:	o_val <= 16'b0010101001100110;
            14'h0dc2 	:	o_val <= 16'b0010101001101001;
            14'h0dc3 	:	o_val <= 16'b0010101001101100;
            14'h0dc4 	:	o_val <= 16'b0010101001101111;
            14'h0dc5 	:	o_val <= 16'b0010101001110001;
            14'h0dc6 	:	o_val <= 16'b0010101001110100;
            14'h0dc7 	:	o_val <= 16'b0010101001110111;
            14'h0dc8 	:	o_val <= 16'b0010101001111010;
            14'h0dc9 	:	o_val <= 16'b0010101001111101;
            14'h0dca 	:	o_val <= 16'b0010101010000000;
            14'h0dcb 	:	o_val <= 16'b0010101010000011;
            14'h0dcc 	:	o_val <= 16'b0010101010000110;
            14'h0dcd 	:	o_val <= 16'b0010101010001001;
            14'h0dce 	:	o_val <= 16'b0010101010001100;
            14'h0dcf 	:	o_val <= 16'b0010101010001111;
            14'h0dd0 	:	o_val <= 16'b0010101010010010;
            14'h0dd1 	:	o_val <= 16'b0010101010010101;
            14'h0dd2 	:	o_val <= 16'b0010101010011000;
            14'h0dd3 	:	o_val <= 16'b0010101010011011;
            14'h0dd4 	:	o_val <= 16'b0010101010011110;
            14'h0dd5 	:	o_val <= 16'b0010101010100001;
            14'h0dd6 	:	o_val <= 16'b0010101010100100;
            14'h0dd7 	:	o_val <= 16'b0010101010100111;
            14'h0dd8 	:	o_val <= 16'b0010101010101010;
            14'h0dd9 	:	o_val <= 16'b0010101010101101;
            14'h0dda 	:	o_val <= 16'b0010101010110000;
            14'h0ddb 	:	o_val <= 16'b0010101010110011;
            14'h0ddc 	:	o_val <= 16'b0010101010110110;
            14'h0ddd 	:	o_val <= 16'b0010101010111001;
            14'h0dde 	:	o_val <= 16'b0010101010111100;
            14'h0ddf 	:	o_val <= 16'b0010101010111111;
            14'h0de0 	:	o_val <= 16'b0010101011000001;
            14'h0de1 	:	o_val <= 16'b0010101011000100;
            14'h0de2 	:	o_val <= 16'b0010101011000111;
            14'h0de3 	:	o_val <= 16'b0010101011001010;
            14'h0de4 	:	o_val <= 16'b0010101011001101;
            14'h0de5 	:	o_val <= 16'b0010101011010000;
            14'h0de6 	:	o_val <= 16'b0010101011010011;
            14'h0de7 	:	o_val <= 16'b0010101011010110;
            14'h0de8 	:	o_val <= 16'b0010101011011001;
            14'h0de9 	:	o_val <= 16'b0010101011011100;
            14'h0dea 	:	o_val <= 16'b0010101011011111;
            14'h0deb 	:	o_val <= 16'b0010101011100010;
            14'h0dec 	:	o_val <= 16'b0010101011100101;
            14'h0ded 	:	o_val <= 16'b0010101011101000;
            14'h0dee 	:	o_val <= 16'b0010101011101011;
            14'h0def 	:	o_val <= 16'b0010101011101110;
            14'h0df0 	:	o_val <= 16'b0010101011110001;
            14'h0df1 	:	o_val <= 16'b0010101011110100;
            14'h0df2 	:	o_val <= 16'b0010101011110111;
            14'h0df3 	:	o_val <= 16'b0010101011111010;
            14'h0df4 	:	o_val <= 16'b0010101011111101;
            14'h0df5 	:	o_val <= 16'b0010101100000000;
            14'h0df6 	:	o_val <= 16'b0010101100000011;
            14'h0df7 	:	o_val <= 16'b0010101100000110;
            14'h0df8 	:	o_val <= 16'b0010101100001001;
            14'h0df9 	:	o_val <= 16'b0010101100001011;
            14'h0dfa 	:	o_val <= 16'b0010101100001110;
            14'h0dfb 	:	o_val <= 16'b0010101100010001;
            14'h0dfc 	:	o_val <= 16'b0010101100010100;
            14'h0dfd 	:	o_val <= 16'b0010101100010111;
            14'h0dfe 	:	o_val <= 16'b0010101100011010;
            14'h0dff 	:	o_val <= 16'b0010101100011101;
            14'h0e00 	:	o_val <= 16'b0010101100100000;
            14'h0e01 	:	o_val <= 16'b0010101100100011;
            14'h0e02 	:	o_val <= 16'b0010101100100110;
            14'h0e03 	:	o_val <= 16'b0010101100101001;
            14'h0e04 	:	o_val <= 16'b0010101100101100;
            14'h0e05 	:	o_val <= 16'b0010101100101111;
            14'h0e06 	:	o_val <= 16'b0010101100110010;
            14'h0e07 	:	o_val <= 16'b0010101100110101;
            14'h0e08 	:	o_val <= 16'b0010101100111000;
            14'h0e09 	:	o_val <= 16'b0010101100111011;
            14'h0e0a 	:	o_val <= 16'b0010101100111110;
            14'h0e0b 	:	o_val <= 16'b0010101101000001;
            14'h0e0c 	:	o_val <= 16'b0010101101000100;
            14'h0e0d 	:	o_val <= 16'b0010101101000111;
            14'h0e0e 	:	o_val <= 16'b0010101101001010;
            14'h0e0f 	:	o_val <= 16'b0010101101001101;
            14'h0e10 	:	o_val <= 16'b0010101101001111;
            14'h0e11 	:	o_val <= 16'b0010101101010010;
            14'h0e12 	:	o_val <= 16'b0010101101010101;
            14'h0e13 	:	o_val <= 16'b0010101101011000;
            14'h0e14 	:	o_val <= 16'b0010101101011011;
            14'h0e15 	:	o_val <= 16'b0010101101011110;
            14'h0e16 	:	o_val <= 16'b0010101101100001;
            14'h0e17 	:	o_val <= 16'b0010101101100100;
            14'h0e18 	:	o_val <= 16'b0010101101100111;
            14'h0e19 	:	o_val <= 16'b0010101101101010;
            14'h0e1a 	:	o_val <= 16'b0010101101101101;
            14'h0e1b 	:	o_val <= 16'b0010101101110000;
            14'h0e1c 	:	o_val <= 16'b0010101101110011;
            14'h0e1d 	:	o_val <= 16'b0010101101110110;
            14'h0e1e 	:	o_val <= 16'b0010101101111001;
            14'h0e1f 	:	o_val <= 16'b0010101101111100;
            14'h0e20 	:	o_val <= 16'b0010101101111111;
            14'h0e21 	:	o_val <= 16'b0010101110000010;
            14'h0e22 	:	o_val <= 16'b0010101110000101;
            14'h0e23 	:	o_val <= 16'b0010101110001000;
            14'h0e24 	:	o_val <= 16'b0010101110001011;
            14'h0e25 	:	o_val <= 16'b0010101110001110;
            14'h0e26 	:	o_val <= 16'b0010101110010001;
            14'h0e27 	:	o_val <= 16'b0010101110010011;
            14'h0e28 	:	o_val <= 16'b0010101110010110;
            14'h0e29 	:	o_val <= 16'b0010101110011001;
            14'h0e2a 	:	o_val <= 16'b0010101110011100;
            14'h0e2b 	:	o_val <= 16'b0010101110011111;
            14'h0e2c 	:	o_val <= 16'b0010101110100010;
            14'h0e2d 	:	o_val <= 16'b0010101110100101;
            14'h0e2e 	:	o_val <= 16'b0010101110101000;
            14'h0e2f 	:	o_val <= 16'b0010101110101011;
            14'h0e30 	:	o_val <= 16'b0010101110101110;
            14'h0e31 	:	o_val <= 16'b0010101110110001;
            14'h0e32 	:	o_val <= 16'b0010101110110100;
            14'h0e33 	:	o_val <= 16'b0010101110110111;
            14'h0e34 	:	o_val <= 16'b0010101110111010;
            14'h0e35 	:	o_val <= 16'b0010101110111101;
            14'h0e36 	:	o_val <= 16'b0010101111000000;
            14'h0e37 	:	o_val <= 16'b0010101111000011;
            14'h0e38 	:	o_val <= 16'b0010101111000110;
            14'h0e39 	:	o_val <= 16'b0010101111001001;
            14'h0e3a 	:	o_val <= 16'b0010101111001100;
            14'h0e3b 	:	o_val <= 16'b0010101111001111;
            14'h0e3c 	:	o_val <= 16'b0010101111010001;
            14'h0e3d 	:	o_val <= 16'b0010101111010100;
            14'h0e3e 	:	o_val <= 16'b0010101111010111;
            14'h0e3f 	:	o_val <= 16'b0010101111011010;
            14'h0e40 	:	o_val <= 16'b0010101111011101;
            14'h0e41 	:	o_val <= 16'b0010101111100000;
            14'h0e42 	:	o_val <= 16'b0010101111100011;
            14'h0e43 	:	o_val <= 16'b0010101111100110;
            14'h0e44 	:	o_val <= 16'b0010101111101001;
            14'h0e45 	:	o_val <= 16'b0010101111101100;
            14'h0e46 	:	o_val <= 16'b0010101111101111;
            14'h0e47 	:	o_val <= 16'b0010101111110010;
            14'h0e48 	:	o_val <= 16'b0010101111110101;
            14'h0e49 	:	o_val <= 16'b0010101111111000;
            14'h0e4a 	:	o_val <= 16'b0010101111111011;
            14'h0e4b 	:	o_val <= 16'b0010101111111110;
            14'h0e4c 	:	o_val <= 16'b0010110000000001;
            14'h0e4d 	:	o_val <= 16'b0010110000000100;
            14'h0e4e 	:	o_val <= 16'b0010110000000111;
            14'h0e4f 	:	o_val <= 16'b0010110000001010;
            14'h0e50 	:	o_val <= 16'b0010110000001100;
            14'h0e51 	:	o_val <= 16'b0010110000001111;
            14'h0e52 	:	o_val <= 16'b0010110000010010;
            14'h0e53 	:	o_val <= 16'b0010110000010101;
            14'h0e54 	:	o_val <= 16'b0010110000011000;
            14'h0e55 	:	o_val <= 16'b0010110000011011;
            14'h0e56 	:	o_val <= 16'b0010110000011110;
            14'h0e57 	:	o_val <= 16'b0010110000100001;
            14'h0e58 	:	o_val <= 16'b0010110000100100;
            14'h0e59 	:	o_val <= 16'b0010110000100111;
            14'h0e5a 	:	o_val <= 16'b0010110000101010;
            14'h0e5b 	:	o_val <= 16'b0010110000101101;
            14'h0e5c 	:	o_val <= 16'b0010110000110000;
            14'h0e5d 	:	o_val <= 16'b0010110000110011;
            14'h0e5e 	:	o_val <= 16'b0010110000110110;
            14'h0e5f 	:	o_val <= 16'b0010110000111001;
            14'h0e60 	:	o_val <= 16'b0010110000111100;
            14'h0e61 	:	o_val <= 16'b0010110000111111;
            14'h0e62 	:	o_val <= 16'b0010110001000010;
            14'h0e63 	:	o_val <= 16'b0010110001000101;
            14'h0e64 	:	o_val <= 16'b0010110001000111;
            14'h0e65 	:	o_val <= 16'b0010110001001010;
            14'h0e66 	:	o_val <= 16'b0010110001001101;
            14'h0e67 	:	o_val <= 16'b0010110001010000;
            14'h0e68 	:	o_val <= 16'b0010110001010011;
            14'h0e69 	:	o_val <= 16'b0010110001010110;
            14'h0e6a 	:	o_val <= 16'b0010110001011001;
            14'h0e6b 	:	o_val <= 16'b0010110001011100;
            14'h0e6c 	:	o_val <= 16'b0010110001011111;
            14'h0e6d 	:	o_val <= 16'b0010110001100010;
            14'h0e6e 	:	o_val <= 16'b0010110001100101;
            14'h0e6f 	:	o_val <= 16'b0010110001101000;
            14'h0e70 	:	o_val <= 16'b0010110001101011;
            14'h0e71 	:	o_val <= 16'b0010110001101110;
            14'h0e72 	:	o_val <= 16'b0010110001110001;
            14'h0e73 	:	o_val <= 16'b0010110001110100;
            14'h0e74 	:	o_val <= 16'b0010110001110111;
            14'h0e75 	:	o_val <= 16'b0010110001111010;
            14'h0e76 	:	o_val <= 16'b0010110001111101;
            14'h0e77 	:	o_val <= 16'b0010110001111111;
            14'h0e78 	:	o_val <= 16'b0010110010000010;
            14'h0e79 	:	o_val <= 16'b0010110010000101;
            14'h0e7a 	:	o_val <= 16'b0010110010001000;
            14'h0e7b 	:	o_val <= 16'b0010110010001011;
            14'h0e7c 	:	o_val <= 16'b0010110010001110;
            14'h0e7d 	:	o_val <= 16'b0010110010010001;
            14'h0e7e 	:	o_val <= 16'b0010110010010100;
            14'h0e7f 	:	o_val <= 16'b0010110010010111;
            14'h0e80 	:	o_val <= 16'b0010110010011010;
            14'h0e81 	:	o_val <= 16'b0010110010011101;
            14'h0e82 	:	o_val <= 16'b0010110010100000;
            14'h0e83 	:	o_val <= 16'b0010110010100011;
            14'h0e84 	:	o_val <= 16'b0010110010100110;
            14'h0e85 	:	o_val <= 16'b0010110010101001;
            14'h0e86 	:	o_val <= 16'b0010110010101100;
            14'h0e87 	:	o_val <= 16'b0010110010101111;
            14'h0e88 	:	o_val <= 16'b0010110010110010;
            14'h0e89 	:	o_val <= 16'b0010110010110100;
            14'h0e8a 	:	o_val <= 16'b0010110010110111;
            14'h0e8b 	:	o_val <= 16'b0010110010111010;
            14'h0e8c 	:	o_val <= 16'b0010110010111101;
            14'h0e8d 	:	o_val <= 16'b0010110011000000;
            14'h0e8e 	:	o_val <= 16'b0010110011000011;
            14'h0e8f 	:	o_val <= 16'b0010110011000110;
            14'h0e90 	:	o_val <= 16'b0010110011001001;
            14'h0e91 	:	o_val <= 16'b0010110011001100;
            14'h0e92 	:	o_val <= 16'b0010110011001111;
            14'h0e93 	:	o_val <= 16'b0010110011010010;
            14'h0e94 	:	o_val <= 16'b0010110011010101;
            14'h0e95 	:	o_val <= 16'b0010110011011000;
            14'h0e96 	:	o_val <= 16'b0010110011011011;
            14'h0e97 	:	o_val <= 16'b0010110011011110;
            14'h0e98 	:	o_val <= 16'b0010110011100001;
            14'h0e99 	:	o_val <= 16'b0010110011100100;
            14'h0e9a 	:	o_val <= 16'b0010110011100110;
            14'h0e9b 	:	o_val <= 16'b0010110011101001;
            14'h0e9c 	:	o_val <= 16'b0010110011101100;
            14'h0e9d 	:	o_val <= 16'b0010110011101111;
            14'h0e9e 	:	o_val <= 16'b0010110011110010;
            14'h0e9f 	:	o_val <= 16'b0010110011110101;
            14'h0ea0 	:	o_val <= 16'b0010110011111000;
            14'h0ea1 	:	o_val <= 16'b0010110011111011;
            14'h0ea2 	:	o_val <= 16'b0010110011111110;
            14'h0ea3 	:	o_val <= 16'b0010110100000001;
            14'h0ea4 	:	o_val <= 16'b0010110100000100;
            14'h0ea5 	:	o_val <= 16'b0010110100000111;
            14'h0ea6 	:	o_val <= 16'b0010110100001010;
            14'h0ea7 	:	o_val <= 16'b0010110100001101;
            14'h0ea8 	:	o_val <= 16'b0010110100010000;
            14'h0ea9 	:	o_val <= 16'b0010110100010011;
            14'h0eaa 	:	o_val <= 16'b0010110100010110;
            14'h0eab 	:	o_val <= 16'b0010110100011000;
            14'h0eac 	:	o_val <= 16'b0010110100011011;
            14'h0ead 	:	o_val <= 16'b0010110100011110;
            14'h0eae 	:	o_val <= 16'b0010110100100001;
            14'h0eaf 	:	o_val <= 16'b0010110100100100;
            14'h0eb0 	:	o_val <= 16'b0010110100100111;
            14'h0eb1 	:	o_val <= 16'b0010110100101010;
            14'h0eb2 	:	o_val <= 16'b0010110100101101;
            14'h0eb3 	:	o_val <= 16'b0010110100110000;
            14'h0eb4 	:	o_val <= 16'b0010110100110011;
            14'h0eb5 	:	o_val <= 16'b0010110100110110;
            14'h0eb6 	:	o_val <= 16'b0010110100111001;
            14'h0eb7 	:	o_val <= 16'b0010110100111100;
            14'h0eb8 	:	o_val <= 16'b0010110100111111;
            14'h0eb9 	:	o_val <= 16'b0010110101000010;
            14'h0eba 	:	o_val <= 16'b0010110101000101;
            14'h0ebb 	:	o_val <= 16'b0010110101001000;
            14'h0ebc 	:	o_val <= 16'b0010110101001010;
            14'h0ebd 	:	o_val <= 16'b0010110101001101;
            14'h0ebe 	:	o_val <= 16'b0010110101010000;
            14'h0ebf 	:	o_val <= 16'b0010110101010011;
            14'h0ec0 	:	o_val <= 16'b0010110101010110;
            14'h0ec1 	:	o_val <= 16'b0010110101011001;
            14'h0ec2 	:	o_val <= 16'b0010110101011100;
            14'h0ec3 	:	o_val <= 16'b0010110101011111;
            14'h0ec4 	:	o_val <= 16'b0010110101100010;
            14'h0ec5 	:	o_val <= 16'b0010110101100101;
            14'h0ec6 	:	o_val <= 16'b0010110101101000;
            14'h0ec7 	:	o_val <= 16'b0010110101101011;
            14'h0ec8 	:	o_val <= 16'b0010110101101110;
            14'h0ec9 	:	o_val <= 16'b0010110101110001;
            14'h0eca 	:	o_val <= 16'b0010110101110100;
            14'h0ecb 	:	o_val <= 16'b0010110101110111;
            14'h0ecc 	:	o_val <= 16'b0010110101111001;
            14'h0ecd 	:	o_val <= 16'b0010110101111100;
            14'h0ece 	:	o_val <= 16'b0010110101111111;
            14'h0ecf 	:	o_val <= 16'b0010110110000010;
            14'h0ed0 	:	o_val <= 16'b0010110110000101;
            14'h0ed1 	:	o_val <= 16'b0010110110001000;
            14'h0ed2 	:	o_val <= 16'b0010110110001011;
            14'h0ed3 	:	o_val <= 16'b0010110110001110;
            14'h0ed4 	:	o_val <= 16'b0010110110010001;
            14'h0ed5 	:	o_val <= 16'b0010110110010100;
            14'h0ed6 	:	o_val <= 16'b0010110110010111;
            14'h0ed7 	:	o_val <= 16'b0010110110011010;
            14'h0ed8 	:	o_val <= 16'b0010110110011101;
            14'h0ed9 	:	o_val <= 16'b0010110110100000;
            14'h0eda 	:	o_val <= 16'b0010110110100011;
            14'h0edb 	:	o_val <= 16'b0010110110100101;
            14'h0edc 	:	o_val <= 16'b0010110110101000;
            14'h0edd 	:	o_val <= 16'b0010110110101011;
            14'h0ede 	:	o_val <= 16'b0010110110101110;
            14'h0edf 	:	o_val <= 16'b0010110110110001;
            14'h0ee0 	:	o_val <= 16'b0010110110110100;
            14'h0ee1 	:	o_val <= 16'b0010110110110111;
            14'h0ee2 	:	o_val <= 16'b0010110110111010;
            14'h0ee3 	:	o_val <= 16'b0010110110111101;
            14'h0ee4 	:	o_val <= 16'b0010110111000000;
            14'h0ee5 	:	o_val <= 16'b0010110111000011;
            14'h0ee6 	:	o_val <= 16'b0010110111000110;
            14'h0ee7 	:	o_val <= 16'b0010110111001001;
            14'h0ee8 	:	o_val <= 16'b0010110111001100;
            14'h0ee9 	:	o_val <= 16'b0010110111001111;
            14'h0eea 	:	o_val <= 16'b0010110111010001;
            14'h0eeb 	:	o_val <= 16'b0010110111010100;
            14'h0eec 	:	o_val <= 16'b0010110111010111;
            14'h0eed 	:	o_val <= 16'b0010110111011010;
            14'h0eee 	:	o_val <= 16'b0010110111011101;
            14'h0eef 	:	o_val <= 16'b0010110111100000;
            14'h0ef0 	:	o_val <= 16'b0010110111100011;
            14'h0ef1 	:	o_val <= 16'b0010110111100110;
            14'h0ef2 	:	o_val <= 16'b0010110111101001;
            14'h0ef3 	:	o_val <= 16'b0010110111101100;
            14'h0ef4 	:	o_val <= 16'b0010110111101111;
            14'h0ef5 	:	o_val <= 16'b0010110111110010;
            14'h0ef6 	:	o_val <= 16'b0010110111110101;
            14'h0ef7 	:	o_val <= 16'b0010110111111000;
            14'h0ef8 	:	o_val <= 16'b0010110111111011;
            14'h0ef9 	:	o_val <= 16'b0010110111111101;
            14'h0efa 	:	o_val <= 16'b0010111000000000;
            14'h0efb 	:	o_val <= 16'b0010111000000011;
            14'h0efc 	:	o_val <= 16'b0010111000000110;
            14'h0efd 	:	o_val <= 16'b0010111000001001;
            14'h0efe 	:	o_val <= 16'b0010111000001100;
            14'h0eff 	:	o_val <= 16'b0010111000001111;
            14'h0f00 	:	o_val <= 16'b0010111000010010;
            14'h0f01 	:	o_val <= 16'b0010111000010101;
            14'h0f02 	:	o_val <= 16'b0010111000011000;
            14'h0f03 	:	o_val <= 16'b0010111000011011;
            14'h0f04 	:	o_val <= 16'b0010111000011110;
            14'h0f05 	:	o_val <= 16'b0010111000100001;
            14'h0f06 	:	o_val <= 16'b0010111000100100;
            14'h0f07 	:	o_val <= 16'b0010111000100111;
            14'h0f08 	:	o_val <= 16'b0010111000101001;
            14'h0f09 	:	o_val <= 16'b0010111000101100;
            14'h0f0a 	:	o_val <= 16'b0010111000101111;
            14'h0f0b 	:	o_val <= 16'b0010111000110010;
            14'h0f0c 	:	o_val <= 16'b0010111000110101;
            14'h0f0d 	:	o_val <= 16'b0010111000111000;
            14'h0f0e 	:	o_val <= 16'b0010111000111011;
            14'h0f0f 	:	o_val <= 16'b0010111000111110;
            14'h0f10 	:	o_val <= 16'b0010111001000001;
            14'h0f11 	:	o_val <= 16'b0010111001000100;
            14'h0f12 	:	o_val <= 16'b0010111001000111;
            14'h0f13 	:	o_val <= 16'b0010111001001010;
            14'h0f14 	:	o_val <= 16'b0010111001001101;
            14'h0f15 	:	o_val <= 16'b0010111001010000;
            14'h0f16 	:	o_val <= 16'b0010111001010010;
            14'h0f17 	:	o_val <= 16'b0010111001010101;
            14'h0f18 	:	o_val <= 16'b0010111001011000;
            14'h0f19 	:	o_val <= 16'b0010111001011011;
            14'h0f1a 	:	o_val <= 16'b0010111001011110;
            14'h0f1b 	:	o_val <= 16'b0010111001100001;
            14'h0f1c 	:	o_val <= 16'b0010111001100100;
            14'h0f1d 	:	o_val <= 16'b0010111001100111;
            14'h0f1e 	:	o_val <= 16'b0010111001101010;
            14'h0f1f 	:	o_val <= 16'b0010111001101101;
            14'h0f20 	:	o_val <= 16'b0010111001110000;
            14'h0f21 	:	o_val <= 16'b0010111001110011;
            14'h0f22 	:	o_val <= 16'b0010111001110110;
            14'h0f23 	:	o_val <= 16'b0010111001111001;
            14'h0f24 	:	o_val <= 16'b0010111001111011;
            14'h0f25 	:	o_val <= 16'b0010111001111110;
            14'h0f26 	:	o_val <= 16'b0010111010000001;
            14'h0f27 	:	o_val <= 16'b0010111010000100;
            14'h0f28 	:	o_val <= 16'b0010111010000111;
            14'h0f29 	:	o_val <= 16'b0010111010001010;
            14'h0f2a 	:	o_val <= 16'b0010111010001101;
            14'h0f2b 	:	o_val <= 16'b0010111010010000;
            14'h0f2c 	:	o_val <= 16'b0010111010010011;
            14'h0f2d 	:	o_val <= 16'b0010111010010110;
            14'h0f2e 	:	o_val <= 16'b0010111010011001;
            14'h0f2f 	:	o_val <= 16'b0010111010011100;
            14'h0f30 	:	o_val <= 16'b0010111010011111;
            14'h0f31 	:	o_val <= 16'b0010111010100001;
            14'h0f32 	:	o_val <= 16'b0010111010100100;
            14'h0f33 	:	o_val <= 16'b0010111010100111;
            14'h0f34 	:	o_val <= 16'b0010111010101010;
            14'h0f35 	:	o_val <= 16'b0010111010101101;
            14'h0f36 	:	o_val <= 16'b0010111010110000;
            14'h0f37 	:	o_val <= 16'b0010111010110011;
            14'h0f38 	:	o_val <= 16'b0010111010110110;
            14'h0f39 	:	o_val <= 16'b0010111010111001;
            14'h0f3a 	:	o_val <= 16'b0010111010111100;
            14'h0f3b 	:	o_val <= 16'b0010111010111111;
            14'h0f3c 	:	o_val <= 16'b0010111011000010;
            14'h0f3d 	:	o_val <= 16'b0010111011000101;
            14'h0f3e 	:	o_val <= 16'b0010111011001000;
            14'h0f3f 	:	o_val <= 16'b0010111011001010;
            14'h0f40 	:	o_val <= 16'b0010111011001101;
            14'h0f41 	:	o_val <= 16'b0010111011010000;
            14'h0f42 	:	o_val <= 16'b0010111011010011;
            14'h0f43 	:	o_val <= 16'b0010111011010110;
            14'h0f44 	:	o_val <= 16'b0010111011011001;
            14'h0f45 	:	o_val <= 16'b0010111011011100;
            14'h0f46 	:	o_val <= 16'b0010111011011111;
            14'h0f47 	:	o_val <= 16'b0010111011100010;
            14'h0f48 	:	o_val <= 16'b0010111011100101;
            14'h0f49 	:	o_val <= 16'b0010111011101000;
            14'h0f4a 	:	o_val <= 16'b0010111011101011;
            14'h0f4b 	:	o_val <= 16'b0010111011101110;
            14'h0f4c 	:	o_val <= 16'b0010111011110000;
            14'h0f4d 	:	o_val <= 16'b0010111011110011;
            14'h0f4e 	:	o_val <= 16'b0010111011110110;
            14'h0f4f 	:	o_val <= 16'b0010111011111001;
            14'h0f50 	:	o_val <= 16'b0010111011111100;
            14'h0f51 	:	o_val <= 16'b0010111011111111;
            14'h0f52 	:	o_val <= 16'b0010111100000010;
            14'h0f53 	:	o_val <= 16'b0010111100000101;
            14'h0f54 	:	o_val <= 16'b0010111100001000;
            14'h0f55 	:	o_val <= 16'b0010111100001011;
            14'h0f56 	:	o_val <= 16'b0010111100001110;
            14'h0f57 	:	o_val <= 16'b0010111100010001;
            14'h0f58 	:	o_val <= 16'b0010111100010100;
            14'h0f59 	:	o_val <= 16'b0010111100010110;
            14'h0f5a 	:	o_val <= 16'b0010111100011001;
            14'h0f5b 	:	o_val <= 16'b0010111100011100;
            14'h0f5c 	:	o_val <= 16'b0010111100011111;
            14'h0f5d 	:	o_val <= 16'b0010111100100010;
            14'h0f5e 	:	o_val <= 16'b0010111100100101;
            14'h0f5f 	:	o_val <= 16'b0010111100101000;
            14'h0f60 	:	o_val <= 16'b0010111100101011;
            14'h0f61 	:	o_val <= 16'b0010111100101110;
            14'h0f62 	:	o_val <= 16'b0010111100110001;
            14'h0f63 	:	o_val <= 16'b0010111100110100;
            14'h0f64 	:	o_val <= 16'b0010111100110111;
            14'h0f65 	:	o_val <= 16'b0010111100111001;
            14'h0f66 	:	o_val <= 16'b0010111100111100;
            14'h0f67 	:	o_val <= 16'b0010111100111111;
            14'h0f68 	:	o_val <= 16'b0010111101000010;
            14'h0f69 	:	o_val <= 16'b0010111101000101;
            14'h0f6a 	:	o_val <= 16'b0010111101001000;
            14'h0f6b 	:	o_val <= 16'b0010111101001011;
            14'h0f6c 	:	o_val <= 16'b0010111101001110;
            14'h0f6d 	:	o_val <= 16'b0010111101010001;
            14'h0f6e 	:	o_val <= 16'b0010111101010100;
            14'h0f6f 	:	o_val <= 16'b0010111101010111;
            14'h0f70 	:	o_val <= 16'b0010111101011010;
            14'h0f71 	:	o_val <= 16'b0010111101011101;
            14'h0f72 	:	o_val <= 16'b0010111101011111;
            14'h0f73 	:	o_val <= 16'b0010111101100010;
            14'h0f74 	:	o_val <= 16'b0010111101100101;
            14'h0f75 	:	o_val <= 16'b0010111101101000;
            14'h0f76 	:	o_val <= 16'b0010111101101011;
            14'h0f77 	:	o_val <= 16'b0010111101101110;
            14'h0f78 	:	o_val <= 16'b0010111101110001;
            14'h0f79 	:	o_val <= 16'b0010111101110100;
            14'h0f7a 	:	o_val <= 16'b0010111101110111;
            14'h0f7b 	:	o_val <= 16'b0010111101111010;
            14'h0f7c 	:	o_val <= 16'b0010111101111101;
            14'h0f7d 	:	o_val <= 16'b0010111110000000;
            14'h0f7e 	:	o_val <= 16'b0010111110000010;
            14'h0f7f 	:	o_val <= 16'b0010111110000101;
            14'h0f80 	:	o_val <= 16'b0010111110001000;
            14'h0f81 	:	o_val <= 16'b0010111110001011;
            14'h0f82 	:	o_val <= 16'b0010111110001110;
            14'h0f83 	:	o_val <= 16'b0010111110010001;
            14'h0f84 	:	o_val <= 16'b0010111110010100;
            14'h0f85 	:	o_val <= 16'b0010111110010111;
            14'h0f86 	:	o_val <= 16'b0010111110011010;
            14'h0f87 	:	o_val <= 16'b0010111110011101;
            14'h0f88 	:	o_val <= 16'b0010111110100000;
            14'h0f89 	:	o_val <= 16'b0010111110100011;
            14'h0f8a 	:	o_val <= 16'b0010111110100101;
            14'h0f8b 	:	o_val <= 16'b0010111110101000;
            14'h0f8c 	:	o_val <= 16'b0010111110101011;
            14'h0f8d 	:	o_val <= 16'b0010111110101110;
            14'h0f8e 	:	o_val <= 16'b0010111110110001;
            14'h0f8f 	:	o_val <= 16'b0010111110110100;
            14'h0f90 	:	o_val <= 16'b0010111110110111;
            14'h0f91 	:	o_val <= 16'b0010111110111010;
            14'h0f92 	:	o_val <= 16'b0010111110111101;
            14'h0f93 	:	o_val <= 16'b0010111111000000;
            14'h0f94 	:	o_val <= 16'b0010111111000011;
            14'h0f95 	:	o_val <= 16'b0010111111000110;
            14'h0f96 	:	o_val <= 16'b0010111111001000;
            14'h0f97 	:	o_val <= 16'b0010111111001011;
            14'h0f98 	:	o_val <= 16'b0010111111001110;
            14'h0f99 	:	o_val <= 16'b0010111111010001;
            14'h0f9a 	:	o_val <= 16'b0010111111010100;
            14'h0f9b 	:	o_val <= 16'b0010111111010111;
            14'h0f9c 	:	o_val <= 16'b0010111111011010;
            14'h0f9d 	:	o_val <= 16'b0010111111011101;
            14'h0f9e 	:	o_val <= 16'b0010111111100000;
            14'h0f9f 	:	o_val <= 16'b0010111111100011;
            14'h0fa0 	:	o_val <= 16'b0010111111100110;
            14'h0fa1 	:	o_val <= 16'b0010111111101000;
            14'h0fa2 	:	o_val <= 16'b0010111111101011;
            14'h0fa3 	:	o_val <= 16'b0010111111101110;
            14'h0fa4 	:	o_val <= 16'b0010111111110001;
            14'h0fa5 	:	o_val <= 16'b0010111111110100;
            14'h0fa6 	:	o_val <= 16'b0010111111110111;
            14'h0fa7 	:	o_val <= 16'b0010111111111010;
            14'h0fa8 	:	o_val <= 16'b0010111111111101;
            14'h0fa9 	:	o_val <= 16'b0011000000000000;
            14'h0faa 	:	o_val <= 16'b0011000000000011;
            14'h0fab 	:	o_val <= 16'b0011000000000110;
            14'h0fac 	:	o_val <= 16'b0011000000001001;
            14'h0fad 	:	o_val <= 16'b0011000000001011;
            14'h0fae 	:	o_val <= 16'b0011000000001110;
            14'h0faf 	:	o_val <= 16'b0011000000010001;
            14'h0fb0 	:	o_val <= 16'b0011000000010100;
            14'h0fb1 	:	o_val <= 16'b0011000000010111;
            14'h0fb2 	:	o_val <= 16'b0011000000011010;
            14'h0fb3 	:	o_val <= 16'b0011000000011101;
            14'h0fb4 	:	o_val <= 16'b0011000000100000;
            14'h0fb5 	:	o_val <= 16'b0011000000100011;
            14'h0fb6 	:	o_val <= 16'b0011000000100110;
            14'h0fb7 	:	o_val <= 16'b0011000000101001;
            14'h0fb8 	:	o_val <= 16'b0011000000101011;
            14'h0fb9 	:	o_val <= 16'b0011000000101110;
            14'h0fba 	:	o_val <= 16'b0011000000110001;
            14'h0fbb 	:	o_val <= 16'b0011000000110100;
            14'h0fbc 	:	o_val <= 16'b0011000000110111;
            14'h0fbd 	:	o_val <= 16'b0011000000111010;
            14'h0fbe 	:	o_val <= 16'b0011000000111101;
            14'h0fbf 	:	o_val <= 16'b0011000001000000;
            14'h0fc0 	:	o_val <= 16'b0011000001000011;
            14'h0fc1 	:	o_val <= 16'b0011000001000110;
            14'h0fc2 	:	o_val <= 16'b0011000001001001;
            14'h0fc3 	:	o_val <= 16'b0011000001001011;
            14'h0fc4 	:	o_val <= 16'b0011000001001110;
            14'h0fc5 	:	o_val <= 16'b0011000001010001;
            14'h0fc6 	:	o_val <= 16'b0011000001010100;
            14'h0fc7 	:	o_val <= 16'b0011000001010111;
            14'h0fc8 	:	o_val <= 16'b0011000001011010;
            14'h0fc9 	:	o_val <= 16'b0011000001011101;
            14'h0fca 	:	o_val <= 16'b0011000001100000;
            14'h0fcb 	:	o_val <= 16'b0011000001100011;
            14'h0fcc 	:	o_val <= 16'b0011000001100110;
            14'h0fcd 	:	o_val <= 16'b0011000001101001;
            14'h0fce 	:	o_val <= 16'b0011000001101011;
            14'h0fcf 	:	o_val <= 16'b0011000001101110;
            14'h0fd0 	:	o_val <= 16'b0011000001110001;
            14'h0fd1 	:	o_val <= 16'b0011000001110100;
            14'h0fd2 	:	o_val <= 16'b0011000001110111;
            14'h0fd3 	:	o_val <= 16'b0011000001111010;
            14'h0fd4 	:	o_val <= 16'b0011000001111101;
            14'h0fd5 	:	o_val <= 16'b0011000010000000;
            14'h0fd6 	:	o_val <= 16'b0011000010000011;
            14'h0fd7 	:	o_val <= 16'b0011000010000110;
            14'h0fd8 	:	o_val <= 16'b0011000010001001;
            14'h0fd9 	:	o_val <= 16'b0011000010001011;
            14'h0fda 	:	o_val <= 16'b0011000010001110;
            14'h0fdb 	:	o_val <= 16'b0011000010010001;
            14'h0fdc 	:	o_val <= 16'b0011000010010100;
            14'h0fdd 	:	o_val <= 16'b0011000010010111;
            14'h0fde 	:	o_val <= 16'b0011000010011010;
            14'h0fdf 	:	o_val <= 16'b0011000010011101;
            14'h0fe0 	:	o_val <= 16'b0011000010100000;
            14'h0fe1 	:	o_val <= 16'b0011000010100011;
            14'h0fe2 	:	o_val <= 16'b0011000010100110;
            14'h0fe3 	:	o_val <= 16'b0011000010101001;
            14'h0fe4 	:	o_val <= 16'b0011000010101011;
            14'h0fe5 	:	o_val <= 16'b0011000010101110;
            14'h0fe6 	:	o_val <= 16'b0011000010110001;
            14'h0fe7 	:	o_val <= 16'b0011000010110100;
            14'h0fe8 	:	o_val <= 16'b0011000010110111;
            14'h0fe9 	:	o_val <= 16'b0011000010111010;
            14'h0fea 	:	o_val <= 16'b0011000010111101;
            14'h0feb 	:	o_val <= 16'b0011000011000000;
            14'h0fec 	:	o_val <= 16'b0011000011000011;
            14'h0fed 	:	o_val <= 16'b0011000011000110;
            14'h0fee 	:	o_val <= 16'b0011000011001000;
            14'h0fef 	:	o_val <= 16'b0011000011001011;
            14'h0ff0 	:	o_val <= 16'b0011000011001110;
            14'h0ff1 	:	o_val <= 16'b0011000011010001;
            14'h0ff2 	:	o_val <= 16'b0011000011010100;
            14'h0ff3 	:	o_val <= 16'b0011000011010111;
            14'h0ff4 	:	o_val <= 16'b0011000011011010;
            14'h0ff5 	:	o_val <= 16'b0011000011011101;
            14'h0ff6 	:	o_val <= 16'b0011000011100000;
            14'h0ff7 	:	o_val <= 16'b0011000011100011;
            14'h0ff8 	:	o_val <= 16'b0011000011100101;
            14'h0ff9 	:	o_val <= 16'b0011000011101000;
            14'h0ffa 	:	o_val <= 16'b0011000011101011;
            14'h0ffb 	:	o_val <= 16'b0011000011101110;
            14'h0ffc 	:	o_val <= 16'b0011000011110001;
            14'h0ffd 	:	o_val <= 16'b0011000011110100;
            14'h0ffe 	:	o_val <= 16'b0011000011110111;
            14'h0fff 	:	o_val <= 16'b0011000011111010;
            14'h1000 	:	o_val <= 16'b0011000011111101;
            14'h1001 	:	o_val <= 16'b0011000100000000;
            14'h1002 	:	o_val <= 16'b0011000100000011;
            14'h1003 	:	o_val <= 16'b0011000100000101;
            14'h1004 	:	o_val <= 16'b0011000100001000;
            14'h1005 	:	o_val <= 16'b0011000100001011;
            14'h1006 	:	o_val <= 16'b0011000100001110;
            14'h1007 	:	o_val <= 16'b0011000100010001;
            14'h1008 	:	o_val <= 16'b0011000100010100;
            14'h1009 	:	o_val <= 16'b0011000100010111;
            14'h100a 	:	o_val <= 16'b0011000100011010;
            14'h100b 	:	o_val <= 16'b0011000100011101;
            14'h100c 	:	o_val <= 16'b0011000100100000;
            14'h100d 	:	o_val <= 16'b0011000100100010;
            14'h100e 	:	o_val <= 16'b0011000100100101;
            14'h100f 	:	o_val <= 16'b0011000100101000;
            14'h1010 	:	o_val <= 16'b0011000100101011;
            14'h1011 	:	o_val <= 16'b0011000100101110;
            14'h1012 	:	o_val <= 16'b0011000100110001;
            14'h1013 	:	o_val <= 16'b0011000100110100;
            14'h1014 	:	o_val <= 16'b0011000100110111;
            14'h1015 	:	o_val <= 16'b0011000100111010;
            14'h1016 	:	o_val <= 16'b0011000100111101;
            14'h1017 	:	o_val <= 16'b0011000100111111;
            14'h1018 	:	o_val <= 16'b0011000101000010;
            14'h1019 	:	o_val <= 16'b0011000101000101;
            14'h101a 	:	o_val <= 16'b0011000101001000;
            14'h101b 	:	o_val <= 16'b0011000101001011;
            14'h101c 	:	o_val <= 16'b0011000101001110;
            14'h101d 	:	o_val <= 16'b0011000101010001;
            14'h101e 	:	o_val <= 16'b0011000101010100;
            14'h101f 	:	o_val <= 16'b0011000101010111;
            14'h1020 	:	o_val <= 16'b0011000101011010;
            14'h1021 	:	o_val <= 16'b0011000101011100;
            14'h1022 	:	o_val <= 16'b0011000101011111;
            14'h1023 	:	o_val <= 16'b0011000101100010;
            14'h1024 	:	o_val <= 16'b0011000101100101;
            14'h1025 	:	o_val <= 16'b0011000101101000;
            14'h1026 	:	o_val <= 16'b0011000101101011;
            14'h1027 	:	o_val <= 16'b0011000101101110;
            14'h1028 	:	o_val <= 16'b0011000101110001;
            14'h1029 	:	o_val <= 16'b0011000101110100;
            14'h102a 	:	o_val <= 16'b0011000101110111;
            14'h102b 	:	o_val <= 16'b0011000101111001;
            14'h102c 	:	o_val <= 16'b0011000101111100;
            14'h102d 	:	o_val <= 16'b0011000101111111;
            14'h102e 	:	o_val <= 16'b0011000110000010;
            14'h102f 	:	o_val <= 16'b0011000110000101;
            14'h1030 	:	o_val <= 16'b0011000110001000;
            14'h1031 	:	o_val <= 16'b0011000110001011;
            14'h1032 	:	o_val <= 16'b0011000110001110;
            14'h1033 	:	o_val <= 16'b0011000110010001;
            14'h1034 	:	o_val <= 16'b0011000110010011;
            14'h1035 	:	o_val <= 16'b0011000110010110;
            14'h1036 	:	o_val <= 16'b0011000110011001;
            14'h1037 	:	o_val <= 16'b0011000110011100;
            14'h1038 	:	o_val <= 16'b0011000110011111;
            14'h1039 	:	o_val <= 16'b0011000110100010;
            14'h103a 	:	o_val <= 16'b0011000110100101;
            14'h103b 	:	o_val <= 16'b0011000110101000;
            14'h103c 	:	o_val <= 16'b0011000110101011;
            14'h103d 	:	o_val <= 16'b0011000110101110;
            14'h103e 	:	o_val <= 16'b0011000110110000;
            14'h103f 	:	o_val <= 16'b0011000110110011;
            14'h1040 	:	o_val <= 16'b0011000110110110;
            14'h1041 	:	o_val <= 16'b0011000110111001;
            14'h1042 	:	o_val <= 16'b0011000110111100;
            14'h1043 	:	o_val <= 16'b0011000110111111;
            14'h1044 	:	o_val <= 16'b0011000111000010;
            14'h1045 	:	o_val <= 16'b0011000111000101;
            14'h1046 	:	o_val <= 16'b0011000111001000;
            14'h1047 	:	o_val <= 16'b0011000111001010;
            14'h1048 	:	o_val <= 16'b0011000111001101;
            14'h1049 	:	o_val <= 16'b0011000111010000;
            14'h104a 	:	o_val <= 16'b0011000111010011;
            14'h104b 	:	o_val <= 16'b0011000111010110;
            14'h104c 	:	o_val <= 16'b0011000111011001;
            14'h104d 	:	o_val <= 16'b0011000111011100;
            14'h104e 	:	o_val <= 16'b0011000111011111;
            14'h104f 	:	o_val <= 16'b0011000111100010;
            14'h1050 	:	o_val <= 16'b0011000111100101;
            14'h1051 	:	o_val <= 16'b0011000111100111;
            14'h1052 	:	o_val <= 16'b0011000111101010;
            14'h1053 	:	o_val <= 16'b0011000111101101;
            14'h1054 	:	o_val <= 16'b0011000111110000;
            14'h1055 	:	o_val <= 16'b0011000111110011;
            14'h1056 	:	o_val <= 16'b0011000111110110;
            14'h1057 	:	o_val <= 16'b0011000111111001;
            14'h1058 	:	o_val <= 16'b0011000111111100;
            14'h1059 	:	o_val <= 16'b0011000111111111;
            14'h105a 	:	o_val <= 16'b0011001000000001;
            14'h105b 	:	o_val <= 16'b0011001000000100;
            14'h105c 	:	o_val <= 16'b0011001000000111;
            14'h105d 	:	o_val <= 16'b0011001000001010;
            14'h105e 	:	o_val <= 16'b0011001000001101;
            14'h105f 	:	o_val <= 16'b0011001000010000;
            14'h1060 	:	o_val <= 16'b0011001000010011;
            14'h1061 	:	o_val <= 16'b0011001000010110;
            14'h1062 	:	o_val <= 16'b0011001000011001;
            14'h1063 	:	o_val <= 16'b0011001000011011;
            14'h1064 	:	o_val <= 16'b0011001000011110;
            14'h1065 	:	o_val <= 16'b0011001000100001;
            14'h1066 	:	o_val <= 16'b0011001000100100;
            14'h1067 	:	o_val <= 16'b0011001000100111;
            14'h1068 	:	o_val <= 16'b0011001000101010;
            14'h1069 	:	o_val <= 16'b0011001000101101;
            14'h106a 	:	o_val <= 16'b0011001000110000;
            14'h106b 	:	o_val <= 16'b0011001000110011;
            14'h106c 	:	o_val <= 16'b0011001000110110;
            14'h106d 	:	o_val <= 16'b0011001000111000;
            14'h106e 	:	o_val <= 16'b0011001000111011;
            14'h106f 	:	o_val <= 16'b0011001000111110;
            14'h1070 	:	o_val <= 16'b0011001001000001;
            14'h1071 	:	o_val <= 16'b0011001001000100;
            14'h1072 	:	o_val <= 16'b0011001001000111;
            14'h1073 	:	o_val <= 16'b0011001001001010;
            14'h1074 	:	o_val <= 16'b0011001001001101;
            14'h1075 	:	o_val <= 16'b0011001001010000;
            14'h1076 	:	o_val <= 16'b0011001001010010;
            14'h1077 	:	o_val <= 16'b0011001001010101;
            14'h1078 	:	o_val <= 16'b0011001001011000;
            14'h1079 	:	o_val <= 16'b0011001001011011;
            14'h107a 	:	o_val <= 16'b0011001001011110;
            14'h107b 	:	o_val <= 16'b0011001001100001;
            14'h107c 	:	o_val <= 16'b0011001001100100;
            14'h107d 	:	o_val <= 16'b0011001001100111;
            14'h107e 	:	o_val <= 16'b0011001001101001;
            14'h107f 	:	o_val <= 16'b0011001001101100;
            14'h1080 	:	o_val <= 16'b0011001001101111;
            14'h1081 	:	o_val <= 16'b0011001001110010;
            14'h1082 	:	o_val <= 16'b0011001001110101;
            14'h1083 	:	o_val <= 16'b0011001001111000;
            14'h1084 	:	o_val <= 16'b0011001001111011;
            14'h1085 	:	o_val <= 16'b0011001001111110;
            14'h1086 	:	o_val <= 16'b0011001010000001;
            14'h1087 	:	o_val <= 16'b0011001010000011;
            14'h1088 	:	o_val <= 16'b0011001010000110;
            14'h1089 	:	o_val <= 16'b0011001010001001;
            14'h108a 	:	o_val <= 16'b0011001010001100;
            14'h108b 	:	o_val <= 16'b0011001010001111;
            14'h108c 	:	o_val <= 16'b0011001010010010;
            14'h108d 	:	o_val <= 16'b0011001010010101;
            14'h108e 	:	o_val <= 16'b0011001010011000;
            14'h108f 	:	o_val <= 16'b0011001010011011;
            14'h1090 	:	o_val <= 16'b0011001010011101;
            14'h1091 	:	o_val <= 16'b0011001010100000;
            14'h1092 	:	o_val <= 16'b0011001010100011;
            14'h1093 	:	o_val <= 16'b0011001010100110;
            14'h1094 	:	o_val <= 16'b0011001010101001;
            14'h1095 	:	o_val <= 16'b0011001010101100;
            14'h1096 	:	o_val <= 16'b0011001010101111;
            14'h1097 	:	o_val <= 16'b0011001010110010;
            14'h1098 	:	o_val <= 16'b0011001010110101;
            14'h1099 	:	o_val <= 16'b0011001010110111;
            14'h109a 	:	o_val <= 16'b0011001010111010;
            14'h109b 	:	o_val <= 16'b0011001010111101;
            14'h109c 	:	o_val <= 16'b0011001011000000;
            14'h109d 	:	o_val <= 16'b0011001011000011;
            14'h109e 	:	o_val <= 16'b0011001011000110;
            14'h109f 	:	o_val <= 16'b0011001011001001;
            14'h10a0 	:	o_val <= 16'b0011001011001100;
            14'h10a1 	:	o_val <= 16'b0011001011001110;
            14'h10a2 	:	o_val <= 16'b0011001011010001;
            14'h10a3 	:	o_val <= 16'b0011001011010100;
            14'h10a4 	:	o_val <= 16'b0011001011010111;
            14'h10a5 	:	o_val <= 16'b0011001011011010;
            14'h10a6 	:	o_val <= 16'b0011001011011101;
            14'h10a7 	:	o_val <= 16'b0011001011100000;
            14'h10a8 	:	o_val <= 16'b0011001011100011;
            14'h10a9 	:	o_val <= 16'b0011001011100110;
            14'h10aa 	:	o_val <= 16'b0011001011101000;
            14'h10ab 	:	o_val <= 16'b0011001011101011;
            14'h10ac 	:	o_val <= 16'b0011001011101110;
            14'h10ad 	:	o_val <= 16'b0011001011110001;
            14'h10ae 	:	o_val <= 16'b0011001011110100;
            14'h10af 	:	o_val <= 16'b0011001011110111;
            14'h10b0 	:	o_val <= 16'b0011001011111010;
            14'h10b1 	:	o_val <= 16'b0011001011111101;
            14'h10b2 	:	o_val <= 16'b0011001011111111;
            14'h10b3 	:	o_val <= 16'b0011001100000010;
            14'h10b4 	:	o_val <= 16'b0011001100000101;
            14'h10b5 	:	o_val <= 16'b0011001100001000;
            14'h10b6 	:	o_val <= 16'b0011001100001011;
            14'h10b7 	:	o_val <= 16'b0011001100001110;
            14'h10b8 	:	o_val <= 16'b0011001100010001;
            14'h10b9 	:	o_val <= 16'b0011001100010100;
            14'h10ba 	:	o_val <= 16'b0011001100010111;
            14'h10bb 	:	o_val <= 16'b0011001100011001;
            14'h10bc 	:	o_val <= 16'b0011001100011100;
            14'h10bd 	:	o_val <= 16'b0011001100011111;
            14'h10be 	:	o_val <= 16'b0011001100100010;
            14'h10bf 	:	o_val <= 16'b0011001100100101;
            14'h10c0 	:	o_val <= 16'b0011001100101000;
            14'h10c1 	:	o_val <= 16'b0011001100101011;
            14'h10c2 	:	o_val <= 16'b0011001100101110;
            14'h10c3 	:	o_val <= 16'b0011001100110000;
            14'h10c4 	:	o_val <= 16'b0011001100110011;
            14'h10c5 	:	o_val <= 16'b0011001100110110;
            14'h10c6 	:	o_val <= 16'b0011001100111001;
            14'h10c7 	:	o_val <= 16'b0011001100111100;
            14'h10c8 	:	o_val <= 16'b0011001100111111;
            14'h10c9 	:	o_val <= 16'b0011001101000010;
            14'h10ca 	:	o_val <= 16'b0011001101000101;
            14'h10cb 	:	o_val <= 16'b0011001101000111;
            14'h10cc 	:	o_val <= 16'b0011001101001010;
            14'h10cd 	:	o_val <= 16'b0011001101001101;
            14'h10ce 	:	o_val <= 16'b0011001101010000;
            14'h10cf 	:	o_val <= 16'b0011001101010011;
            14'h10d0 	:	o_val <= 16'b0011001101010110;
            14'h10d1 	:	o_val <= 16'b0011001101011001;
            14'h10d2 	:	o_val <= 16'b0011001101011100;
            14'h10d3 	:	o_val <= 16'b0011001101011111;
            14'h10d4 	:	o_val <= 16'b0011001101100001;
            14'h10d5 	:	o_val <= 16'b0011001101100100;
            14'h10d6 	:	o_val <= 16'b0011001101100111;
            14'h10d7 	:	o_val <= 16'b0011001101101010;
            14'h10d8 	:	o_val <= 16'b0011001101101101;
            14'h10d9 	:	o_val <= 16'b0011001101110000;
            14'h10da 	:	o_val <= 16'b0011001101110011;
            14'h10db 	:	o_val <= 16'b0011001101110110;
            14'h10dc 	:	o_val <= 16'b0011001101111000;
            14'h10dd 	:	o_val <= 16'b0011001101111011;
            14'h10de 	:	o_val <= 16'b0011001101111110;
            14'h10df 	:	o_val <= 16'b0011001110000001;
            14'h10e0 	:	o_val <= 16'b0011001110000100;
            14'h10e1 	:	o_val <= 16'b0011001110000111;
            14'h10e2 	:	o_val <= 16'b0011001110001010;
            14'h10e3 	:	o_val <= 16'b0011001110001101;
            14'h10e4 	:	o_val <= 16'b0011001110001111;
            14'h10e5 	:	o_val <= 16'b0011001110010010;
            14'h10e6 	:	o_val <= 16'b0011001110010101;
            14'h10e7 	:	o_val <= 16'b0011001110011000;
            14'h10e8 	:	o_val <= 16'b0011001110011011;
            14'h10e9 	:	o_val <= 16'b0011001110011110;
            14'h10ea 	:	o_val <= 16'b0011001110100001;
            14'h10eb 	:	o_val <= 16'b0011001110100100;
            14'h10ec 	:	o_val <= 16'b0011001110100110;
            14'h10ed 	:	o_val <= 16'b0011001110101001;
            14'h10ee 	:	o_val <= 16'b0011001110101100;
            14'h10ef 	:	o_val <= 16'b0011001110101111;
            14'h10f0 	:	o_val <= 16'b0011001110110010;
            14'h10f1 	:	o_val <= 16'b0011001110110101;
            14'h10f2 	:	o_val <= 16'b0011001110111000;
            14'h10f3 	:	o_val <= 16'b0011001110111011;
            14'h10f4 	:	o_val <= 16'b0011001110111101;
            14'h10f5 	:	o_val <= 16'b0011001111000000;
            14'h10f6 	:	o_val <= 16'b0011001111000011;
            14'h10f7 	:	o_val <= 16'b0011001111000110;
            14'h10f8 	:	o_val <= 16'b0011001111001001;
            14'h10f9 	:	o_val <= 16'b0011001111001100;
            14'h10fa 	:	o_val <= 16'b0011001111001111;
            14'h10fb 	:	o_val <= 16'b0011001111010010;
            14'h10fc 	:	o_val <= 16'b0011001111010100;
            14'h10fd 	:	o_val <= 16'b0011001111010111;
            14'h10fe 	:	o_val <= 16'b0011001111011010;
            14'h10ff 	:	o_val <= 16'b0011001111011101;
            14'h1100 	:	o_val <= 16'b0011001111100000;
            14'h1101 	:	o_val <= 16'b0011001111100011;
            14'h1102 	:	o_val <= 16'b0011001111100110;
            14'h1103 	:	o_val <= 16'b0011001111101000;
            14'h1104 	:	o_val <= 16'b0011001111101011;
            14'h1105 	:	o_val <= 16'b0011001111101110;
            14'h1106 	:	o_val <= 16'b0011001111110001;
            14'h1107 	:	o_val <= 16'b0011001111110100;
            14'h1108 	:	o_val <= 16'b0011001111110111;
            14'h1109 	:	o_val <= 16'b0011001111111010;
            14'h110a 	:	o_val <= 16'b0011001111111101;
            14'h110b 	:	o_val <= 16'b0011001111111111;
            14'h110c 	:	o_val <= 16'b0011010000000010;
            14'h110d 	:	o_val <= 16'b0011010000000101;
            14'h110e 	:	o_val <= 16'b0011010000001000;
            14'h110f 	:	o_val <= 16'b0011010000001011;
            14'h1110 	:	o_val <= 16'b0011010000001110;
            14'h1111 	:	o_val <= 16'b0011010000010001;
            14'h1112 	:	o_val <= 16'b0011010000010100;
            14'h1113 	:	o_val <= 16'b0011010000010110;
            14'h1114 	:	o_val <= 16'b0011010000011001;
            14'h1115 	:	o_val <= 16'b0011010000011100;
            14'h1116 	:	o_val <= 16'b0011010000011111;
            14'h1117 	:	o_val <= 16'b0011010000100010;
            14'h1118 	:	o_val <= 16'b0011010000100101;
            14'h1119 	:	o_val <= 16'b0011010000101000;
            14'h111a 	:	o_val <= 16'b0011010000101011;
            14'h111b 	:	o_val <= 16'b0011010000101101;
            14'h111c 	:	o_val <= 16'b0011010000110000;
            14'h111d 	:	o_val <= 16'b0011010000110011;
            14'h111e 	:	o_val <= 16'b0011010000110110;
            14'h111f 	:	o_val <= 16'b0011010000111001;
            14'h1120 	:	o_val <= 16'b0011010000111100;
            14'h1121 	:	o_val <= 16'b0011010000111111;
            14'h1122 	:	o_val <= 16'b0011010001000001;
            14'h1123 	:	o_val <= 16'b0011010001000100;
            14'h1124 	:	o_val <= 16'b0011010001000111;
            14'h1125 	:	o_val <= 16'b0011010001001010;
            14'h1126 	:	o_val <= 16'b0011010001001101;
            14'h1127 	:	o_val <= 16'b0011010001010000;
            14'h1128 	:	o_val <= 16'b0011010001010011;
            14'h1129 	:	o_val <= 16'b0011010001010110;
            14'h112a 	:	o_val <= 16'b0011010001011000;
            14'h112b 	:	o_val <= 16'b0011010001011011;
            14'h112c 	:	o_val <= 16'b0011010001011110;
            14'h112d 	:	o_val <= 16'b0011010001100001;
            14'h112e 	:	o_val <= 16'b0011010001100100;
            14'h112f 	:	o_val <= 16'b0011010001100111;
            14'h1130 	:	o_val <= 16'b0011010001101010;
            14'h1131 	:	o_val <= 16'b0011010001101100;
            14'h1132 	:	o_val <= 16'b0011010001101111;
            14'h1133 	:	o_val <= 16'b0011010001110010;
            14'h1134 	:	o_val <= 16'b0011010001110101;
            14'h1135 	:	o_val <= 16'b0011010001111000;
            14'h1136 	:	o_val <= 16'b0011010001111011;
            14'h1137 	:	o_val <= 16'b0011010001111110;
            14'h1138 	:	o_val <= 16'b0011010010000001;
            14'h1139 	:	o_val <= 16'b0011010010000011;
            14'h113a 	:	o_val <= 16'b0011010010000110;
            14'h113b 	:	o_val <= 16'b0011010010001001;
            14'h113c 	:	o_val <= 16'b0011010010001100;
            14'h113d 	:	o_val <= 16'b0011010010001111;
            14'h113e 	:	o_val <= 16'b0011010010010010;
            14'h113f 	:	o_val <= 16'b0011010010010101;
            14'h1140 	:	o_val <= 16'b0011010010010111;
            14'h1141 	:	o_val <= 16'b0011010010011010;
            14'h1142 	:	o_val <= 16'b0011010010011101;
            14'h1143 	:	o_val <= 16'b0011010010100000;
            14'h1144 	:	o_val <= 16'b0011010010100011;
            14'h1145 	:	o_val <= 16'b0011010010100110;
            14'h1146 	:	o_val <= 16'b0011010010101001;
            14'h1147 	:	o_val <= 16'b0011010010101011;
            14'h1148 	:	o_val <= 16'b0011010010101110;
            14'h1149 	:	o_val <= 16'b0011010010110001;
            14'h114a 	:	o_val <= 16'b0011010010110100;
            14'h114b 	:	o_val <= 16'b0011010010110111;
            14'h114c 	:	o_val <= 16'b0011010010111010;
            14'h114d 	:	o_val <= 16'b0011010010111101;
            14'h114e 	:	o_val <= 16'b0011010011000000;
            14'h114f 	:	o_val <= 16'b0011010011000010;
            14'h1150 	:	o_val <= 16'b0011010011000101;
            14'h1151 	:	o_val <= 16'b0011010011001000;
            14'h1152 	:	o_val <= 16'b0011010011001011;
            14'h1153 	:	o_val <= 16'b0011010011001110;
            14'h1154 	:	o_val <= 16'b0011010011010001;
            14'h1155 	:	o_val <= 16'b0011010011010100;
            14'h1156 	:	o_val <= 16'b0011010011010110;
            14'h1157 	:	o_val <= 16'b0011010011011001;
            14'h1158 	:	o_val <= 16'b0011010011011100;
            14'h1159 	:	o_val <= 16'b0011010011011111;
            14'h115a 	:	o_val <= 16'b0011010011100010;
            14'h115b 	:	o_val <= 16'b0011010011100101;
            14'h115c 	:	o_val <= 16'b0011010011101000;
            14'h115d 	:	o_val <= 16'b0011010011101010;
            14'h115e 	:	o_val <= 16'b0011010011101101;
            14'h115f 	:	o_val <= 16'b0011010011110000;
            14'h1160 	:	o_val <= 16'b0011010011110011;
            14'h1161 	:	o_val <= 16'b0011010011110110;
            14'h1162 	:	o_val <= 16'b0011010011111001;
            14'h1163 	:	o_val <= 16'b0011010011111100;
            14'h1164 	:	o_val <= 16'b0011010011111110;
            14'h1165 	:	o_val <= 16'b0011010100000001;
            14'h1166 	:	o_val <= 16'b0011010100000100;
            14'h1167 	:	o_val <= 16'b0011010100000111;
            14'h1168 	:	o_val <= 16'b0011010100001010;
            14'h1169 	:	o_val <= 16'b0011010100001101;
            14'h116a 	:	o_val <= 16'b0011010100010000;
            14'h116b 	:	o_val <= 16'b0011010100010010;
            14'h116c 	:	o_val <= 16'b0011010100010101;
            14'h116d 	:	o_val <= 16'b0011010100011000;
            14'h116e 	:	o_val <= 16'b0011010100011011;
            14'h116f 	:	o_val <= 16'b0011010100011110;
            14'h1170 	:	o_val <= 16'b0011010100100001;
            14'h1171 	:	o_val <= 16'b0011010100100100;
            14'h1172 	:	o_val <= 16'b0011010100100110;
            14'h1173 	:	o_val <= 16'b0011010100101001;
            14'h1174 	:	o_val <= 16'b0011010100101100;
            14'h1175 	:	o_val <= 16'b0011010100101111;
            14'h1176 	:	o_val <= 16'b0011010100110010;
            14'h1177 	:	o_val <= 16'b0011010100110101;
            14'h1178 	:	o_val <= 16'b0011010100111000;
            14'h1179 	:	o_val <= 16'b0011010100111010;
            14'h117a 	:	o_val <= 16'b0011010100111101;
            14'h117b 	:	o_val <= 16'b0011010101000000;
            14'h117c 	:	o_val <= 16'b0011010101000011;
            14'h117d 	:	o_val <= 16'b0011010101000110;
            14'h117e 	:	o_val <= 16'b0011010101001001;
            14'h117f 	:	o_val <= 16'b0011010101001100;
            14'h1180 	:	o_val <= 16'b0011010101001110;
            14'h1181 	:	o_val <= 16'b0011010101010001;
            14'h1182 	:	o_val <= 16'b0011010101010100;
            14'h1183 	:	o_val <= 16'b0011010101010111;
            14'h1184 	:	o_val <= 16'b0011010101011010;
            14'h1185 	:	o_val <= 16'b0011010101011101;
            14'h1186 	:	o_val <= 16'b0011010101100000;
            14'h1187 	:	o_val <= 16'b0011010101100010;
            14'h1188 	:	o_val <= 16'b0011010101100101;
            14'h1189 	:	o_val <= 16'b0011010101101000;
            14'h118a 	:	o_val <= 16'b0011010101101011;
            14'h118b 	:	o_val <= 16'b0011010101101110;
            14'h118c 	:	o_val <= 16'b0011010101110001;
            14'h118d 	:	o_val <= 16'b0011010101110100;
            14'h118e 	:	o_val <= 16'b0011010101110110;
            14'h118f 	:	o_val <= 16'b0011010101111001;
            14'h1190 	:	o_val <= 16'b0011010101111100;
            14'h1191 	:	o_val <= 16'b0011010101111111;
            14'h1192 	:	o_val <= 16'b0011010110000010;
            14'h1193 	:	o_val <= 16'b0011010110000101;
            14'h1194 	:	o_val <= 16'b0011010110001000;
            14'h1195 	:	o_val <= 16'b0011010110001010;
            14'h1196 	:	o_val <= 16'b0011010110001101;
            14'h1197 	:	o_val <= 16'b0011010110010000;
            14'h1198 	:	o_val <= 16'b0011010110010011;
            14'h1199 	:	o_val <= 16'b0011010110010110;
            14'h119a 	:	o_val <= 16'b0011010110011001;
            14'h119b 	:	o_val <= 16'b0011010110011100;
            14'h119c 	:	o_val <= 16'b0011010110011110;
            14'h119d 	:	o_val <= 16'b0011010110100001;
            14'h119e 	:	o_val <= 16'b0011010110100100;
            14'h119f 	:	o_val <= 16'b0011010110100111;
            14'h11a0 	:	o_val <= 16'b0011010110101010;
            14'h11a1 	:	o_val <= 16'b0011010110101101;
            14'h11a2 	:	o_val <= 16'b0011010110110000;
            14'h11a3 	:	o_val <= 16'b0011010110110010;
            14'h11a4 	:	o_val <= 16'b0011010110110101;
            14'h11a5 	:	o_val <= 16'b0011010110111000;
            14'h11a6 	:	o_val <= 16'b0011010110111011;
            14'h11a7 	:	o_val <= 16'b0011010110111110;
            14'h11a8 	:	o_val <= 16'b0011010111000001;
            14'h11a9 	:	o_val <= 16'b0011010111000011;
            14'h11aa 	:	o_val <= 16'b0011010111000110;
            14'h11ab 	:	o_val <= 16'b0011010111001001;
            14'h11ac 	:	o_val <= 16'b0011010111001100;
            14'h11ad 	:	o_val <= 16'b0011010111001111;
            14'h11ae 	:	o_val <= 16'b0011010111010010;
            14'h11af 	:	o_val <= 16'b0011010111010101;
            14'h11b0 	:	o_val <= 16'b0011010111010111;
            14'h11b1 	:	o_val <= 16'b0011010111011010;
            14'h11b2 	:	o_val <= 16'b0011010111011101;
            14'h11b3 	:	o_val <= 16'b0011010111100000;
            14'h11b4 	:	o_val <= 16'b0011010111100011;
            14'h11b5 	:	o_val <= 16'b0011010111100110;
            14'h11b6 	:	o_val <= 16'b0011010111101001;
            14'h11b7 	:	o_val <= 16'b0011010111101011;
            14'h11b8 	:	o_val <= 16'b0011010111101110;
            14'h11b9 	:	o_val <= 16'b0011010111110001;
            14'h11ba 	:	o_val <= 16'b0011010111110100;
            14'h11bb 	:	o_val <= 16'b0011010111110111;
            14'h11bc 	:	o_val <= 16'b0011010111111010;
            14'h11bd 	:	o_val <= 16'b0011010111111100;
            14'h11be 	:	o_val <= 16'b0011010111111111;
            14'h11bf 	:	o_val <= 16'b0011011000000010;
            14'h11c0 	:	o_val <= 16'b0011011000000101;
            14'h11c1 	:	o_val <= 16'b0011011000001000;
            14'h11c2 	:	o_val <= 16'b0011011000001011;
            14'h11c3 	:	o_val <= 16'b0011011000001110;
            14'h11c4 	:	o_val <= 16'b0011011000010000;
            14'h11c5 	:	o_val <= 16'b0011011000010011;
            14'h11c6 	:	o_val <= 16'b0011011000010110;
            14'h11c7 	:	o_val <= 16'b0011011000011001;
            14'h11c8 	:	o_val <= 16'b0011011000011100;
            14'h11c9 	:	o_val <= 16'b0011011000011111;
            14'h11ca 	:	o_val <= 16'b0011011000100010;
            14'h11cb 	:	o_val <= 16'b0011011000100100;
            14'h11cc 	:	o_val <= 16'b0011011000100111;
            14'h11cd 	:	o_val <= 16'b0011011000101010;
            14'h11ce 	:	o_val <= 16'b0011011000101101;
            14'h11cf 	:	o_val <= 16'b0011011000110000;
            14'h11d0 	:	o_val <= 16'b0011011000110011;
            14'h11d1 	:	o_val <= 16'b0011011000110101;
            14'h11d2 	:	o_val <= 16'b0011011000111000;
            14'h11d3 	:	o_val <= 16'b0011011000111011;
            14'h11d4 	:	o_val <= 16'b0011011000111110;
            14'h11d5 	:	o_val <= 16'b0011011001000001;
            14'h11d6 	:	o_val <= 16'b0011011001000100;
            14'h11d7 	:	o_val <= 16'b0011011001000111;
            14'h11d8 	:	o_val <= 16'b0011011001001001;
            14'h11d9 	:	o_val <= 16'b0011011001001100;
            14'h11da 	:	o_val <= 16'b0011011001001111;
            14'h11db 	:	o_val <= 16'b0011011001010010;
            14'h11dc 	:	o_val <= 16'b0011011001010101;
            14'h11dd 	:	o_val <= 16'b0011011001011000;
            14'h11de 	:	o_val <= 16'b0011011001011010;
            14'h11df 	:	o_val <= 16'b0011011001011101;
            14'h11e0 	:	o_val <= 16'b0011011001100000;
            14'h11e1 	:	o_val <= 16'b0011011001100011;
            14'h11e2 	:	o_val <= 16'b0011011001100110;
            14'h11e3 	:	o_val <= 16'b0011011001101001;
            14'h11e4 	:	o_val <= 16'b0011011001101011;
            14'h11e5 	:	o_val <= 16'b0011011001101110;
            14'h11e6 	:	o_val <= 16'b0011011001110001;
            14'h11e7 	:	o_val <= 16'b0011011001110100;
            14'h11e8 	:	o_val <= 16'b0011011001110111;
            14'h11e9 	:	o_val <= 16'b0011011001111010;
            14'h11ea 	:	o_val <= 16'b0011011001111101;
            14'h11eb 	:	o_val <= 16'b0011011001111111;
            14'h11ec 	:	o_val <= 16'b0011011010000010;
            14'h11ed 	:	o_val <= 16'b0011011010000101;
            14'h11ee 	:	o_val <= 16'b0011011010001000;
            14'h11ef 	:	o_val <= 16'b0011011010001011;
            14'h11f0 	:	o_val <= 16'b0011011010001110;
            14'h11f1 	:	o_val <= 16'b0011011010010000;
            14'h11f2 	:	o_val <= 16'b0011011010010011;
            14'h11f3 	:	o_val <= 16'b0011011010010110;
            14'h11f4 	:	o_val <= 16'b0011011010011001;
            14'h11f5 	:	o_val <= 16'b0011011010011100;
            14'h11f6 	:	o_val <= 16'b0011011010011111;
            14'h11f7 	:	o_val <= 16'b0011011010100001;
            14'h11f8 	:	o_val <= 16'b0011011010100100;
            14'h11f9 	:	o_val <= 16'b0011011010100111;
            14'h11fa 	:	o_val <= 16'b0011011010101010;
            14'h11fb 	:	o_val <= 16'b0011011010101101;
            14'h11fc 	:	o_val <= 16'b0011011010110000;
            14'h11fd 	:	o_val <= 16'b0011011010110011;
            14'h11fe 	:	o_val <= 16'b0011011010110101;
            14'h11ff 	:	o_val <= 16'b0011011010111000;
            14'h1200 	:	o_val <= 16'b0011011010111011;
            14'h1201 	:	o_val <= 16'b0011011010111110;
            14'h1202 	:	o_val <= 16'b0011011011000001;
            14'h1203 	:	o_val <= 16'b0011011011000100;
            14'h1204 	:	o_val <= 16'b0011011011000110;
            14'h1205 	:	o_val <= 16'b0011011011001001;
            14'h1206 	:	o_val <= 16'b0011011011001100;
            14'h1207 	:	o_val <= 16'b0011011011001111;
            14'h1208 	:	o_val <= 16'b0011011011010010;
            14'h1209 	:	o_val <= 16'b0011011011010101;
            14'h120a 	:	o_val <= 16'b0011011011010111;
            14'h120b 	:	o_val <= 16'b0011011011011010;
            14'h120c 	:	o_val <= 16'b0011011011011101;
            14'h120d 	:	o_val <= 16'b0011011011100000;
            14'h120e 	:	o_val <= 16'b0011011011100011;
            14'h120f 	:	o_val <= 16'b0011011011100110;
            14'h1210 	:	o_val <= 16'b0011011011101000;
            14'h1211 	:	o_val <= 16'b0011011011101011;
            14'h1212 	:	o_val <= 16'b0011011011101110;
            14'h1213 	:	o_val <= 16'b0011011011110001;
            14'h1214 	:	o_val <= 16'b0011011011110100;
            14'h1215 	:	o_val <= 16'b0011011011110111;
            14'h1216 	:	o_val <= 16'b0011011011111001;
            14'h1217 	:	o_val <= 16'b0011011011111100;
            14'h1218 	:	o_val <= 16'b0011011011111111;
            14'h1219 	:	o_val <= 16'b0011011100000010;
            14'h121a 	:	o_val <= 16'b0011011100000101;
            14'h121b 	:	o_val <= 16'b0011011100001000;
            14'h121c 	:	o_val <= 16'b0011011100001011;
            14'h121d 	:	o_val <= 16'b0011011100001101;
            14'h121e 	:	o_val <= 16'b0011011100010000;
            14'h121f 	:	o_val <= 16'b0011011100010011;
            14'h1220 	:	o_val <= 16'b0011011100010110;
            14'h1221 	:	o_val <= 16'b0011011100011001;
            14'h1222 	:	o_val <= 16'b0011011100011100;
            14'h1223 	:	o_val <= 16'b0011011100011110;
            14'h1224 	:	o_val <= 16'b0011011100100001;
            14'h1225 	:	o_val <= 16'b0011011100100100;
            14'h1226 	:	o_val <= 16'b0011011100100111;
            14'h1227 	:	o_val <= 16'b0011011100101010;
            14'h1228 	:	o_val <= 16'b0011011100101101;
            14'h1229 	:	o_val <= 16'b0011011100101111;
            14'h122a 	:	o_val <= 16'b0011011100110010;
            14'h122b 	:	o_val <= 16'b0011011100110101;
            14'h122c 	:	o_val <= 16'b0011011100111000;
            14'h122d 	:	o_val <= 16'b0011011100111011;
            14'h122e 	:	o_val <= 16'b0011011100111110;
            14'h122f 	:	o_val <= 16'b0011011101000000;
            14'h1230 	:	o_val <= 16'b0011011101000011;
            14'h1231 	:	o_val <= 16'b0011011101000110;
            14'h1232 	:	o_val <= 16'b0011011101001001;
            14'h1233 	:	o_val <= 16'b0011011101001100;
            14'h1234 	:	o_val <= 16'b0011011101001111;
            14'h1235 	:	o_val <= 16'b0011011101010001;
            14'h1236 	:	o_val <= 16'b0011011101010100;
            14'h1237 	:	o_val <= 16'b0011011101010111;
            14'h1238 	:	o_val <= 16'b0011011101011010;
            14'h1239 	:	o_val <= 16'b0011011101011101;
            14'h123a 	:	o_val <= 16'b0011011101100000;
            14'h123b 	:	o_val <= 16'b0011011101100010;
            14'h123c 	:	o_val <= 16'b0011011101100101;
            14'h123d 	:	o_val <= 16'b0011011101101000;
            14'h123e 	:	o_val <= 16'b0011011101101011;
            14'h123f 	:	o_val <= 16'b0011011101101110;
            14'h1240 	:	o_val <= 16'b0011011101110001;
            14'h1241 	:	o_val <= 16'b0011011101110011;
            14'h1242 	:	o_val <= 16'b0011011101110110;
            14'h1243 	:	o_val <= 16'b0011011101111001;
            14'h1244 	:	o_val <= 16'b0011011101111100;
            14'h1245 	:	o_val <= 16'b0011011101111111;
            14'h1246 	:	o_val <= 16'b0011011110000010;
            14'h1247 	:	o_val <= 16'b0011011110000100;
            14'h1248 	:	o_val <= 16'b0011011110000111;
            14'h1249 	:	o_val <= 16'b0011011110001010;
            14'h124a 	:	o_val <= 16'b0011011110001101;
            14'h124b 	:	o_val <= 16'b0011011110010000;
            14'h124c 	:	o_val <= 16'b0011011110010011;
            14'h124d 	:	o_val <= 16'b0011011110010101;
            14'h124e 	:	o_val <= 16'b0011011110011000;
            14'h124f 	:	o_val <= 16'b0011011110011011;
            14'h1250 	:	o_val <= 16'b0011011110011110;
            14'h1251 	:	o_val <= 16'b0011011110100001;
            14'h1252 	:	o_val <= 16'b0011011110100011;
            14'h1253 	:	o_val <= 16'b0011011110100110;
            14'h1254 	:	o_val <= 16'b0011011110101001;
            14'h1255 	:	o_val <= 16'b0011011110101100;
            14'h1256 	:	o_val <= 16'b0011011110101111;
            14'h1257 	:	o_val <= 16'b0011011110110010;
            14'h1258 	:	o_val <= 16'b0011011110110100;
            14'h1259 	:	o_val <= 16'b0011011110110111;
            14'h125a 	:	o_val <= 16'b0011011110111010;
            14'h125b 	:	o_val <= 16'b0011011110111101;
            14'h125c 	:	o_val <= 16'b0011011111000000;
            14'h125d 	:	o_val <= 16'b0011011111000011;
            14'h125e 	:	o_val <= 16'b0011011111000101;
            14'h125f 	:	o_val <= 16'b0011011111001000;
            14'h1260 	:	o_val <= 16'b0011011111001011;
            14'h1261 	:	o_val <= 16'b0011011111001110;
            14'h1262 	:	o_val <= 16'b0011011111010001;
            14'h1263 	:	o_val <= 16'b0011011111010100;
            14'h1264 	:	o_val <= 16'b0011011111010110;
            14'h1265 	:	o_val <= 16'b0011011111011001;
            14'h1266 	:	o_val <= 16'b0011011111011100;
            14'h1267 	:	o_val <= 16'b0011011111011111;
            14'h1268 	:	o_val <= 16'b0011011111100010;
            14'h1269 	:	o_val <= 16'b0011011111100101;
            14'h126a 	:	o_val <= 16'b0011011111100111;
            14'h126b 	:	o_val <= 16'b0011011111101010;
            14'h126c 	:	o_val <= 16'b0011011111101101;
            14'h126d 	:	o_val <= 16'b0011011111110000;
            14'h126e 	:	o_val <= 16'b0011011111110011;
            14'h126f 	:	o_val <= 16'b0011011111110101;
            14'h1270 	:	o_val <= 16'b0011011111111000;
            14'h1271 	:	o_val <= 16'b0011011111111011;
            14'h1272 	:	o_val <= 16'b0011011111111110;
            14'h1273 	:	o_val <= 16'b0011100000000001;
            14'h1274 	:	o_val <= 16'b0011100000000100;
            14'h1275 	:	o_val <= 16'b0011100000000110;
            14'h1276 	:	o_val <= 16'b0011100000001001;
            14'h1277 	:	o_val <= 16'b0011100000001100;
            14'h1278 	:	o_val <= 16'b0011100000001111;
            14'h1279 	:	o_val <= 16'b0011100000010010;
            14'h127a 	:	o_val <= 16'b0011100000010101;
            14'h127b 	:	o_val <= 16'b0011100000010111;
            14'h127c 	:	o_val <= 16'b0011100000011010;
            14'h127d 	:	o_val <= 16'b0011100000011101;
            14'h127e 	:	o_val <= 16'b0011100000100000;
            14'h127f 	:	o_val <= 16'b0011100000100011;
            14'h1280 	:	o_val <= 16'b0011100000100101;
            14'h1281 	:	o_val <= 16'b0011100000101000;
            14'h1282 	:	o_val <= 16'b0011100000101011;
            14'h1283 	:	o_val <= 16'b0011100000101110;
            14'h1284 	:	o_val <= 16'b0011100000110001;
            14'h1285 	:	o_val <= 16'b0011100000110100;
            14'h1286 	:	o_val <= 16'b0011100000110110;
            14'h1287 	:	o_val <= 16'b0011100000111001;
            14'h1288 	:	o_val <= 16'b0011100000111100;
            14'h1289 	:	o_val <= 16'b0011100000111111;
            14'h128a 	:	o_val <= 16'b0011100001000010;
            14'h128b 	:	o_val <= 16'b0011100001000101;
            14'h128c 	:	o_val <= 16'b0011100001000111;
            14'h128d 	:	o_val <= 16'b0011100001001010;
            14'h128e 	:	o_val <= 16'b0011100001001101;
            14'h128f 	:	o_val <= 16'b0011100001010000;
            14'h1290 	:	o_val <= 16'b0011100001010011;
            14'h1291 	:	o_val <= 16'b0011100001010101;
            14'h1292 	:	o_val <= 16'b0011100001011000;
            14'h1293 	:	o_val <= 16'b0011100001011011;
            14'h1294 	:	o_val <= 16'b0011100001011110;
            14'h1295 	:	o_val <= 16'b0011100001100001;
            14'h1296 	:	o_val <= 16'b0011100001100100;
            14'h1297 	:	o_val <= 16'b0011100001100110;
            14'h1298 	:	o_val <= 16'b0011100001101001;
            14'h1299 	:	o_val <= 16'b0011100001101100;
            14'h129a 	:	o_val <= 16'b0011100001101111;
            14'h129b 	:	o_val <= 16'b0011100001110010;
            14'h129c 	:	o_val <= 16'b0011100001110100;
            14'h129d 	:	o_val <= 16'b0011100001110111;
            14'h129e 	:	o_val <= 16'b0011100001111010;
            14'h129f 	:	o_val <= 16'b0011100001111101;
            14'h12a0 	:	o_val <= 16'b0011100010000000;
            14'h12a1 	:	o_val <= 16'b0011100010000011;
            14'h12a2 	:	o_val <= 16'b0011100010000101;
            14'h12a3 	:	o_val <= 16'b0011100010001000;
            14'h12a4 	:	o_val <= 16'b0011100010001011;
            14'h12a5 	:	o_val <= 16'b0011100010001110;
            14'h12a6 	:	o_val <= 16'b0011100010010001;
            14'h12a7 	:	o_val <= 16'b0011100010010011;
            14'h12a8 	:	o_val <= 16'b0011100010010110;
            14'h12a9 	:	o_val <= 16'b0011100010011001;
            14'h12aa 	:	o_val <= 16'b0011100010011100;
            14'h12ab 	:	o_val <= 16'b0011100010011111;
            14'h12ac 	:	o_val <= 16'b0011100010100010;
            14'h12ad 	:	o_val <= 16'b0011100010100100;
            14'h12ae 	:	o_val <= 16'b0011100010100111;
            14'h12af 	:	o_val <= 16'b0011100010101010;
            14'h12b0 	:	o_val <= 16'b0011100010101101;
            14'h12b1 	:	o_val <= 16'b0011100010110000;
            14'h12b2 	:	o_val <= 16'b0011100010110010;
            14'h12b3 	:	o_val <= 16'b0011100010110101;
            14'h12b4 	:	o_val <= 16'b0011100010111000;
            14'h12b5 	:	o_val <= 16'b0011100010111011;
            14'h12b6 	:	o_val <= 16'b0011100010111110;
            14'h12b7 	:	o_val <= 16'b0011100011000001;
            14'h12b8 	:	o_val <= 16'b0011100011000011;
            14'h12b9 	:	o_val <= 16'b0011100011000110;
            14'h12ba 	:	o_val <= 16'b0011100011001001;
            14'h12bb 	:	o_val <= 16'b0011100011001100;
            14'h12bc 	:	o_val <= 16'b0011100011001111;
            14'h12bd 	:	o_val <= 16'b0011100011010001;
            14'h12be 	:	o_val <= 16'b0011100011010100;
            14'h12bf 	:	o_val <= 16'b0011100011010111;
            14'h12c0 	:	o_val <= 16'b0011100011011010;
            14'h12c1 	:	o_val <= 16'b0011100011011101;
            14'h12c2 	:	o_val <= 16'b0011100011100000;
            14'h12c3 	:	o_val <= 16'b0011100011100010;
            14'h12c4 	:	o_val <= 16'b0011100011100101;
            14'h12c5 	:	o_val <= 16'b0011100011101000;
            14'h12c6 	:	o_val <= 16'b0011100011101011;
            14'h12c7 	:	o_val <= 16'b0011100011101110;
            14'h12c8 	:	o_val <= 16'b0011100011110000;
            14'h12c9 	:	o_val <= 16'b0011100011110011;
            14'h12ca 	:	o_val <= 16'b0011100011110110;
            14'h12cb 	:	o_val <= 16'b0011100011111001;
            14'h12cc 	:	o_val <= 16'b0011100011111100;
            14'h12cd 	:	o_val <= 16'b0011100011111110;
            14'h12ce 	:	o_val <= 16'b0011100100000001;
            14'h12cf 	:	o_val <= 16'b0011100100000100;
            14'h12d0 	:	o_val <= 16'b0011100100000111;
            14'h12d1 	:	o_val <= 16'b0011100100001010;
            14'h12d2 	:	o_val <= 16'b0011100100001101;
            14'h12d3 	:	o_val <= 16'b0011100100001111;
            14'h12d4 	:	o_val <= 16'b0011100100010010;
            14'h12d5 	:	o_val <= 16'b0011100100010101;
            14'h12d6 	:	o_val <= 16'b0011100100011000;
            14'h12d7 	:	o_val <= 16'b0011100100011011;
            14'h12d8 	:	o_val <= 16'b0011100100011101;
            14'h12d9 	:	o_val <= 16'b0011100100100000;
            14'h12da 	:	o_val <= 16'b0011100100100011;
            14'h12db 	:	o_val <= 16'b0011100100100110;
            14'h12dc 	:	o_val <= 16'b0011100100101001;
            14'h12dd 	:	o_val <= 16'b0011100100101011;
            14'h12de 	:	o_val <= 16'b0011100100101110;
            14'h12df 	:	o_val <= 16'b0011100100110001;
            14'h12e0 	:	o_val <= 16'b0011100100110100;
            14'h12e1 	:	o_val <= 16'b0011100100110111;
            14'h12e2 	:	o_val <= 16'b0011100100111010;
            14'h12e3 	:	o_val <= 16'b0011100100111100;
            14'h12e4 	:	o_val <= 16'b0011100100111111;
            14'h12e5 	:	o_val <= 16'b0011100101000010;
            14'h12e6 	:	o_val <= 16'b0011100101000101;
            14'h12e7 	:	o_val <= 16'b0011100101001000;
            14'h12e8 	:	o_val <= 16'b0011100101001010;
            14'h12e9 	:	o_val <= 16'b0011100101001101;
            14'h12ea 	:	o_val <= 16'b0011100101010000;
            14'h12eb 	:	o_val <= 16'b0011100101010011;
            14'h12ec 	:	o_val <= 16'b0011100101010110;
            14'h12ed 	:	o_val <= 16'b0011100101011000;
            14'h12ee 	:	o_val <= 16'b0011100101011011;
            14'h12ef 	:	o_val <= 16'b0011100101011110;
            14'h12f0 	:	o_val <= 16'b0011100101100001;
            14'h12f1 	:	o_val <= 16'b0011100101100100;
            14'h12f2 	:	o_val <= 16'b0011100101100110;
            14'h12f3 	:	o_val <= 16'b0011100101101001;
            14'h12f4 	:	o_val <= 16'b0011100101101100;
            14'h12f5 	:	o_val <= 16'b0011100101101111;
            14'h12f6 	:	o_val <= 16'b0011100101110010;
            14'h12f7 	:	o_val <= 16'b0011100101110101;
            14'h12f8 	:	o_val <= 16'b0011100101110111;
            14'h12f9 	:	o_val <= 16'b0011100101111010;
            14'h12fa 	:	o_val <= 16'b0011100101111101;
            14'h12fb 	:	o_val <= 16'b0011100110000000;
            14'h12fc 	:	o_val <= 16'b0011100110000011;
            14'h12fd 	:	o_val <= 16'b0011100110000101;
            14'h12fe 	:	o_val <= 16'b0011100110001000;
            14'h12ff 	:	o_val <= 16'b0011100110001011;
            14'h1300 	:	o_val <= 16'b0011100110001110;
            14'h1301 	:	o_val <= 16'b0011100110010001;
            14'h1302 	:	o_val <= 16'b0011100110010011;
            14'h1303 	:	o_val <= 16'b0011100110010110;
            14'h1304 	:	o_val <= 16'b0011100110011001;
            14'h1305 	:	o_val <= 16'b0011100110011100;
            14'h1306 	:	o_val <= 16'b0011100110011111;
            14'h1307 	:	o_val <= 16'b0011100110100001;
            14'h1308 	:	o_val <= 16'b0011100110100100;
            14'h1309 	:	o_val <= 16'b0011100110100111;
            14'h130a 	:	o_val <= 16'b0011100110101010;
            14'h130b 	:	o_val <= 16'b0011100110101101;
            14'h130c 	:	o_val <= 16'b0011100110101111;
            14'h130d 	:	o_val <= 16'b0011100110110010;
            14'h130e 	:	o_val <= 16'b0011100110110101;
            14'h130f 	:	o_val <= 16'b0011100110111000;
            14'h1310 	:	o_val <= 16'b0011100110111011;
            14'h1311 	:	o_val <= 16'b0011100110111101;
            14'h1312 	:	o_val <= 16'b0011100111000000;
            14'h1313 	:	o_val <= 16'b0011100111000011;
            14'h1314 	:	o_val <= 16'b0011100111000110;
            14'h1315 	:	o_val <= 16'b0011100111001001;
            14'h1316 	:	o_val <= 16'b0011100111001011;
            14'h1317 	:	o_val <= 16'b0011100111001110;
            14'h1318 	:	o_val <= 16'b0011100111010001;
            14'h1319 	:	o_val <= 16'b0011100111010100;
            14'h131a 	:	o_val <= 16'b0011100111010111;
            14'h131b 	:	o_val <= 16'b0011100111011001;
            14'h131c 	:	o_val <= 16'b0011100111011100;
            14'h131d 	:	o_val <= 16'b0011100111011111;
            14'h131e 	:	o_val <= 16'b0011100111100010;
            14'h131f 	:	o_val <= 16'b0011100111100101;
            14'h1320 	:	o_val <= 16'b0011100111100111;
            14'h1321 	:	o_val <= 16'b0011100111101010;
            14'h1322 	:	o_val <= 16'b0011100111101101;
            14'h1323 	:	o_val <= 16'b0011100111110000;
            14'h1324 	:	o_val <= 16'b0011100111110011;
            14'h1325 	:	o_val <= 16'b0011100111110101;
            14'h1326 	:	o_val <= 16'b0011100111111000;
            14'h1327 	:	o_val <= 16'b0011100111111011;
            14'h1328 	:	o_val <= 16'b0011100111111110;
            14'h1329 	:	o_val <= 16'b0011101000000001;
            14'h132a 	:	o_val <= 16'b0011101000000100;
            14'h132b 	:	o_val <= 16'b0011101000000110;
            14'h132c 	:	o_val <= 16'b0011101000001001;
            14'h132d 	:	o_val <= 16'b0011101000001100;
            14'h132e 	:	o_val <= 16'b0011101000001111;
            14'h132f 	:	o_val <= 16'b0011101000010010;
            14'h1330 	:	o_val <= 16'b0011101000010100;
            14'h1331 	:	o_val <= 16'b0011101000010111;
            14'h1332 	:	o_val <= 16'b0011101000011010;
            14'h1333 	:	o_val <= 16'b0011101000011101;
            14'h1334 	:	o_val <= 16'b0011101000011111;
            14'h1335 	:	o_val <= 16'b0011101000100010;
            14'h1336 	:	o_val <= 16'b0011101000100101;
            14'h1337 	:	o_val <= 16'b0011101000101000;
            14'h1338 	:	o_val <= 16'b0011101000101011;
            14'h1339 	:	o_val <= 16'b0011101000101101;
            14'h133a 	:	o_val <= 16'b0011101000110000;
            14'h133b 	:	o_val <= 16'b0011101000110011;
            14'h133c 	:	o_val <= 16'b0011101000110110;
            14'h133d 	:	o_val <= 16'b0011101000111001;
            14'h133e 	:	o_val <= 16'b0011101000111011;
            14'h133f 	:	o_val <= 16'b0011101000111110;
            14'h1340 	:	o_val <= 16'b0011101001000001;
            14'h1341 	:	o_val <= 16'b0011101001000100;
            14'h1342 	:	o_val <= 16'b0011101001000111;
            14'h1343 	:	o_val <= 16'b0011101001001001;
            14'h1344 	:	o_val <= 16'b0011101001001100;
            14'h1345 	:	o_val <= 16'b0011101001001111;
            14'h1346 	:	o_val <= 16'b0011101001010010;
            14'h1347 	:	o_val <= 16'b0011101001010101;
            14'h1348 	:	o_val <= 16'b0011101001010111;
            14'h1349 	:	o_val <= 16'b0011101001011010;
            14'h134a 	:	o_val <= 16'b0011101001011101;
            14'h134b 	:	o_val <= 16'b0011101001100000;
            14'h134c 	:	o_val <= 16'b0011101001100011;
            14'h134d 	:	o_val <= 16'b0011101001100101;
            14'h134e 	:	o_val <= 16'b0011101001101000;
            14'h134f 	:	o_val <= 16'b0011101001101011;
            14'h1350 	:	o_val <= 16'b0011101001101110;
            14'h1351 	:	o_val <= 16'b0011101001110001;
            14'h1352 	:	o_val <= 16'b0011101001110011;
            14'h1353 	:	o_val <= 16'b0011101001110110;
            14'h1354 	:	o_val <= 16'b0011101001111001;
            14'h1355 	:	o_val <= 16'b0011101001111100;
            14'h1356 	:	o_val <= 16'b0011101001111111;
            14'h1357 	:	o_val <= 16'b0011101010000001;
            14'h1358 	:	o_val <= 16'b0011101010000100;
            14'h1359 	:	o_val <= 16'b0011101010000111;
            14'h135a 	:	o_val <= 16'b0011101010001010;
            14'h135b 	:	o_val <= 16'b0011101010001101;
            14'h135c 	:	o_val <= 16'b0011101010001111;
            14'h135d 	:	o_val <= 16'b0011101010010010;
            14'h135e 	:	o_val <= 16'b0011101010010101;
            14'h135f 	:	o_val <= 16'b0011101010011000;
            14'h1360 	:	o_val <= 16'b0011101010011011;
            14'h1361 	:	o_val <= 16'b0011101010011101;
            14'h1362 	:	o_val <= 16'b0011101010100000;
            14'h1363 	:	o_val <= 16'b0011101010100011;
            14'h1364 	:	o_val <= 16'b0011101010100110;
            14'h1365 	:	o_val <= 16'b0011101010101000;
            14'h1366 	:	o_val <= 16'b0011101010101011;
            14'h1367 	:	o_val <= 16'b0011101010101110;
            14'h1368 	:	o_val <= 16'b0011101010110001;
            14'h1369 	:	o_val <= 16'b0011101010110100;
            14'h136a 	:	o_val <= 16'b0011101010110110;
            14'h136b 	:	o_val <= 16'b0011101010111001;
            14'h136c 	:	o_val <= 16'b0011101010111100;
            14'h136d 	:	o_val <= 16'b0011101010111111;
            14'h136e 	:	o_val <= 16'b0011101011000010;
            14'h136f 	:	o_val <= 16'b0011101011000100;
            14'h1370 	:	o_val <= 16'b0011101011000111;
            14'h1371 	:	o_val <= 16'b0011101011001010;
            14'h1372 	:	o_val <= 16'b0011101011001101;
            14'h1373 	:	o_val <= 16'b0011101011010000;
            14'h1374 	:	o_val <= 16'b0011101011010010;
            14'h1375 	:	o_val <= 16'b0011101011010101;
            14'h1376 	:	o_val <= 16'b0011101011011000;
            14'h1377 	:	o_val <= 16'b0011101011011011;
            14'h1378 	:	o_val <= 16'b0011101011011110;
            14'h1379 	:	o_val <= 16'b0011101011100000;
            14'h137a 	:	o_val <= 16'b0011101011100011;
            14'h137b 	:	o_val <= 16'b0011101011100110;
            14'h137c 	:	o_val <= 16'b0011101011101001;
            14'h137d 	:	o_val <= 16'b0011101011101011;
            14'h137e 	:	o_val <= 16'b0011101011101110;
            14'h137f 	:	o_val <= 16'b0011101011110001;
            14'h1380 	:	o_val <= 16'b0011101011110100;
            14'h1381 	:	o_val <= 16'b0011101011110111;
            14'h1382 	:	o_val <= 16'b0011101011111001;
            14'h1383 	:	o_val <= 16'b0011101011111100;
            14'h1384 	:	o_val <= 16'b0011101011111111;
            14'h1385 	:	o_val <= 16'b0011101100000010;
            14'h1386 	:	o_val <= 16'b0011101100000101;
            14'h1387 	:	o_val <= 16'b0011101100000111;
            14'h1388 	:	o_val <= 16'b0011101100001010;
            14'h1389 	:	o_val <= 16'b0011101100001101;
            14'h138a 	:	o_val <= 16'b0011101100010000;
            14'h138b 	:	o_val <= 16'b0011101100010010;
            14'h138c 	:	o_val <= 16'b0011101100010101;
            14'h138d 	:	o_val <= 16'b0011101100011000;
            14'h138e 	:	o_val <= 16'b0011101100011011;
            14'h138f 	:	o_val <= 16'b0011101100011110;
            14'h1390 	:	o_val <= 16'b0011101100100000;
            14'h1391 	:	o_val <= 16'b0011101100100011;
            14'h1392 	:	o_val <= 16'b0011101100100110;
            14'h1393 	:	o_val <= 16'b0011101100101001;
            14'h1394 	:	o_val <= 16'b0011101100101100;
            14'h1395 	:	o_val <= 16'b0011101100101110;
            14'h1396 	:	o_val <= 16'b0011101100110001;
            14'h1397 	:	o_val <= 16'b0011101100110100;
            14'h1398 	:	o_val <= 16'b0011101100110111;
            14'h1399 	:	o_val <= 16'b0011101100111001;
            14'h139a 	:	o_val <= 16'b0011101100111100;
            14'h139b 	:	o_val <= 16'b0011101100111111;
            14'h139c 	:	o_val <= 16'b0011101101000010;
            14'h139d 	:	o_val <= 16'b0011101101000101;
            14'h139e 	:	o_val <= 16'b0011101101000111;
            14'h139f 	:	o_val <= 16'b0011101101001010;
            14'h13a0 	:	o_val <= 16'b0011101101001101;
            14'h13a1 	:	o_val <= 16'b0011101101010000;
            14'h13a2 	:	o_val <= 16'b0011101101010011;
            14'h13a3 	:	o_val <= 16'b0011101101010101;
            14'h13a4 	:	o_val <= 16'b0011101101011000;
            14'h13a5 	:	o_val <= 16'b0011101101011011;
            14'h13a6 	:	o_val <= 16'b0011101101011110;
            14'h13a7 	:	o_val <= 16'b0011101101100000;
            14'h13a8 	:	o_val <= 16'b0011101101100011;
            14'h13a9 	:	o_val <= 16'b0011101101100110;
            14'h13aa 	:	o_val <= 16'b0011101101101001;
            14'h13ab 	:	o_val <= 16'b0011101101101100;
            14'h13ac 	:	o_val <= 16'b0011101101101110;
            14'h13ad 	:	o_val <= 16'b0011101101110001;
            14'h13ae 	:	o_val <= 16'b0011101101110100;
            14'h13af 	:	o_val <= 16'b0011101101110111;
            14'h13b0 	:	o_val <= 16'b0011101101111010;
            14'h13b1 	:	o_val <= 16'b0011101101111100;
            14'h13b2 	:	o_val <= 16'b0011101101111111;
            14'h13b3 	:	o_val <= 16'b0011101110000010;
            14'h13b4 	:	o_val <= 16'b0011101110000101;
            14'h13b5 	:	o_val <= 16'b0011101110000111;
            14'h13b6 	:	o_val <= 16'b0011101110001010;
            14'h13b7 	:	o_val <= 16'b0011101110001101;
            14'h13b8 	:	o_val <= 16'b0011101110010000;
            14'h13b9 	:	o_val <= 16'b0011101110010011;
            14'h13ba 	:	o_val <= 16'b0011101110010101;
            14'h13bb 	:	o_val <= 16'b0011101110011000;
            14'h13bc 	:	o_val <= 16'b0011101110011011;
            14'h13bd 	:	o_val <= 16'b0011101110011110;
            14'h13be 	:	o_val <= 16'b0011101110100000;
            14'h13bf 	:	o_val <= 16'b0011101110100011;
            14'h13c0 	:	o_val <= 16'b0011101110100110;
            14'h13c1 	:	o_val <= 16'b0011101110101001;
            14'h13c2 	:	o_val <= 16'b0011101110101100;
            14'h13c3 	:	o_val <= 16'b0011101110101110;
            14'h13c4 	:	o_val <= 16'b0011101110110001;
            14'h13c5 	:	o_val <= 16'b0011101110110100;
            14'h13c6 	:	o_val <= 16'b0011101110110111;
            14'h13c7 	:	o_val <= 16'b0011101110111001;
            14'h13c8 	:	o_val <= 16'b0011101110111100;
            14'h13c9 	:	o_val <= 16'b0011101110111111;
            14'h13ca 	:	o_val <= 16'b0011101111000010;
            14'h13cb 	:	o_val <= 16'b0011101111000101;
            14'h13cc 	:	o_val <= 16'b0011101111000111;
            14'h13cd 	:	o_val <= 16'b0011101111001010;
            14'h13ce 	:	o_val <= 16'b0011101111001101;
            14'h13cf 	:	o_val <= 16'b0011101111010000;
            14'h13d0 	:	o_val <= 16'b0011101111010010;
            14'h13d1 	:	o_val <= 16'b0011101111010101;
            14'h13d2 	:	o_val <= 16'b0011101111011000;
            14'h13d3 	:	o_val <= 16'b0011101111011011;
            14'h13d4 	:	o_val <= 16'b0011101111011110;
            14'h13d5 	:	o_val <= 16'b0011101111100000;
            14'h13d6 	:	o_val <= 16'b0011101111100011;
            14'h13d7 	:	o_val <= 16'b0011101111100110;
            14'h13d8 	:	o_val <= 16'b0011101111101001;
            14'h13d9 	:	o_val <= 16'b0011101111101011;
            14'h13da 	:	o_val <= 16'b0011101111101110;
            14'h13db 	:	o_val <= 16'b0011101111110001;
            14'h13dc 	:	o_val <= 16'b0011101111110100;
            14'h13dd 	:	o_val <= 16'b0011101111110111;
            14'h13de 	:	o_val <= 16'b0011101111111001;
            14'h13df 	:	o_val <= 16'b0011101111111100;
            14'h13e0 	:	o_val <= 16'b0011101111111111;
            14'h13e1 	:	o_val <= 16'b0011110000000010;
            14'h13e2 	:	o_val <= 16'b0011110000000100;
            14'h13e3 	:	o_val <= 16'b0011110000000111;
            14'h13e4 	:	o_val <= 16'b0011110000001010;
            14'h13e5 	:	o_val <= 16'b0011110000001101;
            14'h13e6 	:	o_val <= 16'b0011110000010000;
            14'h13e7 	:	o_val <= 16'b0011110000010010;
            14'h13e8 	:	o_val <= 16'b0011110000010101;
            14'h13e9 	:	o_val <= 16'b0011110000011000;
            14'h13ea 	:	o_val <= 16'b0011110000011011;
            14'h13eb 	:	o_val <= 16'b0011110000011101;
            14'h13ec 	:	o_val <= 16'b0011110000100000;
            14'h13ed 	:	o_val <= 16'b0011110000100011;
            14'h13ee 	:	o_val <= 16'b0011110000100110;
            14'h13ef 	:	o_val <= 16'b0011110000101000;
            14'h13f0 	:	o_val <= 16'b0011110000101011;
            14'h13f1 	:	o_val <= 16'b0011110000101110;
            14'h13f2 	:	o_val <= 16'b0011110000110001;
            14'h13f3 	:	o_val <= 16'b0011110000110100;
            14'h13f4 	:	o_val <= 16'b0011110000110110;
            14'h13f5 	:	o_val <= 16'b0011110000111001;
            14'h13f6 	:	o_val <= 16'b0011110000111100;
            14'h13f7 	:	o_val <= 16'b0011110000111111;
            14'h13f8 	:	o_val <= 16'b0011110001000001;
            14'h13f9 	:	o_val <= 16'b0011110001000100;
            14'h13fa 	:	o_val <= 16'b0011110001000111;
            14'h13fb 	:	o_val <= 16'b0011110001001010;
            14'h13fc 	:	o_val <= 16'b0011110001001101;
            14'h13fd 	:	o_val <= 16'b0011110001001111;
            14'h13fe 	:	o_val <= 16'b0011110001010010;
            14'h13ff 	:	o_val <= 16'b0011110001010101;
            14'h1400 	:	o_val <= 16'b0011110001011000;
            14'h1401 	:	o_val <= 16'b0011110001011010;
            14'h1402 	:	o_val <= 16'b0011110001011101;
            14'h1403 	:	o_val <= 16'b0011110001100000;
            14'h1404 	:	o_val <= 16'b0011110001100011;
            14'h1405 	:	o_val <= 16'b0011110001100101;
            14'h1406 	:	o_val <= 16'b0011110001101000;
            14'h1407 	:	o_val <= 16'b0011110001101011;
            14'h1408 	:	o_val <= 16'b0011110001101110;
            14'h1409 	:	o_val <= 16'b0011110001110001;
            14'h140a 	:	o_val <= 16'b0011110001110011;
            14'h140b 	:	o_val <= 16'b0011110001110110;
            14'h140c 	:	o_val <= 16'b0011110001111001;
            14'h140d 	:	o_val <= 16'b0011110001111100;
            14'h140e 	:	o_val <= 16'b0011110001111110;
            14'h140f 	:	o_val <= 16'b0011110010000001;
            14'h1410 	:	o_val <= 16'b0011110010000100;
            14'h1411 	:	o_val <= 16'b0011110010000111;
            14'h1412 	:	o_val <= 16'b0011110010001001;
            14'h1413 	:	o_val <= 16'b0011110010001100;
            14'h1414 	:	o_val <= 16'b0011110010001111;
            14'h1415 	:	o_val <= 16'b0011110010010010;
            14'h1416 	:	o_val <= 16'b0011110010010101;
            14'h1417 	:	o_val <= 16'b0011110010010111;
            14'h1418 	:	o_val <= 16'b0011110010011010;
            14'h1419 	:	o_val <= 16'b0011110010011101;
            14'h141a 	:	o_val <= 16'b0011110010100000;
            14'h141b 	:	o_val <= 16'b0011110010100010;
            14'h141c 	:	o_val <= 16'b0011110010100101;
            14'h141d 	:	o_val <= 16'b0011110010101000;
            14'h141e 	:	o_val <= 16'b0011110010101011;
            14'h141f 	:	o_val <= 16'b0011110010101101;
            14'h1420 	:	o_val <= 16'b0011110010110000;
            14'h1421 	:	o_val <= 16'b0011110010110011;
            14'h1422 	:	o_val <= 16'b0011110010110110;
            14'h1423 	:	o_val <= 16'b0011110010111000;
            14'h1424 	:	o_val <= 16'b0011110010111011;
            14'h1425 	:	o_val <= 16'b0011110010111110;
            14'h1426 	:	o_val <= 16'b0011110011000001;
            14'h1427 	:	o_val <= 16'b0011110011000100;
            14'h1428 	:	o_val <= 16'b0011110011000110;
            14'h1429 	:	o_val <= 16'b0011110011001001;
            14'h142a 	:	o_val <= 16'b0011110011001100;
            14'h142b 	:	o_val <= 16'b0011110011001111;
            14'h142c 	:	o_val <= 16'b0011110011010001;
            14'h142d 	:	o_val <= 16'b0011110011010100;
            14'h142e 	:	o_val <= 16'b0011110011010111;
            14'h142f 	:	o_val <= 16'b0011110011011010;
            14'h1430 	:	o_val <= 16'b0011110011011100;
            14'h1431 	:	o_val <= 16'b0011110011011111;
            14'h1432 	:	o_val <= 16'b0011110011100010;
            14'h1433 	:	o_val <= 16'b0011110011100101;
            14'h1434 	:	o_val <= 16'b0011110011100111;
            14'h1435 	:	o_val <= 16'b0011110011101010;
            14'h1436 	:	o_val <= 16'b0011110011101101;
            14'h1437 	:	o_val <= 16'b0011110011110000;
            14'h1438 	:	o_val <= 16'b0011110011110011;
            14'h1439 	:	o_val <= 16'b0011110011110101;
            14'h143a 	:	o_val <= 16'b0011110011111000;
            14'h143b 	:	o_val <= 16'b0011110011111011;
            14'h143c 	:	o_val <= 16'b0011110011111110;
            14'h143d 	:	o_val <= 16'b0011110100000000;
            14'h143e 	:	o_val <= 16'b0011110100000011;
            14'h143f 	:	o_val <= 16'b0011110100000110;
            14'h1440 	:	o_val <= 16'b0011110100001001;
            14'h1441 	:	o_val <= 16'b0011110100001011;
            14'h1442 	:	o_val <= 16'b0011110100001110;
            14'h1443 	:	o_val <= 16'b0011110100010001;
            14'h1444 	:	o_val <= 16'b0011110100010100;
            14'h1445 	:	o_val <= 16'b0011110100010110;
            14'h1446 	:	o_val <= 16'b0011110100011001;
            14'h1447 	:	o_val <= 16'b0011110100011100;
            14'h1448 	:	o_val <= 16'b0011110100011111;
            14'h1449 	:	o_val <= 16'b0011110100100001;
            14'h144a 	:	o_val <= 16'b0011110100100100;
            14'h144b 	:	o_val <= 16'b0011110100100111;
            14'h144c 	:	o_val <= 16'b0011110100101010;
            14'h144d 	:	o_val <= 16'b0011110100101101;
            14'h144e 	:	o_val <= 16'b0011110100101111;
            14'h144f 	:	o_val <= 16'b0011110100110010;
            14'h1450 	:	o_val <= 16'b0011110100110101;
            14'h1451 	:	o_val <= 16'b0011110100111000;
            14'h1452 	:	o_val <= 16'b0011110100111010;
            14'h1453 	:	o_val <= 16'b0011110100111101;
            14'h1454 	:	o_val <= 16'b0011110101000000;
            14'h1455 	:	o_val <= 16'b0011110101000011;
            14'h1456 	:	o_val <= 16'b0011110101000101;
            14'h1457 	:	o_val <= 16'b0011110101001000;
            14'h1458 	:	o_val <= 16'b0011110101001011;
            14'h1459 	:	o_val <= 16'b0011110101001110;
            14'h145a 	:	o_val <= 16'b0011110101010000;
            14'h145b 	:	o_val <= 16'b0011110101010011;
            14'h145c 	:	o_val <= 16'b0011110101010110;
            14'h145d 	:	o_val <= 16'b0011110101011001;
            14'h145e 	:	o_val <= 16'b0011110101011011;
            14'h145f 	:	o_val <= 16'b0011110101011110;
            14'h1460 	:	o_val <= 16'b0011110101100001;
            14'h1461 	:	o_val <= 16'b0011110101100100;
            14'h1462 	:	o_val <= 16'b0011110101100110;
            14'h1463 	:	o_val <= 16'b0011110101101001;
            14'h1464 	:	o_val <= 16'b0011110101101100;
            14'h1465 	:	o_val <= 16'b0011110101101111;
            14'h1466 	:	o_val <= 16'b0011110101110001;
            14'h1467 	:	o_val <= 16'b0011110101110100;
            14'h1468 	:	o_val <= 16'b0011110101110111;
            14'h1469 	:	o_val <= 16'b0011110101111010;
            14'h146a 	:	o_val <= 16'b0011110101111100;
            14'h146b 	:	o_val <= 16'b0011110101111111;
            14'h146c 	:	o_val <= 16'b0011110110000010;
            14'h146d 	:	o_val <= 16'b0011110110000101;
            14'h146e 	:	o_val <= 16'b0011110110001000;
            14'h146f 	:	o_val <= 16'b0011110110001010;
            14'h1470 	:	o_val <= 16'b0011110110001101;
            14'h1471 	:	o_val <= 16'b0011110110010000;
            14'h1472 	:	o_val <= 16'b0011110110010011;
            14'h1473 	:	o_val <= 16'b0011110110010101;
            14'h1474 	:	o_val <= 16'b0011110110011000;
            14'h1475 	:	o_val <= 16'b0011110110011011;
            14'h1476 	:	o_val <= 16'b0011110110011110;
            14'h1477 	:	o_val <= 16'b0011110110100000;
            14'h1478 	:	o_val <= 16'b0011110110100011;
            14'h1479 	:	o_val <= 16'b0011110110100110;
            14'h147a 	:	o_val <= 16'b0011110110101001;
            14'h147b 	:	o_val <= 16'b0011110110101011;
            14'h147c 	:	o_val <= 16'b0011110110101110;
            14'h147d 	:	o_val <= 16'b0011110110110001;
            14'h147e 	:	o_val <= 16'b0011110110110100;
            14'h147f 	:	o_val <= 16'b0011110110110110;
            14'h1480 	:	o_val <= 16'b0011110110111001;
            14'h1481 	:	o_val <= 16'b0011110110111100;
            14'h1482 	:	o_val <= 16'b0011110110111111;
            14'h1483 	:	o_val <= 16'b0011110111000001;
            14'h1484 	:	o_val <= 16'b0011110111000100;
            14'h1485 	:	o_val <= 16'b0011110111000111;
            14'h1486 	:	o_val <= 16'b0011110111001010;
            14'h1487 	:	o_val <= 16'b0011110111001100;
            14'h1488 	:	o_val <= 16'b0011110111001111;
            14'h1489 	:	o_val <= 16'b0011110111010010;
            14'h148a 	:	o_val <= 16'b0011110111010101;
            14'h148b 	:	o_val <= 16'b0011110111010111;
            14'h148c 	:	o_val <= 16'b0011110111011010;
            14'h148d 	:	o_val <= 16'b0011110111011101;
            14'h148e 	:	o_val <= 16'b0011110111100000;
            14'h148f 	:	o_val <= 16'b0011110111100010;
            14'h1490 	:	o_val <= 16'b0011110111100101;
            14'h1491 	:	o_val <= 16'b0011110111101000;
            14'h1492 	:	o_val <= 16'b0011110111101011;
            14'h1493 	:	o_val <= 16'b0011110111101101;
            14'h1494 	:	o_val <= 16'b0011110111110000;
            14'h1495 	:	o_val <= 16'b0011110111110011;
            14'h1496 	:	o_val <= 16'b0011110111110110;
            14'h1497 	:	o_val <= 16'b0011110111111000;
            14'h1498 	:	o_val <= 16'b0011110111111011;
            14'h1499 	:	o_val <= 16'b0011110111111110;
            14'h149a 	:	o_val <= 16'b0011111000000001;
            14'h149b 	:	o_val <= 16'b0011111000000011;
            14'h149c 	:	o_val <= 16'b0011111000000110;
            14'h149d 	:	o_val <= 16'b0011111000001001;
            14'h149e 	:	o_val <= 16'b0011111000001100;
            14'h149f 	:	o_val <= 16'b0011111000001110;
            14'h14a0 	:	o_val <= 16'b0011111000010001;
            14'h14a1 	:	o_val <= 16'b0011111000010100;
            14'h14a2 	:	o_val <= 16'b0011111000010111;
            14'h14a3 	:	o_val <= 16'b0011111000011001;
            14'h14a4 	:	o_val <= 16'b0011111000011100;
            14'h14a5 	:	o_val <= 16'b0011111000011111;
            14'h14a6 	:	o_val <= 16'b0011111000100010;
            14'h14a7 	:	o_val <= 16'b0011111000100100;
            14'h14a8 	:	o_val <= 16'b0011111000100111;
            14'h14a9 	:	o_val <= 16'b0011111000101010;
            14'h14aa 	:	o_val <= 16'b0011111000101101;
            14'h14ab 	:	o_val <= 16'b0011111000101111;
            14'h14ac 	:	o_val <= 16'b0011111000110010;
            14'h14ad 	:	o_val <= 16'b0011111000110101;
            14'h14ae 	:	o_val <= 16'b0011111000111000;
            14'h14af 	:	o_val <= 16'b0011111000111010;
            14'h14b0 	:	o_val <= 16'b0011111000111101;
            14'h14b1 	:	o_val <= 16'b0011111001000000;
            14'h14b2 	:	o_val <= 16'b0011111001000011;
            14'h14b3 	:	o_val <= 16'b0011111001000101;
            14'h14b4 	:	o_val <= 16'b0011111001001000;
            14'h14b5 	:	o_val <= 16'b0011111001001011;
            14'h14b6 	:	o_val <= 16'b0011111001001101;
            14'h14b7 	:	o_val <= 16'b0011111001010000;
            14'h14b8 	:	o_val <= 16'b0011111001010011;
            14'h14b9 	:	o_val <= 16'b0011111001010110;
            14'h14ba 	:	o_val <= 16'b0011111001011000;
            14'h14bb 	:	o_val <= 16'b0011111001011011;
            14'h14bc 	:	o_val <= 16'b0011111001011110;
            14'h14bd 	:	o_val <= 16'b0011111001100001;
            14'h14be 	:	o_val <= 16'b0011111001100011;
            14'h14bf 	:	o_val <= 16'b0011111001100110;
            14'h14c0 	:	o_val <= 16'b0011111001101001;
            14'h14c1 	:	o_val <= 16'b0011111001101100;
            14'h14c2 	:	o_val <= 16'b0011111001101110;
            14'h14c3 	:	o_val <= 16'b0011111001110001;
            14'h14c4 	:	o_val <= 16'b0011111001110100;
            14'h14c5 	:	o_val <= 16'b0011111001110111;
            14'h14c6 	:	o_val <= 16'b0011111001111001;
            14'h14c7 	:	o_val <= 16'b0011111001111100;
            14'h14c8 	:	o_val <= 16'b0011111001111111;
            14'h14c9 	:	o_val <= 16'b0011111010000010;
            14'h14ca 	:	o_val <= 16'b0011111010000100;
            14'h14cb 	:	o_val <= 16'b0011111010000111;
            14'h14cc 	:	o_val <= 16'b0011111010001010;
            14'h14cd 	:	o_val <= 16'b0011111010001101;
            14'h14ce 	:	o_val <= 16'b0011111010001111;
            14'h14cf 	:	o_val <= 16'b0011111010010010;
            14'h14d0 	:	o_val <= 16'b0011111010010101;
            14'h14d1 	:	o_val <= 16'b0011111010011000;
            14'h14d2 	:	o_val <= 16'b0011111010011010;
            14'h14d3 	:	o_val <= 16'b0011111010011101;
            14'h14d4 	:	o_val <= 16'b0011111010100000;
            14'h14d5 	:	o_val <= 16'b0011111010100010;
            14'h14d6 	:	o_val <= 16'b0011111010100101;
            14'h14d7 	:	o_val <= 16'b0011111010101000;
            14'h14d8 	:	o_val <= 16'b0011111010101011;
            14'h14d9 	:	o_val <= 16'b0011111010101101;
            14'h14da 	:	o_val <= 16'b0011111010110000;
            14'h14db 	:	o_val <= 16'b0011111010110011;
            14'h14dc 	:	o_val <= 16'b0011111010110110;
            14'h14dd 	:	o_val <= 16'b0011111010111000;
            14'h14de 	:	o_val <= 16'b0011111010111011;
            14'h14df 	:	o_val <= 16'b0011111010111110;
            14'h14e0 	:	o_val <= 16'b0011111011000001;
            14'h14e1 	:	o_val <= 16'b0011111011000011;
            14'h14e2 	:	o_val <= 16'b0011111011000110;
            14'h14e3 	:	o_val <= 16'b0011111011001001;
            14'h14e4 	:	o_val <= 16'b0011111011001100;
            14'h14e5 	:	o_val <= 16'b0011111011001110;
            14'h14e6 	:	o_val <= 16'b0011111011010001;
            14'h14e7 	:	o_val <= 16'b0011111011010100;
            14'h14e8 	:	o_val <= 16'b0011111011010111;
            14'h14e9 	:	o_val <= 16'b0011111011011001;
            14'h14ea 	:	o_val <= 16'b0011111011011100;
            14'h14eb 	:	o_val <= 16'b0011111011011111;
            14'h14ec 	:	o_val <= 16'b0011111011100001;
            14'h14ed 	:	o_val <= 16'b0011111011100100;
            14'h14ee 	:	o_val <= 16'b0011111011100111;
            14'h14ef 	:	o_val <= 16'b0011111011101010;
            14'h14f0 	:	o_val <= 16'b0011111011101100;
            14'h14f1 	:	o_val <= 16'b0011111011101111;
            14'h14f2 	:	o_val <= 16'b0011111011110010;
            14'h14f3 	:	o_val <= 16'b0011111011110101;
            14'h14f4 	:	o_val <= 16'b0011111011110111;
            14'h14f5 	:	o_val <= 16'b0011111011111010;
            14'h14f6 	:	o_val <= 16'b0011111011111101;
            14'h14f7 	:	o_val <= 16'b0011111100000000;
            14'h14f8 	:	o_val <= 16'b0011111100000010;
            14'h14f9 	:	o_val <= 16'b0011111100000101;
            14'h14fa 	:	o_val <= 16'b0011111100001000;
            14'h14fb 	:	o_val <= 16'b0011111100001010;
            14'h14fc 	:	o_val <= 16'b0011111100001101;
            14'h14fd 	:	o_val <= 16'b0011111100010000;
            14'h14fe 	:	o_val <= 16'b0011111100010011;
            14'h14ff 	:	o_val <= 16'b0011111100010101;
            14'h1500 	:	o_val <= 16'b0011111100011000;
            14'h1501 	:	o_val <= 16'b0011111100011011;
            14'h1502 	:	o_val <= 16'b0011111100011110;
            14'h1503 	:	o_val <= 16'b0011111100100000;
            14'h1504 	:	o_val <= 16'b0011111100100011;
            14'h1505 	:	o_val <= 16'b0011111100100110;
            14'h1506 	:	o_val <= 16'b0011111100101001;
            14'h1507 	:	o_val <= 16'b0011111100101011;
            14'h1508 	:	o_val <= 16'b0011111100101110;
            14'h1509 	:	o_val <= 16'b0011111100110001;
            14'h150a 	:	o_val <= 16'b0011111100110011;
            14'h150b 	:	o_val <= 16'b0011111100110110;
            14'h150c 	:	o_val <= 16'b0011111100111001;
            14'h150d 	:	o_val <= 16'b0011111100111100;
            14'h150e 	:	o_val <= 16'b0011111100111110;
            14'h150f 	:	o_val <= 16'b0011111101000001;
            14'h1510 	:	o_val <= 16'b0011111101000100;
            14'h1511 	:	o_val <= 16'b0011111101000111;
            14'h1512 	:	o_val <= 16'b0011111101001001;
            14'h1513 	:	o_val <= 16'b0011111101001100;
            14'h1514 	:	o_val <= 16'b0011111101001111;
            14'h1515 	:	o_val <= 16'b0011111101010010;
            14'h1516 	:	o_val <= 16'b0011111101010100;
            14'h1517 	:	o_val <= 16'b0011111101010111;
            14'h1518 	:	o_val <= 16'b0011111101011010;
            14'h1519 	:	o_val <= 16'b0011111101011100;
            14'h151a 	:	o_val <= 16'b0011111101011111;
            14'h151b 	:	o_val <= 16'b0011111101100010;
            14'h151c 	:	o_val <= 16'b0011111101100101;
            14'h151d 	:	o_val <= 16'b0011111101100111;
            14'h151e 	:	o_val <= 16'b0011111101101010;
            14'h151f 	:	o_val <= 16'b0011111101101101;
            14'h1520 	:	o_val <= 16'b0011111101110000;
            14'h1521 	:	o_val <= 16'b0011111101110010;
            14'h1522 	:	o_val <= 16'b0011111101110101;
            14'h1523 	:	o_val <= 16'b0011111101111000;
            14'h1524 	:	o_val <= 16'b0011111101111010;
            14'h1525 	:	o_val <= 16'b0011111101111101;
            14'h1526 	:	o_val <= 16'b0011111110000000;
            14'h1527 	:	o_val <= 16'b0011111110000011;
            14'h1528 	:	o_val <= 16'b0011111110000101;
            14'h1529 	:	o_val <= 16'b0011111110001000;
            14'h152a 	:	o_val <= 16'b0011111110001011;
            14'h152b 	:	o_val <= 16'b0011111110001110;
            14'h152c 	:	o_val <= 16'b0011111110010000;
            14'h152d 	:	o_val <= 16'b0011111110010011;
            14'h152e 	:	o_val <= 16'b0011111110010110;
            14'h152f 	:	o_val <= 16'b0011111110011000;
            14'h1530 	:	o_val <= 16'b0011111110011011;
            14'h1531 	:	o_val <= 16'b0011111110011110;
            14'h1532 	:	o_val <= 16'b0011111110100001;
            14'h1533 	:	o_val <= 16'b0011111110100011;
            14'h1534 	:	o_val <= 16'b0011111110100110;
            14'h1535 	:	o_val <= 16'b0011111110101001;
            14'h1536 	:	o_val <= 16'b0011111110101100;
            14'h1537 	:	o_val <= 16'b0011111110101110;
            14'h1538 	:	o_val <= 16'b0011111110110001;
            14'h1539 	:	o_val <= 16'b0011111110110100;
            14'h153a 	:	o_val <= 16'b0011111110110110;
            14'h153b 	:	o_val <= 16'b0011111110111001;
            14'h153c 	:	o_val <= 16'b0011111110111100;
            14'h153d 	:	o_val <= 16'b0011111110111111;
            14'h153e 	:	o_val <= 16'b0011111111000001;
            14'h153f 	:	o_val <= 16'b0011111111000100;
            14'h1540 	:	o_val <= 16'b0011111111000111;
            14'h1541 	:	o_val <= 16'b0011111111001010;
            14'h1542 	:	o_val <= 16'b0011111111001100;
            14'h1543 	:	o_val <= 16'b0011111111001111;
            14'h1544 	:	o_val <= 16'b0011111111010010;
            14'h1545 	:	o_val <= 16'b0011111111010100;
            14'h1546 	:	o_val <= 16'b0011111111010111;
            14'h1547 	:	o_val <= 16'b0011111111011010;
            14'h1548 	:	o_val <= 16'b0011111111011101;
            14'h1549 	:	o_val <= 16'b0011111111011111;
            14'h154a 	:	o_val <= 16'b0011111111100010;
            14'h154b 	:	o_val <= 16'b0011111111100101;
            14'h154c 	:	o_val <= 16'b0011111111100111;
            14'h154d 	:	o_val <= 16'b0011111111101010;
            14'h154e 	:	o_val <= 16'b0011111111101101;
            14'h154f 	:	o_val <= 16'b0011111111110000;
            14'h1550 	:	o_val <= 16'b0011111111110010;
            14'h1551 	:	o_val <= 16'b0011111111110101;
            14'h1552 	:	o_val <= 16'b0011111111111000;
            14'h1553 	:	o_val <= 16'b0011111111111011;
            14'h1554 	:	o_val <= 16'b0011111111111101;
            14'h1555 	:	o_val <= 16'b0100000000000000;
            14'h1556 	:	o_val <= 16'b0100000000000011;
            14'h1557 	:	o_val <= 16'b0100000000000101;
            14'h1558 	:	o_val <= 16'b0100000000001000;
            14'h1559 	:	o_val <= 16'b0100000000001011;
            14'h155a 	:	o_val <= 16'b0100000000001110;
            14'h155b 	:	o_val <= 16'b0100000000010000;
            14'h155c 	:	o_val <= 16'b0100000000010011;
            14'h155d 	:	o_val <= 16'b0100000000010110;
            14'h155e 	:	o_val <= 16'b0100000000011000;
            14'h155f 	:	o_val <= 16'b0100000000011011;
            14'h1560 	:	o_val <= 16'b0100000000011110;
            14'h1561 	:	o_val <= 16'b0100000000100001;
            14'h1562 	:	o_val <= 16'b0100000000100011;
            14'h1563 	:	o_val <= 16'b0100000000100110;
            14'h1564 	:	o_val <= 16'b0100000000101001;
            14'h1565 	:	o_val <= 16'b0100000000101011;
            14'h1566 	:	o_val <= 16'b0100000000101110;
            14'h1567 	:	o_val <= 16'b0100000000110001;
            14'h1568 	:	o_val <= 16'b0100000000110100;
            14'h1569 	:	o_val <= 16'b0100000000110110;
            14'h156a 	:	o_val <= 16'b0100000000111001;
            14'h156b 	:	o_val <= 16'b0100000000111100;
            14'h156c 	:	o_val <= 16'b0100000000111110;
            14'h156d 	:	o_val <= 16'b0100000001000001;
            14'h156e 	:	o_val <= 16'b0100000001000100;
            14'h156f 	:	o_val <= 16'b0100000001000111;
            14'h1570 	:	o_val <= 16'b0100000001001001;
            14'h1571 	:	o_val <= 16'b0100000001001100;
            14'h1572 	:	o_val <= 16'b0100000001001111;
            14'h1573 	:	o_val <= 16'b0100000001010010;
            14'h1574 	:	o_val <= 16'b0100000001010100;
            14'h1575 	:	o_val <= 16'b0100000001010111;
            14'h1576 	:	o_val <= 16'b0100000001011010;
            14'h1577 	:	o_val <= 16'b0100000001011100;
            14'h1578 	:	o_val <= 16'b0100000001011111;
            14'h1579 	:	o_val <= 16'b0100000001100010;
            14'h157a 	:	o_val <= 16'b0100000001100101;
            14'h157b 	:	o_val <= 16'b0100000001100111;
            14'h157c 	:	o_val <= 16'b0100000001101010;
            14'h157d 	:	o_val <= 16'b0100000001101101;
            14'h157e 	:	o_val <= 16'b0100000001101111;
            14'h157f 	:	o_val <= 16'b0100000001110010;
            14'h1580 	:	o_val <= 16'b0100000001110101;
            14'h1581 	:	o_val <= 16'b0100000001111000;
            14'h1582 	:	o_val <= 16'b0100000001111010;
            14'h1583 	:	o_val <= 16'b0100000001111101;
            14'h1584 	:	o_val <= 16'b0100000010000000;
            14'h1585 	:	o_val <= 16'b0100000010000010;
            14'h1586 	:	o_val <= 16'b0100000010000101;
            14'h1587 	:	o_val <= 16'b0100000010001000;
            14'h1588 	:	o_val <= 16'b0100000010001011;
            14'h1589 	:	o_val <= 16'b0100000010001101;
            14'h158a 	:	o_val <= 16'b0100000010010000;
            14'h158b 	:	o_val <= 16'b0100000010010011;
            14'h158c 	:	o_val <= 16'b0100000010010101;
            14'h158d 	:	o_val <= 16'b0100000010011000;
            14'h158e 	:	o_val <= 16'b0100000010011011;
            14'h158f 	:	o_val <= 16'b0100000010011101;
            14'h1590 	:	o_val <= 16'b0100000010100000;
            14'h1591 	:	o_val <= 16'b0100000010100011;
            14'h1592 	:	o_val <= 16'b0100000010100110;
            14'h1593 	:	o_val <= 16'b0100000010101000;
            14'h1594 	:	o_val <= 16'b0100000010101011;
            14'h1595 	:	o_val <= 16'b0100000010101110;
            14'h1596 	:	o_val <= 16'b0100000010110000;
            14'h1597 	:	o_val <= 16'b0100000010110011;
            14'h1598 	:	o_val <= 16'b0100000010110110;
            14'h1599 	:	o_val <= 16'b0100000010111001;
            14'h159a 	:	o_val <= 16'b0100000010111011;
            14'h159b 	:	o_val <= 16'b0100000010111110;
            14'h159c 	:	o_val <= 16'b0100000011000001;
            14'h159d 	:	o_val <= 16'b0100000011000011;
            14'h159e 	:	o_val <= 16'b0100000011000110;
            14'h159f 	:	o_val <= 16'b0100000011001001;
            14'h15a0 	:	o_val <= 16'b0100000011001100;
            14'h15a1 	:	o_val <= 16'b0100000011001110;
            14'h15a2 	:	o_val <= 16'b0100000011010001;
            14'h15a3 	:	o_val <= 16'b0100000011010100;
            14'h15a4 	:	o_val <= 16'b0100000011010110;
            14'h15a5 	:	o_val <= 16'b0100000011011001;
            14'h15a6 	:	o_val <= 16'b0100000011011100;
            14'h15a7 	:	o_val <= 16'b0100000011011111;
            14'h15a8 	:	o_val <= 16'b0100000011100001;
            14'h15a9 	:	o_val <= 16'b0100000011100100;
            14'h15aa 	:	o_val <= 16'b0100000011100111;
            14'h15ab 	:	o_val <= 16'b0100000011101001;
            14'h15ac 	:	o_val <= 16'b0100000011101100;
            14'h15ad 	:	o_val <= 16'b0100000011101111;
            14'h15ae 	:	o_val <= 16'b0100000011110001;
            14'h15af 	:	o_val <= 16'b0100000011110100;
            14'h15b0 	:	o_val <= 16'b0100000011110111;
            14'h15b1 	:	o_val <= 16'b0100000011111010;
            14'h15b2 	:	o_val <= 16'b0100000011111100;
            14'h15b3 	:	o_val <= 16'b0100000011111111;
            14'h15b4 	:	o_val <= 16'b0100000100000010;
            14'h15b5 	:	o_val <= 16'b0100000100000100;
            14'h15b6 	:	o_val <= 16'b0100000100000111;
            14'h15b7 	:	o_val <= 16'b0100000100001010;
            14'h15b8 	:	o_val <= 16'b0100000100001101;
            14'h15b9 	:	o_val <= 16'b0100000100001111;
            14'h15ba 	:	o_val <= 16'b0100000100010010;
            14'h15bb 	:	o_val <= 16'b0100000100010101;
            14'h15bc 	:	o_val <= 16'b0100000100010111;
            14'h15bd 	:	o_val <= 16'b0100000100011010;
            14'h15be 	:	o_val <= 16'b0100000100011101;
            14'h15bf 	:	o_val <= 16'b0100000100011111;
            14'h15c0 	:	o_val <= 16'b0100000100100010;
            14'h15c1 	:	o_val <= 16'b0100000100100101;
            14'h15c2 	:	o_val <= 16'b0100000100101000;
            14'h15c3 	:	o_val <= 16'b0100000100101010;
            14'h15c4 	:	o_val <= 16'b0100000100101101;
            14'h15c5 	:	o_val <= 16'b0100000100110000;
            14'h15c6 	:	o_val <= 16'b0100000100110010;
            14'h15c7 	:	o_val <= 16'b0100000100110101;
            14'h15c8 	:	o_val <= 16'b0100000100111000;
            14'h15c9 	:	o_val <= 16'b0100000100111011;
            14'h15ca 	:	o_val <= 16'b0100000100111101;
            14'h15cb 	:	o_val <= 16'b0100000101000000;
            14'h15cc 	:	o_val <= 16'b0100000101000011;
            14'h15cd 	:	o_val <= 16'b0100000101000101;
            14'h15ce 	:	o_val <= 16'b0100000101001000;
            14'h15cf 	:	o_val <= 16'b0100000101001011;
            14'h15d0 	:	o_val <= 16'b0100000101001101;
            14'h15d1 	:	o_val <= 16'b0100000101010000;
            14'h15d2 	:	o_val <= 16'b0100000101010011;
            14'h15d3 	:	o_val <= 16'b0100000101010110;
            14'h15d4 	:	o_val <= 16'b0100000101011000;
            14'h15d5 	:	o_val <= 16'b0100000101011011;
            14'h15d6 	:	o_val <= 16'b0100000101011110;
            14'h15d7 	:	o_val <= 16'b0100000101100000;
            14'h15d8 	:	o_val <= 16'b0100000101100011;
            14'h15d9 	:	o_val <= 16'b0100000101100110;
            14'h15da 	:	o_val <= 16'b0100000101101000;
            14'h15db 	:	o_val <= 16'b0100000101101011;
            14'h15dc 	:	o_val <= 16'b0100000101101110;
            14'h15dd 	:	o_val <= 16'b0100000101110001;
            14'h15de 	:	o_val <= 16'b0100000101110011;
            14'h15df 	:	o_val <= 16'b0100000101110110;
            14'h15e0 	:	o_val <= 16'b0100000101111001;
            14'h15e1 	:	o_val <= 16'b0100000101111011;
            14'h15e2 	:	o_val <= 16'b0100000101111110;
            14'h15e3 	:	o_val <= 16'b0100000110000001;
            14'h15e4 	:	o_val <= 16'b0100000110000011;
            14'h15e5 	:	o_val <= 16'b0100000110000110;
            14'h15e6 	:	o_val <= 16'b0100000110001001;
            14'h15e7 	:	o_val <= 16'b0100000110001100;
            14'h15e8 	:	o_val <= 16'b0100000110001110;
            14'h15e9 	:	o_val <= 16'b0100000110010001;
            14'h15ea 	:	o_val <= 16'b0100000110010100;
            14'h15eb 	:	o_val <= 16'b0100000110010110;
            14'h15ec 	:	o_val <= 16'b0100000110011001;
            14'h15ed 	:	o_val <= 16'b0100000110011100;
            14'h15ee 	:	o_val <= 16'b0100000110011110;
            14'h15ef 	:	o_val <= 16'b0100000110100001;
            14'h15f0 	:	o_val <= 16'b0100000110100100;
            14'h15f1 	:	o_val <= 16'b0100000110100111;
            14'h15f2 	:	o_val <= 16'b0100000110101001;
            14'h15f3 	:	o_val <= 16'b0100000110101100;
            14'h15f4 	:	o_val <= 16'b0100000110101111;
            14'h15f5 	:	o_val <= 16'b0100000110110001;
            14'h15f6 	:	o_val <= 16'b0100000110110100;
            14'h15f7 	:	o_val <= 16'b0100000110110111;
            14'h15f8 	:	o_val <= 16'b0100000110111001;
            14'h15f9 	:	o_val <= 16'b0100000110111100;
            14'h15fa 	:	o_val <= 16'b0100000110111111;
            14'h15fb 	:	o_val <= 16'b0100000111000001;
            14'h15fc 	:	o_val <= 16'b0100000111000100;
            14'h15fd 	:	o_val <= 16'b0100000111000111;
            14'h15fe 	:	o_val <= 16'b0100000111001010;
            14'h15ff 	:	o_val <= 16'b0100000111001100;
            14'h1600 	:	o_val <= 16'b0100000111001111;
            14'h1601 	:	o_val <= 16'b0100000111010010;
            14'h1602 	:	o_val <= 16'b0100000111010100;
            14'h1603 	:	o_val <= 16'b0100000111010111;
            14'h1604 	:	o_val <= 16'b0100000111011010;
            14'h1605 	:	o_val <= 16'b0100000111011100;
            14'h1606 	:	o_val <= 16'b0100000111011111;
            14'h1607 	:	o_val <= 16'b0100000111100010;
            14'h1608 	:	o_val <= 16'b0100000111100101;
            14'h1609 	:	o_val <= 16'b0100000111100111;
            14'h160a 	:	o_val <= 16'b0100000111101010;
            14'h160b 	:	o_val <= 16'b0100000111101101;
            14'h160c 	:	o_val <= 16'b0100000111101111;
            14'h160d 	:	o_val <= 16'b0100000111110010;
            14'h160e 	:	o_val <= 16'b0100000111110101;
            14'h160f 	:	o_val <= 16'b0100000111110111;
            14'h1610 	:	o_val <= 16'b0100000111111010;
            14'h1611 	:	o_val <= 16'b0100000111111101;
            14'h1612 	:	o_val <= 16'b0100000111111111;
            14'h1613 	:	o_val <= 16'b0100001000000010;
            14'h1614 	:	o_val <= 16'b0100001000000101;
            14'h1615 	:	o_val <= 16'b0100001000001000;
            14'h1616 	:	o_val <= 16'b0100001000001010;
            14'h1617 	:	o_val <= 16'b0100001000001101;
            14'h1618 	:	o_val <= 16'b0100001000010000;
            14'h1619 	:	o_val <= 16'b0100001000010010;
            14'h161a 	:	o_val <= 16'b0100001000010101;
            14'h161b 	:	o_val <= 16'b0100001000011000;
            14'h161c 	:	o_val <= 16'b0100001000011010;
            14'h161d 	:	o_val <= 16'b0100001000011101;
            14'h161e 	:	o_val <= 16'b0100001000100000;
            14'h161f 	:	o_val <= 16'b0100001000100010;
            14'h1620 	:	o_val <= 16'b0100001000100101;
            14'h1621 	:	o_val <= 16'b0100001000101000;
            14'h1622 	:	o_val <= 16'b0100001000101010;
            14'h1623 	:	o_val <= 16'b0100001000101101;
            14'h1624 	:	o_val <= 16'b0100001000110000;
            14'h1625 	:	o_val <= 16'b0100001000110011;
            14'h1626 	:	o_val <= 16'b0100001000110101;
            14'h1627 	:	o_val <= 16'b0100001000111000;
            14'h1628 	:	o_val <= 16'b0100001000111011;
            14'h1629 	:	o_val <= 16'b0100001000111101;
            14'h162a 	:	o_val <= 16'b0100001001000000;
            14'h162b 	:	o_val <= 16'b0100001001000011;
            14'h162c 	:	o_val <= 16'b0100001001000101;
            14'h162d 	:	o_val <= 16'b0100001001001000;
            14'h162e 	:	o_val <= 16'b0100001001001011;
            14'h162f 	:	o_val <= 16'b0100001001001101;
            14'h1630 	:	o_val <= 16'b0100001001010000;
            14'h1631 	:	o_val <= 16'b0100001001010011;
            14'h1632 	:	o_val <= 16'b0100001001010101;
            14'h1633 	:	o_val <= 16'b0100001001011000;
            14'h1634 	:	o_val <= 16'b0100001001011011;
            14'h1635 	:	o_val <= 16'b0100001001011110;
            14'h1636 	:	o_val <= 16'b0100001001100000;
            14'h1637 	:	o_val <= 16'b0100001001100011;
            14'h1638 	:	o_val <= 16'b0100001001100110;
            14'h1639 	:	o_val <= 16'b0100001001101000;
            14'h163a 	:	o_val <= 16'b0100001001101011;
            14'h163b 	:	o_val <= 16'b0100001001101110;
            14'h163c 	:	o_val <= 16'b0100001001110000;
            14'h163d 	:	o_val <= 16'b0100001001110011;
            14'h163e 	:	o_val <= 16'b0100001001110110;
            14'h163f 	:	o_val <= 16'b0100001001111000;
            14'h1640 	:	o_val <= 16'b0100001001111011;
            14'h1641 	:	o_val <= 16'b0100001001111110;
            14'h1642 	:	o_val <= 16'b0100001010000000;
            14'h1643 	:	o_val <= 16'b0100001010000011;
            14'h1644 	:	o_val <= 16'b0100001010000110;
            14'h1645 	:	o_val <= 16'b0100001010001001;
            14'h1646 	:	o_val <= 16'b0100001010001011;
            14'h1647 	:	o_val <= 16'b0100001010001110;
            14'h1648 	:	o_val <= 16'b0100001010010001;
            14'h1649 	:	o_val <= 16'b0100001010010011;
            14'h164a 	:	o_val <= 16'b0100001010010110;
            14'h164b 	:	o_val <= 16'b0100001010011001;
            14'h164c 	:	o_val <= 16'b0100001010011011;
            14'h164d 	:	o_val <= 16'b0100001010011110;
            14'h164e 	:	o_val <= 16'b0100001010100001;
            14'h164f 	:	o_val <= 16'b0100001010100011;
            14'h1650 	:	o_val <= 16'b0100001010100110;
            14'h1651 	:	o_val <= 16'b0100001010101001;
            14'h1652 	:	o_val <= 16'b0100001010101011;
            14'h1653 	:	o_val <= 16'b0100001010101110;
            14'h1654 	:	o_val <= 16'b0100001010110001;
            14'h1655 	:	o_val <= 16'b0100001010110011;
            14'h1656 	:	o_val <= 16'b0100001010110110;
            14'h1657 	:	o_val <= 16'b0100001010111001;
            14'h1658 	:	o_val <= 16'b0100001010111011;
            14'h1659 	:	o_val <= 16'b0100001010111110;
            14'h165a 	:	o_val <= 16'b0100001011000001;
            14'h165b 	:	o_val <= 16'b0100001011000100;
            14'h165c 	:	o_val <= 16'b0100001011000110;
            14'h165d 	:	o_val <= 16'b0100001011001001;
            14'h165e 	:	o_val <= 16'b0100001011001100;
            14'h165f 	:	o_val <= 16'b0100001011001110;
            14'h1660 	:	o_val <= 16'b0100001011010001;
            14'h1661 	:	o_val <= 16'b0100001011010100;
            14'h1662 	:	o_val <= 16'b0100001011010110;
            14'h1663 	:	o_val <= 16'b0100001011011001;
            14'h1664 	:	o_val <= 16'b0100001011011100;
            14'h1665 	:	o_val <= 16'b0100001011011110;
            14'h1666 	:	o_val <= 16'b0100001011100001;
            14'h1667 	:	o_val <= 16'b0100001011100100;
            14'h1668 	:	o_val <= 16'b0100001011100110;
            14'h1669 	:	o_val <= 16'b0100001011101001;
            14'h166a 	:	o_val <= 16'b0100001011101100;
            14'h166b 	:	o_val <= 16'b0100001011101110;
            14'h166c 	:	o_val <= 16'b0100001011110001;
            14'h166d 	:	o_val <= 16'b0100001011110100;
            14'h166e 	:	o_val <= 16'b0100001011110110;
            14'h166f 	:	o_val <= 16'b0100001011111001;
            14'h1670 	:	o_val <= 16'b0100001011111100;
            14'h1671 	:	o_val <= 16'b0100001011111110;
            14'h1672 	:	o_val <= 16'b0100001100000001;
            14'h1673 	:	o_val <= 16'b0100001100000100;
            14'h1674 	:	o_val <= 16'b0100001100000110;
            14'h1675 	:	o_val <= 16'b0100001100001001;
            14'h1676 	:	o_val <= 16'b0100001100001100;
            14'h1677 	:	o_val <= 16'b0100001100001111;
            14'h1678 	:	o_val <= 16'b0100001100010001;
            14'h1679 	:	o_val <= 16'b0100001100010100;
            14'h167a 	:	o_val <= 16'b0100001100010111;
            14'h167b 	:	o_val <= 16'b0100001100011001;
            14'h167c 	:	o_val <= 16'b0100001100011100;
            14'h167d 	:	o_val <= 16'b0100001100011111;
            14'h167e 	:	o_val <= 16'b0100001100100001;
            14'h167f 	:	o_val <= 16'b0100001100100100;
            14'h1680 	:	o_val <= 16'b0100001100100111;
            14'h1681 	:	o_val <= 16'b0100001100101001;
            14'h1682 	:	o_val <= 16'b0100001100101100;
            14'h1683 	:	o_val <= 16'b0100001100101111;
            14'h1684 	:	o_val <= 16'b0100001100110001;
            14'h1685 	:	o_val <= 16'b0100001100110100;
            14'h1686 	:	o_val <= 16'b0100001100110111;
            14'h1687 	:	o_val <= 16'b0100001100111001;
            14'h1688 	:	o_val <= 16'b0100001100111100;
            14'h1689 	:	o_val <= 16'b0100001100111111;
            14'h168a 	:	o_val <= 16'b0100001101000001;
            14'h168b 	:	o_val <= 16'b0100001101000100;
            14'h168c 	:	o_val <= 16'b0100001101000111;
            14'h168d 	:	o_val <= 16'b0100001101001001;
            14'h168e 	:	o_val <= 16'b0100001101001100;
            14'h168f 	:	o_val <= 16'b0100001101001111;
            14'h1690 	:	o_val <= 16'b0100001101010001;
            14'h1691 	:	o_val <= 16'b0100001101010100;
            14'h1692 	:	o_val <= 16'b0100001101010111;
            14'h1693 	:	o_val <= 16'b0100001101011001;
            14'h1694 	:	o_val <= 16'b0100001101011100;
            14'h1695 	:	o_val <= 16'b0100001101011111;
            14'h1696 	:	o_val <= 16'b0100001101100001;
            14'h1697 	:	o_val <= 16'b0100001101100100;
            14'h1698 	:	o_val <= 16'b0100001101100111;
            14'h1699 	:	o_val <= 16'b0100001101101001;
            14'h169a 	:	o_val <= 16'b0100001101101100;
            14'h169b 	:	o_val <= 16'b0100001101101111;
            14'h169c 	:	o_val <= 16'b0100001101110001;
            14'h169d 	:	o_val <= 16'b0100001101110100;
            14'h169e 	:	o_val <= 16'b0100001101110111;
            14'h169f 	:	o_val <= 16'b0100001101111001;
            14'h16a0 	:	o_val <= 16'b0100001101111100;
            14'h16a1 	:	o_val <= 16'b0100001101111111;
            14'h16a2 	:	o_val <= 16'b0100001110000001;
            14'h16a3 	:	o_val <= 16'b0100001110000100;
            14'h16a4 	:	o_val <= 16'b0100001110000111;
            14'h16a5 	:	o_val <= 16'b0100001110001001;
            14'h16a6 	:	o_val <= 16'b0100001110001100;
            14'h16a7 	:	o_val <= 16'b0100001110001111;
            14'h16a8 	:	o_val <= 16'b0100001110010001;
            14'h16a9 	:	o_val <= 16'b0100001110010100;
            14'h16aa 	:	o_val <= 16'b0100001110010111;
            14'h16ab 	:	o_val <= 16'b0100001110011001;
            14'h16ac 	:	o_val <= 16'b0100001110011100;
            14'h16ad 	:	o_val <= 16'b0100001110011111;
            14'h16ae 	:	o_val <= 16'b0100001110100001;
            14'h16af 	:	o_val <= 16'b0100001110100100;
            14'h16b0 	:	o_val <= 16'b0100001110100111;
            14'h16b1 	:	o_val <= 16'b0100001110101001;
            14'h16b2 	:	o_val <= 16'b0100001110101100;
            14'h16b3 	:	o_val <= 16'b0100001110101111;
            14'h16b4 	:	o_val <= 16'b0100001110110001;
            14'h16b5 	:	o_val <= 16'b0100001110110100;
            14'h16b6 	:	o_val <= 16'b0100001110110111;
            14'h16b7 	:	o_val <= 16'b0100001110111001;
            14'h16b8 	:	o_val <= 16'b0100001110111100;
            14'h16b9 	:	o_val <= 16'b0100001110111111;
            14'h16ba 	:	o_val <= 16'b0100001111000001;
            14'h16bb 	:	o_val <= 16'b0100001111000100;
            14'h16bc 	:	o_val <= 16'b0100001111000111;
            14'h16bd 	:	o_val <= 16'b0100001111001001;
            14'h16be 	:	o_val <= 16'b0100001111001100;
            14'h16bf 	:	o_val <= 16'b0100001111001111;
            14'h16c0 	:	o_val <= 16'b0100001111010001;
            14'h16c1 	:	o_val <= 16'b0100001111010100;
            14'h16c2 	:	o_val <= 16'b0100001111010111;
            14'h16c3 	:	o_val <= 16'b0100001111011001;
            14'h16c4 	:	o_val <= 16'b0100001111011100;
            14'h16c5 	:	o_val <= 16'b0100001111011111;
            14'h16c6 	:	o_val <= 16'b0100001111100001;
            14'h16c7 	:	o_val <= 16'b0100001111100100;
            14'h16c8 	:	o_val <= 16'b0100001111100111;
            14'h16c9 	:	o_val <= 16'b0100001111101001;
            14'h16ca 	:	o_val <= 16'b0100001111101100;
            14'h16cb 	:	o_val <= 16'b0100001111101111;
            14'h16cc 	:	o_val <= 16'b0100001111110001;
            14'h16cd 	:	o_val <= 16'b0100001111110100;
            14'h16ce 	:	o_val <= 16'b0100001111110111;
            14'h16cf 	:	o_val <= 16'b0100001111111001;
            14'h16d0 	:	o_val <= 16'b0100001111111100;
            14'h16d1 	:	o_val <= 16'b0100001111111111;
            14'h16d2 	:	o_val <= 16'b0100010000000001;
            14'h16d3 	:	o_val <= 16'b0100010000000100;
            14'h16d4 	:	o_val <= 16'b0100010000000111;
            14'h16d5 	:	o_val <= 16'b0100010000001001;
            14'h16d6 	:	o_val <= 16'b0100010000001100;
            14'h16d7 	:	o_val <= 16'b0100010000001111;
            14'h16d8 	:	o_val <= 16'b0100010000010001;
            14'h16d9 	:	o_val <= 16'b0100010000010100;
            14'h16da 	:	o_val <= 16'b0100010000010111;
            14'h16db 	:	o_val <= 16'b0100010000011001;
            14'h16dc 	:	o_val <= 16'b0100010000011100;
            14'h16dd 	:	o_val <= 16'b0100010000011111;
            14'h16de 	:	o_val <= 16'b0100010000100001;
            14'h16df 	:	o_val <= 16'b0100010000100100;
            14'h16e0 	:	o_val <= 16'b0100010000100111;
            14'h16e1 	:	o_val <= 16'b0100010000101001;
            14'h16e2 	:	o_val <= 16'b0100010000101100;
            14'h16e3 	:	o_val <= 16'b0100010000101111;
            14'h16e4 	:	o_val <= 16'b0100010000110001;
            14'h16e5 	:	o_val <= 16'b0100010000110100;
            14'h16e6 	:	o_val <= 16'b0100010000110111;
            14'h16e7 	:	o_val <= 16'b0100010000111001;
            14'h16e8 	:	o_val <= 16'b0100010000111100;
            14'h16e9 	:	o_val <= 16'b0100010000111111;
            14'h16ea 	:	o_val <= 16'b0100010001000001;
            14'h16eb 	:	o_val <= 16'b0100010001000100;
            14'h16ec 	:	o_val <= 16'b0100010001000111;
            14'h16ed 	:	o_val <= 16'b0100010001001001;
            14'h16ee 	:	o_val <= 16'b0100010001001100;
            14'h16ef 	:	o_val <= 16'b0100010001001110;
            14'h16f0 	:	o_val <= 16'b0100010001010001;
            14'h16f1 	:	o_val <= 16'b0100010001010100;
            14'h16f2 	:	o_val <= 16'b0100010001010110;
            14'h16f3 	:	o_val <= 16'b0100010001011001;
            14'h16f4 	:	o_val <= 16'b0100010001011100;
            14'h16f5 	:	o_val <= 16'b0100010001011110;
            14'h16f6 	:	o_val <= 16'b0100010001100001;
            14'h16f7 	:	o_val <= 16'b0100010001100100;
            14'h16f8 	:	o_val <= 16'b0100010001100110;
            14'h16f9 	:	o_val <= 16'b0100010001101001;
            14'h16fa 	:	o_val <= 16'b0100010001101100;
            14'h16fb 	:	o_val <= 16'b0100010001101110;
            14'h16fc 	:	o_val <= 16'b0100010001110001;
            14'h16fd 	:	o_val <= 16'b0100010001110100;
            14'h16fe 	:	o_val <= 16'b0100010001110110;
            14'h16ff 	:	o_val <= 16'b0100010001111001;
            14'h1700 	:	o_val <= 16'b0100010001111100;
            14'h1701 	:	o_val <= 16'b0100010001111110;
            14'h1702 	:	o_val <= 16'b0100010010000001;
            14'h1703 	:	o_val <= 16'b0100010010000100;
            14'h1704 	:	o_val <= 16'b0100010010000110;
            14'h1705 	:	o_val <= 16'b0100010010001001;
            14'h1706 	:	o_val <= 16'b0100010010001100;
            14'h1707 	:	o_val <= 16'b0100010010001110;
            14'h1708 	:	o_val <= 16'b0100010010010001;
            14'h1709 	:	o_val <= 16'b0100010010010100;
            14'h170a 	:	o_val <= 16'b0100010010010110;
            14'h170b 	:	o_val <= 16'b0100010010011001;
            14'h170c 	:	o_val <= 16'b0100010010011011;
            14'h170d 	:	o_val <= 16'b0100010010011110;
            14'h170e 	:	o_val <= 16'b0100010010100001;
            14'h170f 	:	o_val <= 16'b0100010010100011;
            14'h1710 	:	o_val <= 16'b0100010010100110;
            14'h1711 	:	o_val <= 16'b0100010010101001;
            14'h1712 	:	o_val <= 16'b0100010010101011;
            14'h1713 	:	o_val <= 16'b0100010010101110;
            14'h1714 	:	o_val <= 16'b0100010010110001;
            14'h1715 	:	o_val <= 16'b0100010010110011;
            14'h1716 	:	o_val <= 16'b0100010010110110;
            14'h1717 	:	o_val <= 16'b0100010010111001;
            14'h1718 	:	o_val <= 16'b0100010010111011;
            14'h1719 	:	o_val <= 16'b0100010010111110;
            14'h171a 	:	o_val <= 16'b0100010011000001;
            14'h171b 	:	o_val <= 16'b0100010011000011;
            14'h171c 	:	o_val <= 16'b0100010011000110;
            14'h171d 	:	o_val <= 16'b0100010011001001;
            14'h171e 	:	o_val <= 16'b0100010011001011;
            14'h171f 	:	o_val <= 16'b0100010011001110;
            14'h1720 	:	o_val <= 16'b0100010011010000;
            14'h1721 	:	o_val <= 16'b0100010011010011;
            14'h1722 	:	o_val <= 16'b0100010011010110;
            14'h1723 	:	o_val <= 16'b0100010011011000;
            14'h1724 	:	o_val <= 16'b0100010011011011;
            14'h1725 	:	o_val <= 16'b0100010011011110;
            14'h1726 	:	o_val <= 16'b0100010011100000;
            14'h1727 	:	o_val <= 16'b0100010011100011;
            14'h1728 	:	o_val <= 16'b0100010011100110;
            14'h1729 	:	o_val <= 16'b0100010011101000;
            14'h172a 	:	o_val <= 16'b0100010011101011;
            14'h172b 	:	o_val <= 16'b0100010011101110;
            14'h172c 	:	o_val <= 16'b0100010011110000;
            14'h172d 	:	o_val <= 16'b0100010011110011;
            14'h172e 	:	o_val <= 16'b0100010011110110;
            14'h172f 	:	o_val <= 16'b0100010011111000;
            14'h1730 	:	o_val <= 16'b0100010011111011;
            14'h1731 	:	o_val <= 16'b0100010011111101;
            14'h1732 	:	o_val <= 16'b0100010100000000;
            14'h1733 	:	o_val <= 16'b0100010100000011;
            14'h1734 	:	o_val <= 16'b0100010100000101;
            14'h1735 	:	o_val <= 16'b0100010100001000;
            14'h1736 	:	o_val <= 16'b0100010100001011;
            14'h1737 	:	o_val <= 16'b0100010100001101;
            14'h1738 	:	o_val <= 16'b0100010100010000;
            14'h1739 	:	o_val <= 16'b0100010100010011;
            14'h173a 	:	o_val <= 16'b0100010100010101;
            14'h173b 	:	o_val <= 16'b0100010100011000;
            14'h173c 	:	o_val <= 16'b0100010100011011;
            14'h173d 	:	o_val <= 16'b0100010100011101;
            14'h173e 	:	o_val <= 16'b0100010100100000;
            14'h173f 	:	o_val <= 16'b0100010100100011;
            14'h1740 	:	o_val <= 16'b0100010100100101;
            14'h1741 	:	o_val <= 16'b0100010100101000;
            14'h1742 	:	o_val <= 16'b0100010100101010;
            14'h1743 	:	o_val <= 16'b0100010100101101;
            14'h1744 	:	o_val <= 16'b0100010100110000;
            14'h1745 	:	o_val <= 16'b0100010100110010;
            14'h1746 	:	o_val <= 16'b0100010100110101;
            14'h1747 	:	o_val <= 16'b0100010100111000;
            14'h1748 	:	o_val <= 16'b0100010100111010;
            14'h1749 	:	o_val <= 16'b0100010100111101;
            14'h174a 	:	o_val <= 16'b0100010101000000;
            14'h174b 	:	o_val <= 16'b0100010101000010;
            14'h174c 	:	o_val <= 16'b0100010101000101;
            14'h174d 	:	o_val <= 16'b0100010101001000;
            14'h174e 	:	o_val <= 16'b0100010101001010;
            14'h174f 	:	o_val <= 16'b0100010101001101;
            14'h1750 	:	o_val <= 16'b0100010101001111;
            14'h1751 	:	o_val <= 16'b0100010101010010;
            14'h1752 	:	o_val <= 16'b0100010101010101;
            14'h1753 	:	o_val <= 16'b0100010101010111;
            14'h1754 	:	o_val <= 16'b0100010101011010;
            14'h1755 	:	o_val <= 16'b0100010101011101;
            14'h1756 	:	o_val <= 16'b0100010101011111;
            14'h1757 	:	o_val <= 16'b0100010101100010;
            14'h1758 	:	o_val <= 16'b0100010101100101;
            14'h1759 	:	o_val <= 16'b0100010101100111;
            14'h175a 	:	o_val <= 16'b0100010101101010;
            14'h175b 	:	o_val <= 16'b0100010101101100;
            14'h175c 	:	o_val <= 16'b0100010101101111;
            14'h175d 	:	o_val <= 16'b0100010101110010;
            14'h175e 	:	o_val <= 16'b0100010101110100;
            14'h175f 	:	o_val <= 16'b0100010101110111;
            14'h1760 	:	o_val <= 16'b0100010101111010;
            14'h1761 	:	o_val <= 16'b0100010101111100;
            14'h1762 	:	o_val <= 16'b0100010101111111;
            14'h1763 	:	o_val <= 16'b0100010110000010;
            14'h1764 	:	o_val <= 16'b0100010110000100;
            14'h1765 	:	o_val <= 16'b0100010110000111;
            14'h1766 	:	o_val <= 16'b0100010110001010;
            14'h1767 	:	o_val <= 16'b0100010110001100;
            14'h1768 	:	o_val <= 16'b0100010110001111;
            14'h1769 	:	o_val <= 16'b0100010110010001;
            14'h176a 	:	o_val <= 16'b0100010110010100;
            14'h176b 	:	o_val <= 16'b0100010110010111;
            14'h176c 	:	o_val <= 16'b0100010110011001;
            14'h176d 	:	o_val <= 16'b0100010110011100;
            14'h176e 	:	o_val <= 16'b0100010110011111;
            14'h176f 	:	o_val <= 16'b0100010110100001;
            14'h1770 	:	o_val <= 16'b0100010110100100;
            14'h1771 	:	o_val <= 16'b0100010110100111;
            14'h1772 	:	o_val <= 16'b0100010110101001;
            14'h1773 	:	o_val <= 16'b0100010110101100;
            14'h1774 	:	o_val <= 16'b0100010110101110;
            14'h1775 	:	o_val <= 16'b0100010110110001;
            14'h1776 	:	o_val <= 16'b0100010110110100;
            14'h1777 	:	o_val <= 16'b0100010110110110;
            14'h1778 	:	o_val <= 16'b0100010110111001;
            14'h1779 	:	o_val <= 16'b0100010110111100;
            14'h177a 	:	o_val <= 16'b0100010110111110;
            14'h177b 	:	o_val <= 16'b0100010111000001;
            14'h177c 	:	o_val <= 16'b0100010111000011;
            14'h177d 	:	o_val <= 16'b0100010111000110;
            14'h177e 	:	o_val <= 16'b0100010111001001;
            14'h177f 	:	o_val <= 16'b0100010111001011;
            14'h1780 	:	o_val <= 16'b0100010111001110;
            14'h1781 	:	o_val <= 16'b0100010111010001;
            14'h1782 	:	o_val <= 16'b0100010111010011;
            14'h1783 	:	o_val <= 16'b0100010111010110;
            14'h1784 	:	o_val <= 16'b0100010111011001;
            14'h1785 	:	o_val <= 16'b0100010111011011;
            14'h1786 	:	o_val <= 16'b0100010111011110;
            14'h1787 	:	o_val <= 16'b0100010111100000;
            14'h1788 	:	o_val <= 16'b0100010111100011;
            14'h1789 	:	o_val <= 16'b0100010111100110;
            14'h178a 	:	o_val <= 16'b0100010111101000;
            14'h178b 	:	o_val <= 16'b0100010111101011;
            14'h178c 	:	o_val <= 16'b0100010111101110;
            14'h178d 	:	o_val <= 16'b0100010111110000;
            14'h178e 	:	o_val <= 16'b0100010111110011;
            14'h178f 	:	o_val <= 16'b0100010111110110;
            14'h1790 	:	o_val <= 16'b0100010111111000;
            14'h1791 	:	o_val <= 16'b0100010111111011;
            14'h1792 	:	o_val <= 16'b0100010111111101;
            14'h1793 	:	o_val <= 16'b0100011000000000;
            14'h1794 	:	o_val <= 16'b0100011000000011;
            14'h1795 	:	o_val <= 16'b0100011000000101;
            14'h1796 	:	o_val <= 16'b0100011000001000;
            14'h1797 	:	o_val <= 16'b0100011000001011;
            14'h1798 	:	o_val <= 16'b0100011000001101;
            14'h1799 	:	o_val <= 16'b0100011000010000;
            14'h179a 	:	o_val <= 16'b0100011000010010;
            14'h179b 	:	o_val <= 16'b0100011000010101;
            14'h179c 	:	o_val <= 16'b0100011000011000;
            14'h179d 	:	o_val <= 16'b0100011000011010;
            14'h179e 	:	o_val <= 16'b0100011000011101;
            14'h179f 	:	o_val <= 16'b0100011000100000;
            14'h17a0 	:	o_val <= 16'b0100011000100010;
            14'h17a1 	:	o_val <= 16'b0100011000100101;
            14'h17a2 	:	o_val <= 16'b0100011000100111;
            14'h17a3 	:	o_val <= 16'b0100011000101010;
            14'h17a4 	:	o_val <= 16'b0100011000101101;
            14'h17a5 	:	o_val <= 16'b0100011000101111;
            14'h17a6 	:	o_val <= 16'b0100011000110010;
            14'h17a7 	:	o_val <= 16'b0100011000110101;
            14'h17a8 	:	o_val <= 16'b0100011000110111;
            14'h17a9 	:	o_val <= 16'b0100011000111010;
            14'h17aa 	:	o_val <= 16'b0100011000111100;
            14'h17ab 	:	o_val <= 16'b0100011000111111;
            14'h17ac 	:	o_val <= 16'b0100011001000010;
            14'h17ad 	:	o_val <= 16'b0100011001000100;
            14'h17ae 	:	o_val <= 16'b0100011001000111;
            14'h17af 	:	o_val <= 16'b0100011001001010;
            14'h17b0 	:	o_val <= 16'b0100011001001100;
            14'h17b1 	:	o_val <= 16'b0100011001001111;
            14'h17b2 	:	o_val <= 16'b0100011001010001;
            14'h17b3 	:	o_val <= 16'b0100011001010100;
            14'h17b4 	:	o_val <= 16'b0100011001010111;
            14'h17b5 	:	o_val <= 16'b0100011001011001;
            14'h17b6 	:	o_val <= 16'b0100011001011100;
            14'h17b7 	:	o_val <= 16'b0100011001011111;
            14'h17b8 	:	o_val <= 16'b0100011001100001;
            14'h17b9 	:	o_val <= 16'b0100011001100100;
            14'h17ba 	:	o_val <= 16'b0100011001100110;
            14'h17bb 	:	o_val <= 16'b0100011001101001;
            14'h17bc 	:	o_val <= 16'b0100011001101100;
            14'h17bd 	:	o_val <= 16'b0100011001101110;
            14'h17be 	:	o_val <= 16'b0100011001110001;
            14'h17bf 	:	o_val <= 16'b0100011001110100;
            14'h17c0 	:	o_val <= 16'b0100011001110110;
            14'h17c1 	:	o_val <= 16'b0100011001111001;
            14'h17c2 	:	o_val <= 16'b0100011001111011;
            14'h17c3 	:	o_val <= 16'b0100011001111110;
            14'h17c4 	:	o_val <= 16'b0100011010000001;
            14'h17c5 	:	o_val <= 16'b0100011010000011;
            14'h17c6 	:	o_val <= 16'b0100011010000110;
            14'h17c7 	:	o_val <= 16'b0100011010001001;
            14'h17c8 	:	o_val <= 16'b0100011010001011;
            14'h17c9 	:	o_val <= 16'b0100011010001110;
            14'h17ca 	:	o_val <= 16'b0100011010010000;
            14'h17cb 	:	o_val <= 16'b0100011010010011;
            14'h17cc 	:	o_val <= 16'b0100011010010110;
            14'h17cd 	:	o_val <= 16'b0100011010011000;
            14'h17ce 	:	o_val <= 16'b0100011010011011;
            14'h17cf 	:	o_val <= 16'b0100011010011110;
            14'h17d0 	:	o_val <= 16'b0100011010100000;
            14'h17d1 	:	o_val <= 16'b0100011010100011;
            14'h17d2 	:	o_val <= 16'b0100011010100101;
            14'h17d3 	:	o_val <= 16'b0100011010101000;
            14'h17d4 	:	o_val <= 16'b0100011010101011;
            14'h17d5 	:	o_val <= 16'b0100011010101101;
            14'h17d6 	:	o_val <= 16'b0100011010110000;
            14'h17d7 	:	o_val <= 16'b0100011010110010;
            14'h17d8 	:	o_val <= 16'b0100011010110101;
            14'h17d9 	:	o_val <= 16'b0100011010111000;
            14'h17da 	:	o_val <= 16'b0100011010111010;
            14'h17db 	:	o_val <= 16'b0100011010111101;
            14'h17dc 	:	o_val <= 16'b0100011011000000;
            14'h17dd 	:	o_val <= 16'b0100011011000010;
            14'h17de 	:	o_val <= 16'b0100011011000101;
            14'h17df 	:	o_val <= 16'b0100011011000111;
            14'h17e0 	:	o_val <= 16'b0100011011001010;
            14'h17e1 	:	o_val <= 16'b0100011011001101;
            14'h17e2 	:	o_val <= 16'b0100011011001111;
            14'h17e3 	:	o_val <= 16'b0100011011010010;
            14'h17e4 	:	o_val <= 16'b0100011011010101;
            14'h17e5 	:	o_val <= 16'b0100011011010111;
            14'h17e6 	:	o_val <= 16'b0100011011011010;
            14'h17e7 	:	o_val <= 16'b0100011011011100;
            14'h17e8 	:	o_val <= 16'b0100011011011111;
            14'h17e9 	:	o_val <= 16'b0100011011100010;
            14'h17ea 	:	o_val <= 16'b0100011011100100;
            14'h17eb 	:	o_val <= 16'b0100011011100111;
            14'h17ec 	:	o_val <= 16'b0100011011101001;
            14'h17ed 	:	o_val <= 16'b0100011011101100;
            14'h17ee 	:	o_val <= 16'b0100011011101111;
            14'h17ef 	:	o_val <= 16'b0100011011110001;
            14'h17f0 	:	o_val <= 16'b0100011011110100;
            14'h17f1 	:	o_val <= 16'b0100011011110111;
            14'h17f2 	:	o_val <= 16'b0100011011111001;
            14'h17f3 	:	o_val <= 16'b0100011011111100;
            14'h17f4 	:	o_val <= 16'b0100011011111110;
            14'h17f5 	:	o_val <= 16'b0100011100000001;
            14'h17f6 	:	o_val <= 16'b0100011100000100;
            14'h17f7 	:	o_val <= 16'b0100011100000110;
            14'h17f8 	:	o_val <= 16'b0100011100001001;
            14'h17f9 	:	o_val <= 16'b0100011100001011;
            14'h17fa 	:	o_val <= 16'b0100011100001110;
            14'h17fb 	:	o_val <= 16'b0100011100010001;
            14'h17fc 	:	o_val <= 16'b0100011100010011;
            14'h17fd 	:	o_val <= 16'b0100011100010110;
            14'h17fe 	:	o_val <= 16'b0100011100011001;
            14'h17ff 	:	o_val <= 16'b0100011100011011;
            14'h1800 	:	o_val <= 16'b0100011100011110;
            14'h1801 	:	o_val <= 16'b0100011100100000;
            14'h1802 	:	o_val <= 16'b0100011100100011;
            14'h1803 	:	o_val <= 16'b0100011100100110;
            14'h1804 	:	o_val <= 16'b0100011100101000;
            14'h1805 	:	o_val <= 16'b0100011100101011;
            14'h1806 	:	o_val <= 16'b0100011100101101;
            14'h1807 	:	o_val <= 16'b0100011100110000;
            14'h1808 	:	o_val <= 16'b0100011100110011;
            14'h1809 	:	o_val <= 16'b0100011100110101;
            14'h180a 	:	o_val <= 16'b0100011100111000;
            14'h180b 	:	o_val <= 16'b0100011100111010;
            14'h180c 	:	o_val <= 16'b0100011100111101;
            14'h180d 	:	o_val <= 16'b0100011101000000;
            14'h180e 	:	o_val <= 16'b0100011101000010;
            14'h180f 	:	o_val <= 16'b0100011101000101;
            14'h1810 	:	o_val <= 16'b0100011101001000;
            14'h1811 	:	o_val <= 16'b0100011101001010;
            14'h1812 	:	o_val <= 16'b0100011101001101;
            14'h1813 	:	o_val <= 16'b0100011101001111;
            14'h1814 	:	o_val <= 16'b0100011101010010;
            14'h1815 	:	o_val <= 16'b0100011101010101;
            14'h1816 	:	o_val <= 16'b0100011101010111;
            14'h1817 	:	o_val <= 16'b0100011101011010;
            14'h1818 	:	o_val <= 16'b0100011101011100;
            14'h1819 	:	o_val <= 16'b0100011101011111;
            14'h181a 	:	o_val <= 16'b0100011101100010;
            14'h181b 	:	o_val <= 16'b0100011101100100;
            14'h181c 	:	o_val <= 16'b0100011101100111;
            14'h181d 	:	o_val <= 16'b0100011101101001;
            14'h181e 	:	o_val <= 16'b0100011101101100;
            14'h181f 	:	o_val <= 16'b0100011101101111;
            14'h1820 	:	o_val <= 16'b0100011101110001;
            14'h1821 	:	o_val <= 16'b0100011101110100;
            14'h1822 	:	o_val <= 16'b0100011101110110;
            14'h1823 	:	o_val <= 16'b0100011101111001;
            14'h1824 	:	o_val <= 16'b0100011101111100;
            14'h1825 	:	o_val <= 16'b0100011101111110;
            14'h1826 	:	o_val <= 16'b0100011110000001;
            14'h1827 	:	o_val <= 16'b0100011110000011;
            14'h1828 	:	o_val <= 16'b0100011110000110;
            14'h1829 	:	o_val <= 16'b0100011110001001;
            14'h182a 	:	o_val <= 16'b0100011110001011;
            14'h182b 	:	o_val <= 16'b0100011110001110;
            14'h182c 	:	o_val <= 16'b0100011110010000;
            14'h182d 	:	o_val <= 16'b0100011110010011;
            14'h182e 	:	o_val <= 16'b0100011110010110;
            14'h182f 	:	o_val <= 16'b0100011110011000;
            14'h1830 	:	o_val <= 16'b0100011110011011;
            14'h1831 	:	o_val <= 16'b0100011110011110;
            14'h1832 	:	o_val <= 16'b0100011110100000;
            14'h1833 	:	o_val <= 16'b0100011110100011;
            14'h1834 	:	o_val <= 16'b0100011110100101;
            14'h1835 	:	o_val <= 16'b0100011110101000;
            14'h1836 	:	o_val <= 16'b0100011110101011;
            14'h1837 	:	o_val <= 16'b0100011110101101;
            14'h1838 	:	o_val <= 16'b0100011110110000;
            14'h1839 	:	o_val <= 16'b0100011110110010;
            14'h183a 	:	o_val <= 16'b0100011110110101;
            14'h183b 	:	o_val <= 16'b0100011110111000;
            14'h183c 	:	o_val <= 16'b0100011110111010;
            14'h183d 	:	o_val <= 16'b0100011110111101;
            14'h183e 	:	o_val <= 16'b0100011110111111;
            14'h183f 	:	o_val <= 16'b0100011111000010;
            14'h1840 	:	o_val <= 16'b0100011111000101;
            14'h1841 	:	o_val <= 16'b0100011111000111;
            14'h1842 	:	o_val <= 16'b0100011111001010;
            14'h1843 	:	o_val <= 16'b0100011111001100;
            14'h1844 	:	o_val <= 16'b0100011111001111;
            14'h1845 	:	o_val <= 16'b0100011111010010;
            14'h1846 	:	o_val <= 16'b0100011111010100;
            14'h1847 	:	o_val <= 16'b0100011111010111;
            14'h1848 	:	o_val <= 16'b0100011111011001;
            14'h1849 	:	o_val <= 16'b0100011111011100;
            14'h184a 	:	o_val <= 16'b0100011111011111;
            14'h184b 	:	o_val <= 16'b0100011111100001;
            14'h184c 	:	o_val <= 16'b0100011111100100;
            14'h184d 	:	o_val <= 16'b0100011111100110;
            14'h184e 	:	o_val <= 16'b0100011111101001;
            14'h184f 	:	o_val <= 16'b0100011111101100;
            14'h1850 	:	o_val <= 16'b0100011111101110;
            14'h1851 	:	o_val <= 16'b0100011111110001;
            14'h1852 	:	o_val <= 16'b0100011111110011;
            14'h1853 	:	o_val <= 16'b0100011111110110;
            14'h1854 	:	o_val <= 16'b0100011111111001;
            14'h1855 	:	o_val <= 16'b0100011111111011;
            14'h1856 	:	o_val <= 16'b0100011111111110;
            14'h1857 	:	o_val <= 16'b0100100000000000;
            14'h1858 	:	o_val <= 16'b0100100000000011;
            14'h1859 	:	o_val <= 16'b0100100000000110;
            14'h185a 	:	o_val <= 16'b0100100000001000;
            14'h185b 	:	o_val <= 16'b0100100000001011;
            14'h185c 	:	o_val <= 16'b0100100000001101;
            14'h185d 	:	o_val <= 16'b0100100000010000;
            14'h185e 	:	o_val <= 16'b0100100000010011;
            14'h185f 	:	o_val <= 16'b0100100000010101;
            14'h1860 	:	o_val <= 16'b0100100000011000;
            14'h1861 	:	o_val <= 16'b0100100000011010;
            14'h1862 	:	o_val <= 16'b0100100000011101;
            14'h1863 	:	o_val <= 16'b0100100000100000;
            14'h1864 	:	o_val <= 16'b0100100000100010;
            14'h1865 	:	o_val <= 16'b0100100000100101;
            14'h1866 	:	o_val <= 16'b0100100000100111;
            14'h1867 	:	o_val <= 16'b0100100000101010;
            14'h1868 	:	o_val <= 16'b0100100000101100;
            14'h1869 	:	o_val <= 16'b0100100000101111;
            14'h186a 	:	o_val <= 16'b0100100000110010;
            14'h186b 	:	o_val <= 16'b0100100000110100;
            14'h186c 	:	o_val <= 16'b0100100000110111;
            14'h186d 	:	o_val <= 16'b0100100000111001;
            14'h186e 	:	o_val <= 16'b0100100000111100;
            14'h186f 	:	o_val <= 16'b0100100000111111;
            14'h1870 	:	o_val <= 16'b0100100001000001;
            14'h1871 	:	o_val <= 16'b0100100001000100;
            14'h1872 	:	o_val <= 16'b0100100001000110;
            14'h1873 	:	o_val <= 16'b0100100001001001;
            14'h1874 	:	o_val <= 16'b0100100001001100;
            14'h1875 	:	o_val <= 16'b0100100001001110;
            14'h1876 	:	o_val <= 16'b0100100001010001;
            14'h1877 	:	o_val <= 16'b0100100001010011;
            14'h1878 	:	o_val <= 16'b0100100001010110;
            14'h1879 	:	o_val <= 16'b0100100001011001;
            14'h187a 	:	o_val <= 16'b0100100001011011;
            14'h187b 	:	o_val <= 16'b0100100001011110;
            14'h187c 	:	o_val <= 16'b0100100001100000;
            14'h187d 	:	o_val <= 16'b0100100001100011;
            14'h187e 	:	o_val <= 16'b0100100001100110;
            14'h187f 	:	o_val <= 16'b0100100001101000;
            14'h1880 	:	o_val <= 16'b0100100001101011;
            14'h1881 	:	o_val <= 16'b0100100001101101;
            14'h1882 	:	o_val <= 16'b0100100001110000;
            14'h1883 	:	o_val <= 16'b0100100001110010;
            14'h1884 	:	o_val <= 16'b0100100001110101;
            14'h1885 	:	o_val <= 16'b0100100001111000;
            14'h1886 	:	o_val <= 16'b0100100001111010;
            14'h1887 	:	o_val <= 16'b0100100001111101;
            14'h1888 	:	o_val <= 16'b0100100001111111;
            14'h1889 	:	o_val <= 16'b0100100010000010;
            14'h188a 	:	o_val <= 16'b0100100010000101;
            14'h188b 	:	o_val <= 16'b0100100010000111;
            14'h188c 	:	o_val <= 16'b0100100010001010;
            14'h188d 	:	o_val <= 16'b0100100010001100;
            14'h188e 	:	o_val <= 16'b0100100010001111;
            14'h188f 	:	o_val <= 16'b0100100010010010;
            14'h1890 	:	o_val <= 16'b0100100010010100;
            14'h1891 	:	o_val <= 16'b0100100010010111;
            14'h1892 	:	o_val <= 16'b0100100010011001;
            14'h1893 	:	o_val <= 16'b0100100010011100;
            14'h1894 	:	o_val <= 16'b0100100010011110;
            14'h1895 	:	o_val <= 16'b0100100010100001;
            14'h1896 	:	o_val <= 16'b0100100010100100;
            14'h1897 	:	o_val <= 16'b0100100010100110;
            14'h1898 	:	o_val <= 16'b0100100010101001;
            14'h1899 	:	o_val <= 16'b0100100010101011;
            14'h189a 	:	o_val <= 16'b0100100010101110;
            14'h189b 	:	o_val <= 16'b0100100010110001;
            14'h189c 	:	o_val <= 16'b0100100010110011;
            14'h189d 	:	o_val <= 16'b0100100010110110;
            14'h189e 	:	o_val <= 16'b0100100010111000;
            14'h189f 	:	o_val <= 16'b0100100010111011;
            14'h18a0 	:	o_val <= 16'b0100100010111110;
            14'h18a1 	:	o_val <= 16'b0100100011000000;
            14'h18a2 	:	o_val <= 16'b0100100011000011;
            14'h18a3 	:	o_val <= 16'b0100100011000101;
            14'h18a4 	:	o_val <= 16'b0100100011001000;
            14'h18a5 	:	o_val <= 16'b0100100011001010;
            14'h18a6 	:	o_val <= 16'b0100100011001101;
            14'h18a7 	:	o_val <= 16'b0100100011010000;
            14'h18a8 	:	o_val <= 16'b0100100011010010;
            14'h18a9 	:	o_val <= 16'b0100100011010101;
            14'h18aa 	:	o_val <= 16'b0100100011010111;
            14'h18ab 	:	o_val <= 16'b0100100011011010;
            14'h18ac 	:	o_val <= 16'b0100100011011101;
            14'h18ad 	:	o_val <= 16'b0100100011011111;
            14'h18ae 	:	o_val <= 16'b0100100011100010;
            14'h18af 	:	o_val <= 16'b0100100011100100;
            14'h18b0 	:	o_val <= 16'b0100100011100111;
            14'h18b1 	:	o_val <= 16'b0100100011101001;
            14'h18b2 	:	o_val <= 16'b0100100011101100;
            14'h18b3 	:	o_val <= 16'b0100100011101111;
            14'h18b4 	:	o_val <= 16'b0100100011110001;
            14'h18b5 	:	o_val <= 16'b0100100011110100;
            14'h18b6 	:	o_val <= 16'b0100100011110110;
            14'h18b7 	:	o_val <= 16'b0100100011111001;
            14'h18b8 	:	o_val <= 16'b0100100011111011;
            14'h18b9 	:	o_val <= 16'b0100100011111110;
            14'h18ba 	:	o_val <= 16'b0100100100000001;
            14'h18bb 	:	o_val <= 16'b0100100100000011;
            14'h18bc 	:	o_val <= 16'b0100100100000110;
            14'h18bd 	:	o_val <= 16'b0100100100001000;
            14'h18be 	:	o_val <= 16'b0100100100001011;
            14'h18bf 	:	o_val <= 16'b0100100100001110;
            14'h18c0 	:	o_val <= 16'b0100100100010000;
            14'h18c1 	:	o_val <= 16'b0100100100010011;
            14'h18c2 	:	o_val <= 16'b0100100100010101;
            14'h18c3 	:	o_val <= 16'b0100100100011000;
            14'h18c4 	:	o_val <= 16'b0100100100011010;
            14'h18c5 	:	o_val <= 16'b0100100100011101;
            14'h18c6 	:	o_val <= 16'b0100100100100000;
            14'h18c7 	:	o_val <= 16'b0100100100100010;
            14'h18c8 	:	o_val <= 16'b0100100100100101;
            14'h18c9 	:	o_val <= 16'b0100100100100111;
            14'h18ca 	:	o_val <= 16'b0100100100101010;
            14'h18cb 	:	o_val <= 16'b0100100100101100;
            14'h18cc 	:	o_val <= 16'b0100100100101111;
            14'h18cd 	:	o_val <= 16'b0100100100110010;
            14'h18ce 	:	o_val <= 16'b0100100100110100;
            14'h18cf 	:	o_val <= 16'b0100100100110111;
            14'h18d0 	:	o_val <= 16'b0100100100111001;
            14'h18d1 	:	o_val <= 16'b0100100100111100;
            14'h18d2 	:	o_val <= 16'b0100100100111111;
            14'h18d3 	:	o_val <= 16'b0100100101000001;
            14'h18d4 	:	o_val <= 16'b0100100101000100;
            14'h18d5 	:	o_val <= 16'b0100100101000110;
            14'h18d6 	:	o_val <= 16'b0100100101001001;
            14'h18d7 	:	o_val <= 16'b0100100101001011;
            14'h18d8 	:	o_val <= 16'b0100100101001110;
            14'h18d9 	:	o_val <= 16'b0100100101010001;
            14'h18da 	:	o_val <= 16'b0100100101010011;
            14'h18db 	:	o_val <= 16'b0100100101010110;
            14'h18dc 	:	o_val <= 16'b0100100101011000;
            14'h18dd 	:	o_val <= 16'b0100100101011011;
            14'h18de 	:	o_val <= 16'b0100100101011101;
            14'h18df 	:	o_val <= 16'b0100100101100000;
            14'h18e0 	:	o_val <= 16'b0100100101100011;
            14'h18e1 	:	o_val <= 16'b0100100101100101;
            14'h18e2 	:	o_val <= 16'b0100100101101000;
            14'h18e3 	:	o_val <= 16'b0100100101101010;
            14'h18e4 	:	o_val <= 16'b0100100101101101;
            14'h18e5 	:	o_val <= 16'b0100100101101111;
            14'h18e6 	:	o_val <= 16'b0100100101110010;
            14'h18e7 	:	o_val <= 16'b0100100101110101;
            14'h18e8 	:	o_val <= 16'b0100100101110111;
            14'h18e9 	:	o_val <= 16'b0100100101111010;
            14'h18ea 	:	o_val <= 16'b0100100101111100;
            14'h18eb 	:	o_val <= 16'b0100100101111111;
            14'h18ec 	:	o_val <= 16'b0100100110000001;
            14'h18ed 	:	o_val <= 16'b0100100110000100;
            14'h18ee 	:	o_val <= 16'b0100100110000111;
            14'h18ef 	:	o_val <= 16'b0100100110001001;
            14'h18f0 	:	o_val <= 16'b0100100110001100;
            14'h18f1 	:	o_val <= 16'b0100100110001110;
            14'h18f2 	:	o_val <= 16'b0100100110010001;
            14'h18f3 	:	o_val <= 16'b0100100110010011;
            14'h18f4 	:	o_val <= 16'b0100100110010110;
            14'h18f5 	:	o_val <= 16'b0100100110011001;
            14'h18f6 	:	o_val <= 16'b0100100110011011;
            14'h18f7 	:	o_val <= 16'b0100100110011110;
            14'h18f8 	:	o_val <= 16'b0100100110100000;
            14'h18f9 	:	o_val <= 16'b0100100110100011;
            14'h18fa 	:	o_val <= 16'b0100100110100101;
            14'h18fb 	:	o_val <= 16'b0100100110101000;
            14'h18fc 	:	o_val <= 16'b0100100110101011;
            14'h18fd 	:	o_val <= 16'b0100100110101101;
            14'h18fe 	:	o_val <= 16'b0100100110110000;
            14'h18ff 	:	o_val <= 16'b0100100110110010;
            14'h1900 	:	o_val <= 16'b0100100110110101;
            14'h1901 	:	o_val <= 16'b0100100110110111;
            14'h1902 	:	o_val <= 16'b0100100110111010;
            14'h1903 	:	o_val <= 16'b0100100110111101;
            14'h1904 	:	o_val <= 16'b0100100110111111;
            14'h1905 	:	o_val <= 16'b0100100111000010;
            14'h1906 	:	o_val <= 16'b0100100111000100;
            14'h1907 	:	o_val <= 16'b0100100111000111;
            14'h1908 	:	o_val <= 16'b0100100111001001;
            14'h1909 	:	o_val <= 16'b0100100111001100;
            14'h190a 	:	o_val <= 16'b0100100111001111;
            14'h190b 	:	o_val <= 16'b0100100111010001;
            14'h190c 	:	o_val <= 16'b0100100111010100;
            14'h190d 	:	o_val <= 16'b0100100111010110;
            14'h190e 	:	o_val <= 16'b0100100111011001;
            14'h190f 	:	o_val <= 16'b0100100111011011;
            14'h1910 	:	o_val <= 16'b0100100111011110;
            14'h1911 	:	o_val <= 16'b0100100111100001;
            14'h1912 	:	o_val <= 16'b0100100111100011;
            14'h1913 	:	o_val <= 16'b0100100111100110;
            14'h1914 	:	o_val <= 16'b0100100111101000;
            14'h1915 	:	o_val <= 16'b0100100111101011;
            14'h1916 	:	o_val <= 16'b0100100111101101;
            14'h1917 	:	o_val <= 16'b0100100111110000;
            14'h1918 	:	o_val <= 16'b0100100111110010;
            14'h1919 	:	o_val <= 16'b0100100111110101;
            14'h191a 	:	o_val <= 16'b0100100111111000;
            14'h191b 	:	o_val <= 16'b0100100111111010;
            14'h191c 	:	o_val <= 16'b0100100111111101;
            14'h191d 	:	o_val <= 16'b0100100111111111;
            14'h191e 	:	o_val <= 16'b0100101000000010;
            14'h191f 	:	o_val <= 16'b0100101000000100;
            14'h1920 	:	o_val <= 16'b0100101000000111;
            14'h1921 	:	o_val <= 16'b0100101000001010;
            14'h1922 	:	o_val <= 16'b0100101000001100;
            14'h1923 	:	o_val <= 16'b0100101000001111;
            14'h1924 	:	o_val <= 16'b0100101000010001;
            14'h1925 	:	o_val <= 16'b0100101000010100;
            14'h1926 	:	o_val <= 16'b0100101000010110;
            14'h1927 	:	o_val <= 16'b0100101000011001;
            14'h1928 	:	o_val <= 16'b0100101000011011;
            14'h1929 	:	o_val <= 16'b0100101000011110;
            14'h192a 	:	o_val <= 16'b0100101000100001;
            14'h192b 	:	o_val <= 16'b0100101000100011;
            14'h192c 	:	o_val <= 16'b0100101000100110;
            14'h192d 	:	o_val <= 16'b0100101000101000;
            14'h192e 	:	o_val <= 16'b0100101000101011;
            14'h192f 	:	o_val <= 16'b0100101000101101;
            14'h1930 	:	o_val <= 16'b0100101000110000;
            14'h1931 	:	o_val <= 16'b0100101000110011;
            14'h1932 	:	o_val <= 16'b0100101000110101;
            14'h1933 	:	o_val <= 16'b0100101000111000;
            14'h1934 	:	o_val <= 16'b0100101000111010;
            14'h1935 	:	o_val <= 16'b0100101000111101;
            14'h1936 	:	o_val <= 16'b0100101000111111;
            14'h1937 	:	o_val <= 16'b0100101001000010;
            14'h1938 	:	o_val <= 16'b0100101001000100;
            14'h1939 	:	o_val <= 16'b0100101001000111;
            14'h193a 	:	o_val <= 16'b0100101001001010;
            14'h193b 	:	o_val <= 16'b0100101001001100;
            14'h193c 	:	o_val <= 16'b0100101001001111;
            14'h193d 	:	o_val <= 16'b0100101001010001;
            14'h193e 	:	o_val <= 16'b0100101001010100;
            14'h193f 	:	o_val <= 16'b0100101001010110;
            14'h1940 	:	o_val <= 16'b0100101001011001;
            14'h1941 	:	o_val <= 16'b0100101001011011;
            14'h1942 	:	o_val <= 16'b0100101001011110;
            14'h1943 	:	o_val <= 16'b0100101001100001;
            14'h1944 	:	o_val <= 16'b0100101001100011;
            14'h1945 	:	o_val <= 16'b0100101001100110;
            14'h1946 	:	o_val <= 16'b0100101001101000;
            14'h1947 	:	o_val <= 16'b0100101001101011;
            14'h1948 	:	o_val <= 16'b0100101001101101;
            14'h1949 	:	o_val <= 16'b0100101001110000;
            14'h194a 	:	o_val <= 16'b0100101001110010;
            14'h194b 	:	o_val <= 16'b0100101001110101;
            14'h194c 	:	o_val <= 16'b0100101001111000;
            14'h194d 	:	o_val <= 16'b0100101001111010;
            14'h194e 	:	o_val <= 16'b0100101001111101;
            14'h194f 	:	o_val <= 16'b0100101001111111;
            14'h1950 	:	o_val <= 16'b0100101010000010;
            14'h1951 	:	o_val <= 16'b0100101010000100;
            14'h1952 	:	o_val <= 16'b0100101010000111;
            14'h1953 	:	o_val <= 16'b0100101010001001;
            14'h1954 	:	o_val <= 16'b0100101010001100;
            14'h1955 	:	o_val <= 16'b0100101010001111;
            14'h1956 	:	o_val <= 16'b0100101010010001;
            14'h1957 	:	o_val <= 16'b0100101010010100;
            14'h1958 	:	o_val <= 16'b0100101010010110;
            14'h1959 	:	o_val <= 16'b0100101010011001;
            14'h195a 	:	o_val <= 16'b0100101010011011;
            14'h195b 	:	o_val <= 16'b0100101010011110;
            14'h195c 	:	o_val <= 16'b0100101010100000;
            14'h195d 	:	o_val <= 16'b0100101010100011;
            14'h195e 	:	o_val <= 16'b0100101010100110;
            14'h195f 	:	o_val <= 16'b0100101010101000;
            14'h1960 	:	o_val <= 16'b0100101010101011;
            14'h1961 	:	o_val <= 16'b0100101010101101;
            14'h1962 	:	o_val <= 16'b0100101010110000;
            14'h1963 	:	o_val <= 16'b0100101010110010;
            14'h1964 	:	o_val <= 16'b0100101010110101;
            14'h1965 	:	o_val <= 16'b0100101010110111;
            14'h1966 	:	o_val <= 16'b0100101010111010;
            14'h1967 	:	o_val <= 16'b0100101010111100;
            14'h1968 	:	o_val <= 16'b0100101010111111;
            14'h1969 	:	o_val <= 16'b0100101011000010;
            14'h196a 	:	o_val <= 16'b0100101011000100;
            14'h196b 	:	o_val <= 16'b0100101011000111;
            14'h196c 	:	o_val <= 16'b0100101011001001;
            14'h196d 	:	o_val <= 16'b0100101011001100;
            14'h196e 	:	o_val <= 16'b0100101011001110;
            14'h196f 	:	o_val <= 16'b0100101011010001;
            14'h1970 	:	o_val <= 16'b0100101011010011;
            14'h1971 	:	o_val <= 16'b0100101011010110;
            14'h1972 	:	o_val <= 16'b0100101011011001;
            14'h1973 	:	o_val <= 16'b0100101011011011;
            14'h1974 	:	o_val <= 16'b0100101011011110;
            14'h1975 	:	o_val <= 16'b0100101011100000;
            14'h1976 	:	o_val <= 16'b0100101011100011;
            14'h1977 	:	o_val <= 16'b0100101011100101;
            14'h1978 	:	o_val <= 16'b0100101011101000;
            14'h1979 	:	o_val <= 16'b0100101011101010;
            14'h197a 	:	o_val <= 16'b0100101011101101;
            14'h197b 	:	o_val <= 16'b0100101011101111;
            14'h197c 	:	o_val <= 16'b0100101011110010;
            14'h197d 	:	o_val <= 16'b0100101011110101;
            14'h197e 	:	o_val <= 16'b0100101011110111;
            14'h197f 	:	o_val <= 16'b0100101011111010;
            14'h1980 	:	o_val <= 16'b0100101011111100;
            14'h1981 	:	o_val <= 16'b0100101011111111;
            14'h1982 	:	o_val <= 16'b0100101100000001;
            14'h1983 	:	o_val <= 16'b0100101100000100;
            14'h1984 	:	o_val <= 16'b0100101100000110;
            14'h1985 	:	o_val <= 16'b0100101100001001;
            14'h1986 	:	o_val <= 16'b0100101100001011;
            14'h1987 	:	o_val <= 16'b0100101100001110;
            14'h1988 	:	o_val <= 16'b0100101100010001;
            14'h1989 	:	o_val <= 16'b0100101100010011;
            14'h198a 	:	o_val <= 16'b0100101100010110;
            14'h198b 	:	o_val <= 16'b0100101100011000;
            14'h198c 	:	o_val <= 16'b0100101100011011;
            14'h198d 	:	o_val <= 16'b0100101100011101;
            14'h198e 	:	o_val <= 16'b0100101100100000;
            14'h198f 	:	o_val <= 16'b0100101100100010;
            14'h1990 	:	o_val <= 16'b0100101100100101;
            14'h1991 	:	o_val <= 16'b0100101100100111;
            14'h1992 	:	o_val <= 16'b0100101100101010;
            14'h1993 	:	o_val <= 16'b0100101100101101;
            14'h1994 	:	o_val <= 16'b0100101100101111;
            14'h1995 	:	o_val <= 16'b0100101100110010;
            14'h1996 	:	o_val <= 16'b0100101100110100;
            14'h1997 	:	o_val <= 16'b0100101100110111;
            14'h1998 	:	o_val <= 16'b0100101100111001;
            14'h1999 	:	o_val <= 16'b0100101100111100;
            14'h199a 	:	o_val <= 16'b0100101100111110;
            14'h199b 	:	o_val <= 16'b0100101101000001;
            14'h199c 	:	o_val <= 16'b0100101101000011;
            14'h199d 	:	o_val <= 16'b0100101101000110;
            14'h199e 	:	o_val <= 16'b0100101101001000;
            14'h199f 	:	o_val <= 16'b0100101101001011;
            14'h19a0 	:	o_val <= 16'b0100101101001110;
            14'h19a1 	:	o_val <= 16'b0100101101010000;
            14'h19a2 	:	o_val <= 16'b0100101101010011;
            14'h19a3 	:	o_val <= 16'b0100101101010101;
            14'h19a4 	:	o_val <= 16'b0100101101011000;
            14'h19a5 	:	o_val <= 16'b0100101101011010;
            14'h19a6 	:	o_val <= 16'b0100101101011101;
            14'h19a7 	:	o_val <= 16'b0100101101011111;
            14'h19a8 	:	o_val <= 16'b0100101101100010;
            14'h19a9 	:	o_val <= 16'b0100101101100100;
            14'h19aa 	:	o_val <= 16'b0100101101100111;
            14'h19ab 	:	o_val <= 16'b0100101101101010;
            14'h19ac 	:	o_val <= 16'b0100101101101100;
            14'h19ad 	:	o_val <= 16'b0100101101101111;
            14'h19ae 	:	o_val <= 16'b0100101101110001;
            14'h19af 	:	o_val <= 16'b0100101101110100;
            14'h19b0 	:	o_val <= 16'b0100101101110110;
            14'h19b1 	:	o_val <= 16'b0100101101111001;
            14'h19b2 	:	o_val <= 16'b0100101101111011;
            14'h19b3 	:	o_val <= 16'b0100101101111110;
            14'h19b4 	:	o_val <= 16'b0100101110000000;
            14'h19b5 	:	o_val <= 16'b0100101110000011;
            14'h19b6 	:	o_val <= 16'b0100101110000101;
            14'h19b7 	:	o_val <= 16'b0100101110001000;
            14'h19b8 	:	o_val <= 16'b0100101110001010;
            14'h19b9 	:	o_val <= 16'b0100101110001101;
            14'h19ba 	:	o_val <= 16'b0100101110010000;
            14'h19bb 	:	o_val <= 16'b0100101110010010;
            14'h19bc 	:	o_val <= 16'b0100101110010101;
            14'h19bd 	:	o_val <= 16'b0100101110010111;
            14'h19be 	:	o_val <= 16'b0100101110011010;
            14'h19bf 	:	o_val <= 16'b0100101110011100;
            14'h19c0 	:	o_val <= 16'b0100101110011111;
            14'h19c1 	:	o_val <= 16'b0100101110100001;
            14'h19c2 	:	o_val <= 16'b0100101110100100;
            14'h19c3 	:	o_val <= 16'b0100101110100110;
            14'h19c4 	:	o_val <= 16'b0100101110101001;
            14'h19c5 	:	o_val <= 16'b0100101110101011;
            14'h19c6 	:	o_val <= 16'b0100101110101110;
            14'h19c7 	:	o_val <= 16'b0100101110110001;
            14'h19c8 	:	o_val <= 16'b0100101110110011;
            14'h19c9 	:	o_val <= 16'b0100101110110110;
            14'h19ca 	:	o_val <= 16'b0100101110111000;
            14'h19cb 	:	o_val <= 16'b0100101110111011;
            14'h19cc 	:	o_val <= 16'b0100101110111101;
            14'h19cd 	:	o_val <= 16'b0100101111000000;
            14'h19ce 	:	o_val <= 16'b0100101111000010;
            14'h19cf 	:	o_val <= 16'b0100101111000101;
            14'h19d0 	:	o_val <= 16'b0100101111000111;
            14'h19d1 	:	o_val <= 16'b0100101111001010;
            14'h19d2 	:	o_val <= 16'b0100101111001100;
            14'h19d3 	:	o_val <= 16'b0100101111001111;
            14'h19d4 	:	o_val <= 16'b0100101111010001;
            14'h19d5 	:	o_val <= 16'b0100101111010100;
            14'h19d6 	:	o_val <= 16'b0100101111010111;
            14'h19d7 	:	o_val <= 16'b0100101111011001;
            14'h19d8 	:	o_val <= 16'b0100101111011100;
            14'h19d9 	:	o_val <= 16'b0100101111011110;
            14'h19da 	:	o_val <= 16'b0100101111100001;
            14'h19db 	:	o_val <= 16'b0100101111100011;
            14'h19dc 	:	o_val <= 16'b0100101111100110;
            14'h19dd 	:	o_val <= 16'b0100101111101000;
            14'h19de 	:	o_val <= 16'b0100101111101011;
            14'h19df 	:	o_val <= 16'b0100101111101101;
            14'h19e0 	:	o_val <= 16'b0100101111110000;
            14'h19e1 	:	o_val <= 16'b0100101111110010;
            14'h19e2 	:	o_val <= 16'b0100101111110101;
            14'h19e3 	:	o_val <= 16'b0100101111110111;
            14'h19e4 	:	o_val <= 16'b0100101111111010;
            14'h19e5 	:	o_val <= 16'b0100101111111100;
            14'h19e6 	:	o_val <= 16'b0100101111111111;
            14'h19e7 	:	o_val <= 16'b0100110000000001;
            14'h19e8 	:	o_val <= 16'b0100110000000100;
            14'h19e9 	:	o_val <= 16'b0100110000000111;
            14'h19ea 	:	o_val <= 16'b0100110000001001;
            14'h19eb 	:	o_val <= 16'b0100110000001100;
            14'h19ec 	:	o_val <= 16'b0100110000001110;
            14'h19ed 	:	o_val <= 16'b0100110000010001;
            14'h19ee 	:	o_val <= 16'b0100110000010011;
            14'h19ef 	:	o_val <= 16'b0100110000010110;
            14'h19f0 	:	o_val <= 16'b0100110000011000;
            14'h19f1 	:	o_val <= 16'b0100110000011011;
            14'h19f2 	:	o_val <= 16'b0100110000011101;
            14'h19f3 	:	o_val <= 16'b0100110000100000;
            14'h19f4 	:	o_val <= 16'b0100110000100010;
            14'h19f5 	:	o_val <= 16'b0100110000100101;
            14'h19f6 	:	o_val <= 16'b0100110000100111;
            14'h19f7 	:	o_val <= 16'b0100110000101010;
            14'h19f8 	:	o_val <= 16'b0100110000101100;
            14'h19f9 	:	o_val <= 16'b0100110000101111;
            14'h19fa 	:	o_val <= 16'b0100110000110001;
            14'h19fb 	:	o_val <= 16'b0100110000110100;
            14'h19fc 	:	o_val <= 16'b0100110000110111;
            14'h19fd 	:	o_val <= 16'b0100110000111001;
            14'h19fe 	:	o_val <= 16'b0100110000111100;
            14'h19ff 	:	o_val <= 16'b0100110000111110;
            14'h1a00 	:	o_val <= 16'b0100110001000001;
            14'h1a01 	:	o_val <= 16'b0100110001000011;
            14'h1a02 	:	o_val <= 16'b0100110001000110;
            14'h1a03 	:	o_val <= 16'b0100110001001000;
            14'h1a04 	:	o_val <= 16'b0100110001001011;
            14'h1a05 	:	o_val <= 16'b0100110001001101;
            14'h1a06 	:	o_val <= 16'b0100110001010000;
            14'h1a07 	:	o_val <= 16'b0100110001010010;
            14'h1a08 	:	o_val <= 16'b0100110001010101;
            14'h1a09 	:	o_val <= 16'b0100110001010111;
            14'h1a0a 	:	o_val <= 16'b0100110001011010;
            14'h1a0b 	:	o_val <= 16'b0100110001011100;
            14'h1a0c 	:	o_val <= 16'b0100110001011111;
            14'h1a0d 	:	o_val <= 16'b0100110001100001;
            14'h1a0e 	:	o_val <= 16'b0100110001100100;
            14'h1a0f 	:	o_val <= 16'b0100110001100110;
            14'h1a10 	:	o_val <= 16'b0100110001101001;
            14'h1a11 	:	o_val <= 16'b0100110001101100;
            14'h1a12 	:	o_val <= 16'b0100110001101110;
            14'h1a13 	:	o_val <= 16'b0100110001110001;
            14'h1a14 	:	o_val <= 16'b0100110001110011;
            14'h1a15 	:	o_val <= 16'b0100110001110110;
            14'h1a16 	:	o_val <= 16'b0100110001111000;
            14'h1a17 	:	o_val <= 16'b0100110001111011;
            14'h1a18 	:	o_val <= 16'b0100110001111101;
            14'h1a19 	:	o_val <= 16'b0100110010000000;
            14'h1a1a 	:	o_val <= 16'b0100110010000010;
            14'h1a1b 	:	o_val <= 16'b0100110010000101;
            14'h1a1c 	:	o_val <= 16'b0100110010000111;
            14'h1a1d 	:	o_val <= 16'b0100110010001010;
            14'h1a1e 	:	o_val <= 16'b0100110010001100;
            14'h1a1f 	:	o_val <= 16'b0100110010001111;
            14'h1a20 	:	o_val <= 16'b0100110010010001;
            14'h1a21 	:	o_val <= 16'b0100110010010100;
            14'h1a22 	:	o_val <= 16'b0100110010010110;
            14'h1a23 	:	o_val <= 16'b0100110010011001;
            14'h1a24 	:	o_val <= 16'b0100110010011011;
            14'h1a25 	:	o_val <= 16'b0100110010011110;
            14'h1a26 	:	o_val <= 16'b0100110010100000;
            14'h1a27 	:	o_val <= 16'b0100110010100011;
            14'h1a28 	:	o_val <= 16'b0100110010100101;
            14'h1a29 	:	o_val <= 16'b0100110010101000;
            14'h1a2a 	:	o_val <= 16'b0100110010101010;
            14'h1a2b 	:	o_val <= 16'b0100110010101101;
            14'h1a2c 	:	o_val <= 16'b0100110010101111;
            14'h1a2d 	:	o_val <= 16'b0100110010110010;
            14'h1a2e 	:	o_val <= 16'b0100110010110101;
            14'h1a2f 	:	o_val <= 16'b0100110010110111;
            14'h1a30 	:	o_val <= 16'b0100110010111010;
            14'h1a31 	:	o_val <= 16'b0100110010111100;
            14'h1a32 	:	o_val <= 16'b0100110010111111;
            14'h1a33 	:	o_val <= 16'b0100110011000001;
            14'h1a34 	:	o_val <= 16'b0100110011000100;
            14'h1a35 	:	o_val <= 16'b0100110011000110;
            14'h1a36 	:	o_val <= 16'b0100110011001001;
            14'h1a37 	:	o_val <= 16'b0100110011001011;
            14'h1a38 	:	o_val <= 16'b0100110011001110;
            14'h1a39 	:	o_val <= 16'b0100110011010000;
            14'h1a3a 	:	o_val <= 16'b0100110011010011;
            14'h1a3b 	:	o_val <= 16'b0100110011010101;
            14'h1a3c 	:	o_val <= 16'b0100110011011000;
            14'h1a3d 	:	o_val <= 16'b0100110011011010;
            14'h1a3e 	:	o_val <= 16'b0100110011011101;
            14'h1a3f 	:	o_val <= 16'b0100110011011111;
            14'h1a40 	:	o_val <= 16'b0100110011100010;
            14'h1a41 	:	o_val <= 16'b0100110011100100;
            14'h1a42 	:	o_val <= 16'b0100110011100111;
            14'h1a43 	:	o_val <= 16'b0100110011101001;
            14'h1a44 	:	o_val <= 16'b0100110011101100;
            14'h1a45 	:	o_val <= 16'b0100110011101110;
            14'h1a46 	:	o_val <= 16'b0100110011110001;
            14'h1a47 	:	o_val <= 16'b0100110011110011;
            14'h1a48 	:	o_val <= 16'b0100110011110110;
            14'h1a49 	:	o_val <= 16'b0100110011111000;
            14'h1a4a 	:	o_val <= 16'b0100110011111011;
            14'h1a4b 	:	o_val <= 16'b0100110011111101;
            14'h1a4c 	:	o_val <= 16'b0100110100000000;
            14'h1a4d 	:	o_val <= 16'b0100110100000010;
            14'h1a4e 	:	o_val <= 16'b0100110100000101;
            14'h1a4f 	:	o_val <= 16'b0100110100000111;
            14'h1a50 	:	o_val <= 16'b0100110100001010;
            14'h1a51 	:	o_val <= 16'b0100110100001100;
            14'h1a52 	:	o_val <= 16'b0100110100001111;
            14'h1a53 	:	o_val <= 16'b0100110100010001;
            14'h1a54 	:	o_val <= 16'b0100110100010100;
            14'h1a55 	:	o_val <= 16'b0100110100010110;
            14'h1a56 	:	o_val <= 16'b0100110100011001;
            14'h1a57 	:	o_val <= 16'b0100110100011011;
            14'h1a58 	:	o_val <= 16'b0100110100011110;
            14'h1a59 	:	o_val <= 16'b0100110100100000;
            14'h1a5a 	:	o_val <= 16'b0100110100100011;
            14'h1a5b 	:	o_val <= 16'b0100110100100110;
            14'h1a5c 	:	o_val <= 16'b0100110100101000;
            14'h1a5d 	:	o_val <= 16'b0100110100101011;
            14'h1a5e 	:	o_val <= 16'b0100110100101101;
            14'h1a5f 	:	o_val <= 16'b0100110100110000;
            14'h1a60 	:	o_val <= 16'b0100110100110010;
            14'h1a61 	:	o_val <= 16'b0100110100110101;
            14'h1a62 	:	o_val <= 16'b0100110100110111;
            14'h1a63 	:	o_val <= 16'b0100110100111010;
            14'h1a64 	:	o_val <= 16'b0100110100111100;
            14'h1a65 	:	o_val <= 16'b0100110100111111;
            14'h1a66 	:	o_val <= 16'b0100110101000001;
            14'h1a67 	:	o_val <= 16'b0100110101000100;
            14'h1a68 	:	o_val <= 16'b0100110101000110;
            14'h1a69 	:	o_val <= 16'b0100110101001001;
            14'h1a6a 	:	o_val <= 16'b0100110101001011;
            14'h1a6b 	:	o_val <= 16'b0100110101001110;
            14'h1a6c 	:	o_val <= 16'b0100110101010000;
            14'h1a6d 	:	o_val <= 16'b0100110101010011;
            14'h1a6e 	:	o_val <= 16'b0100110101010101;
            14'h1a6f 	:	o_val <= 16'b0100110101011000;
            14'h1a70 	:	o_val <= 16'b0100110101011010;
            14'h1a71 	:	o_val <= 16'b0100110101011101;
            14'h1a72 	:	o_val <= 16'b0100110101011111;
            14'h1a73 	:	o_val <= 16'b0100110101100010;
            14'h1a74 	:	o_val <= 16'b0100110101100100;
            14'h1a75 	:	o_val <= 16'b0100110101100111;
            14'h1a76 	:	o_val <= 16'b0100110101101001;
            14'h1a77 	:	o_val <= 16'b0100110101101100;
            14'h1a78 	:	o_val <= 16'b0100110101101110;
            14'h1a79 	:	o_val <= 16'b0100110101110001;
            14'h1a7a 	:	o_val <= 16'b0100110101110011;
            14'h1a7b 	:	o_val <= 16'b0100110101110110;
            14'h1a7c 	:	o_val <= 16'b0100110101111000;
            14'h1a7d 	:	o_val <= 16'b0100110101111011;
            14'h1a7e 	:	o_val <= 16'b0100110101111101;
            14'h1a7f 	:	o_val <= 16'b0100110110000000;
            14'h1a80 	:	o_val <= 16'b0100110110000010;
            14'h1a81 	:	o_val <= 16'b0100110110000101;
            14'h1a82 	:	o_val <= 16'b0100110110000111;
            14'h1a83 	:	o_val <= 16'b0100110110001010;
            14'h1a84 	:	o_val <= 16'b0100110110001100;
            14'h1a85 	:	o_val <= 16'b0100110110001111;
            14'h1a86 	:	o_val <= 16'b0100110110010001;
            14'h1a87 	:	o_val <= 16'b0100110110010100;
            14'h1a88 	:	o_val <= 16'b0100110110010110;
            14'h1a89 	:	o_val <= 16'b0100110110011001;
            14'h1a8a 	:	o_val <= 16'b0100110110011011;
            14'h1a8b 	:	o_val <= 16'b0100110110011110;
            14'h1a8c 	:	o_val <= 16'b0100110110100000;
            14'h1a8d 	:	o_val <= 16'b0100110110100011;
            14'h1a8e 	:	o_val <= 16'b0100110110100101;
            14'h1a8f 	:	o_val <= 16'b0100110110101000;
            14'h1a90 	:	o_val <= 16'b0100110110101010;
            14'h1a91 	:	o_val <= 16'b0100110110101101;
            14'h1a92 	:	o_val <= 16'b0100110110101111;
            14'h1a93 	:	o_val <= 16'b0100110110110010;
            14'h1a94 	:	o_val <= 16'b0100110110110100;
            14'h1a95 	:	o_val <= 16'b0100110110110111;
            14'h1a96 	:	o_val <= 16'b0100110110111001;
            14'h1a97 	:	o_val <= 16'b0100110110111100;
            14'h1a98 	:	o_val <= 16'b0100110110111110;
            14'h1a99 	:	o_val <= 16'b0100110111000001;
            14'h1a9a 	:	o_val <= 16'b0100110111000011;
            14'h1a9b 	:	o_val <= 16'b0100110111000110;
            14'h1a9c 	:	o_val <= 16'b0100110111001000;
            14'h1a9d 	:	o_val <= 16'b0100110111001011;
            14'h1a9e 	:	o_val <= 16'b0100110111001101;
            14'h1a9f 	:	o_val <= 16'b0100110111010000;
            14'h1aa0 	:	o_val <= 16'b0100110111010010;
            14'h1aa1 	:	o_val <= 16'b0100110111010101;
            14'h1aa2 	:	o_val <= 16'b0100110111010111;
            14'h1aa3 	:	o_val <= 16'b0100110111011010;
            14'h1aa4 	:	o_val <= 16'b0100110111011100;
            14'h1aa5 	:	o_val <= 16'b0100110111011111;
            14'h1aa6 	:	o_val <= 16'b0100110111100001;
            14'h1aa7 	:	o_val <= 16'b0100110111100100;
            14'h1aa8 	:	o_val <= 16'b0100110111100110;
            14'h1aa9 	:	o_val <= 16'b0100110111101000;
            14'h1aaa 	:	o_val <= 16'b0100110111101011;
            14'h1aab 	:	o_val <= 16'b0100110111101101;
            14'h1aac 	:	o_val <= 16'b0100110111110000;
            14'h1aad 	:	o_val <= 16'b0100110111110010;
            14'h1aae 	:	o_val <= 16'b0100110111110101;
            14'h1aaf 	:	o_val <= 16'b0100110111110111;
            14'h1ab0 	:	o_val <= 16'b0100110111111010;
            14'h1ab1 	:	o_val <= 16'b0100110111111100;
            14'h1ab2 	:	o_val <= 16'b0100110111111111;
            14'h1ab3 	:	o_val <= 16'b0100111000000001;
            14'h1ab4 	:	o_val <= 16'b0100111000000100;
            14'h1ab5 	:	o_val <= 16'b0100111000000110;
            14'h1ab6 	:	o_val <= 16'b0100111000001001;
            14'h1ab7 	:	o_val <= 16'b0100111000001011;
            14'h1ab8 	:	o_val <= 16'b0100111000001110;
            14'h1ab9 	:	o_val <= 16'b0100111000010000;
            14'h1aba 	:	o_val <= 16'b0100111000010011;
            14'h1abb 	:	o_val <= 16'b0100111000010101;
            14'h1abc 	:	o_val <= 16'b0100111000011000;
            14'h1abd 	:	o_val <= 16'b0100111000011010;
            14'h1abe 	:	o_val <= 16'b0100111000011101;
            14'h1abf 	:	o_val <= 16'b0100111000011111;
            14'h1ac0 	:	o_val <= 16'b0100111000100010;
            14'h1ac1 	:	o_val <= 16'b0100111000100100;
            14'h1ac2 	:	o_val <= 16'b0100111000100111;
            14'h1ac3 	:	o_val <= 16'b0100111000101001;
            14'h1ac4 	:	o_val <= 16'b0100111000101100;
            14'h1ac5 	:	o_val <= 16'b0100111000101110;
            14'h1ac6 	:	o_val <= 16'b0100111000110001;
            14'h1ac7 	:	o_val <= 16'b0100111000110011;
            14'h1ac8 	:	o_val <= 16'b0100111000110110;
            14'h1ac9 	:	o_val <= 16'b0100111000111000;
            14'h1aca 	:	o_val <= 16'b0100111000111011;
            14'h1acb 	:	o_val <= 16'b0100111000111101;
            14'h1acc 	:	o_val <= 16'b0100111001000000;
            14'h1acd 	:	o_val <= 16'b0100111001000010;
            14'h1ace 	:	o_val <= 16'b0100111001000101;
            14'h1acf 	:	o_val <= 16'b0100111001000111;
            14'h1ad0 	:	o_val <= 16'b0100111001001010;
            14'h1ad1 	:	o_val <= 16'b0100111001001100;
            14'h1ad2 	:	o_val <= 16'b0100111001001111;
            14'h1ad3 	:	o_val <= 16'b0100111001010001;
            14'h1ad4 	:	o_val <= 16'b0100111001010011;
            14'h1ad5 	:	o_val <= 16'b0100111001010110;
            14'h1ad6 	:	o_val <= 16'b0100111001011000;
            14'h1ad7 	:	o_val <= 16'b0100111001011011;
            14'h1ad8 	:	o_val <= 16'b0100111001011101;
            14'h1ad9 	:	o_val <= 16'b0100111001100000;
            14'h1ada 	:	o_val <= 16'b0100111001100010;
            14'h1adb 	:	o_val <= 16'b0100111001100101;
            14'h1adc 	:	o_val <= 16'b0100111001100111;
            14'h1add 	:	o_val <= 16'b0100111001101010;
            14'h1ade 	:	o_val <= 16'b0100111001101100;
            14'h1adf 	:	o_val <= 16'b0100111001101111;
            14'h1ae0 	:	o_val <= 16'b0100111001110001;
            14'h1ae1 	:	o_val <= 16'b0100111001110100;
            14'h1ae2 	:	o_val <= 16'b0100111001110110;
            14'h1ae3 	:	o_val <= 16'b0100111001111001;
            14'h1ae4 	:	o_val <= 16'b0100111001111011;
            14'h1ae5 	:	o_val <= 16'b0100111001111110;
            14'h1ae6 	:	o_val <= 16'b0100111010000000;
            14'h1ae7 	:	o_val <= 16'b0100111010000011;
            14'h1ae8 	:	o_val <= 16'b0100111010000101;
            14'h1ae9 	:	o_val <= 16'b0100111010001000;
            14'h1aea 	:	o_val <= 16'b0100111010001010;
            14'h1aeb 	:	o_val <= 16'b0100111010001101;
            14'h1aec 	:	o_val <= 16'b0100111010001111;
            14'h1aed 	:	o_val <= 16'b0100111010010010;
            14'h1aee 	:	o_val <= 16'b0100111010010100;
            14'h1aef 	:	o_val <= 16'b0100111010010111;
            14'h1af0 	:	o_val <= 16'b0100111010011001;
            14'h1af1 	:	o_val <= 16'b0100111010011011;
            14'h1af2 	:	o_val <= 16'b0100111010011110;
            14'h1af3 	:	o_val <= 16'b0100111010100000;
            14'h1af4 	:	o_val <= 16'b0100111010100011;
            14'h1af5 	:	o_val <= 16'b0100111010100101;
            14'h1af6 	:	o_val <= 16'b0100111010101000;
            14'h1af7 	:	o_val <= 16'b0100111010101010;
            14'h1af8 	:	o_val <= 16'b0100111010101101;
            14'h1af9 	:	o_val <= 16'b0100111010101111;
            14'h1afa 	:	o_val <= 16'b0100111010110010;
            14'h1afb 	:	o_val <= 16'b0100111010110100;
            14'h1afc 	:	o_val <= 16'b0100111010110111;
            14'h1afd 	:	o_val <= 16'b0100111010111001;
            14'h1afe 	:	o_val <= 16'b0100111010111100;
            14'h1aff 	:	o_val <= 16'b0100111010111110;
            14'h1b00 	:	o_val <= 16'b0100111011000001;
            14'h1b01 	:	o_val <= 16'b0100111011000011;
            14'h1b02 	:	o_val <= 16'b0100111011000110;
            14'h1b03 	:	o_val <= 16'b0100111011001000;
            14'h1b04 	:	o_val <= 16'b0100111011001011;
            14'h1b05 	:	o_val <= 16'b0100111011001101;
            14'h1b06 	:	o_val <= 16'b0100111011010000;
            14'h1b07 	:	o_val <= 16'b0100111011010010;
            14'h1b08 	:	o_val <= 16'b0100111011010100;
            14'h1b09 	:	o_val <= 16'b0100111011010111;
            14'h1b0a 	:	o_val <= 16'b0100111011011001;
            14'h1b0b 	:	o_val <= 16'b0100111011011100;
            14'h1b0c 	:	o_val <= 16'b0100111011011110;
            14'h1b0d 	:	o_val <= 16'b0100111011100001;
            14'h1b0e 	:	o_val <= 16'b0100111011100011;
            14'h1b0f 	:	o_val <= 16'b0100111011100110;
            14'h1b10 	:	o_val <= 16'b0100111011101000;
            14'h1b11 	:	o_val <= 16'b0100111011101011;
            14'h1b12 	:	o_val <= 16'b0100111011101101;
            14'h1b13 	:	o_val <= 16'b0100111011110000;
            14'h1b14 	:	o_val <= 16'b0100111011110010;
            14'h1b15 	:	o_val <= 16'b0100111011110101;
            14'h1b16 	:	o_val <= 16'b0100111011110111;
            14'h1b17 	:	o_val <= 16'b0100111011111010;
            14'h1b18 	:	o_val <= 16'b0100111011111100;
            14'h1b19 	:	o_val <= 16'b0100111011111111;
            14'h1b1a 	:	o_val <= 16'b0100111100000001;
            14'h1b1b 	:	o_val <= 16'b0100111100000011;
            14'h1b1c 	:	o_val <= 16'b0100111100000110;
            14'h1b1d 	:	o_val <= 16'b0100111100001000;
            14'h1b1e 	:	o_val <= 16'b0100111100001011;
            14'h1b1f 	:	o_val <= 16'b0100111100001101;
            14'h1b20 	:	o_val <= 16'b0100111100010000;
            14'h1b21 	:	o_val <= 16'b0100111100010010;
            14'h1b22 	:	o_val <= 16'b0100111100010101;
            14'h1b23 	:	o_val <= 16'b0100111100010111;
            14'h1b24 	:	o_val <= 16'b0100111100011010;
            14'h1b25 	:	o_val <= 16'b0100111100011100;
            14'h1b26 	:	o_val <= 16'b0100111100011111;
            14'h1b27 	:	o_val <= 16'b0100111100100001;
            14'h1b28 	:	o_val <= 16'b0100111100100100;
            14'h1b29 	:	o_val <= 16'b0100111100100110;
            14'h1b2a 	:	o_val <= 16'b0100111100101000;
            14'h1b2b 	:	o_val <= 16'b0100111100101011;
            14'h1b2c 	:	o_val <= 16'b0100111100101101;
            14'h1b2d 	:	o_val <= 16'b0100111100110000;
            14'h1b2e 	:	o_val <= 16'b0100111100110010;
            14'h1b2f 	:	o_val <= 16'b0100111100110101;
            14'h1b30 	:	o_val <= 16'b0100111100110111;
            14'h1b31 	:	o_val <= 16'b0100111100111010;
            14'h1b32 	:	o_val <= 16'b0100111100111100;
            14'h1b33 	:	o_val <= 16'b0100111100111111;
            14'h1b34 	:	o_val <= 16'b0100111101000001;
            14'h1b35 	:	o_val <= 16'b0100111101000100;
            14'h1b36 	:	o_val <= 16'b0100111101000110;
            14'h1b37 	:	o_val <= 16'b0100111101001001;
            14'h1b38 	:	o_val <= 16'b0100111101001011;
            14'h1b39 	:	o_val <= 16'b0100111101001110;
            14'h1b3a 	:	o_val <= 16'b0100111101010000;
            14'h1b3b 	:	o_val <= 16'b0100111101010010;
            14'h1b3c 	:	o_val <= 16'b0100111101010101;
            14'h1b3d 	:	o_val <= 16'b0100111101010111;
            14'h1b3e 	:	o_val <= 16'b0100111101011010;
            14'h1b3f 	:	o_val <= 16'b0100111101011100;
            14'h1b40 	:	o_val <= 16'b0100111101011111;
            14'h1b41 	:	o_val <= 16'b0100111101100001;
            14'h1b42 	:	o_val <= 16'b0100111101100100;
            14'h1b43 	:	o_val <= 16'b0100111101100110;
            14'h1b44 	:	o_val <= 16'b0100111101101001;
            14'h1b45 	:	o_val <= 16'b0100111101101011;
            14'h1b46 	:	o_val <= 16'b0100111101101110;
            14'h1b47 	:	o_val <= 16'b0100111101110000;
            14'h1b48 	:	o_val <= 16'b0100111101110010;
            14'h1b49 	:	o_val <= 16'b0100111101110101;
            14'h1b4a 	:	o_val <= 16'b0100111101110111;
            14'h1b4b 	:	o_val <= 16'b0100111101111010;
            14'h1b4c 	:	o_val <= 16'b0100111101111100;
            14'h1b4d 	:	o_val <= 16'b0100111101111111;
            14'h1b4e 	:	o_val <= 16'b0100111110000001;
            14'h1b4f 	:	o_val <= 16'b0100111110000100;
            14'h1b50 	:	o_val <= 16'b0100111110000110;
            14'h1b51 	:	o_val <= 16'b0100111110001001;
            14'h1b52 	:	o_val <= 16'b0100111110001011;
            14'h1b53 	:	o_val <= 16'b0100111110001110;
            14'h1b54 	:	o_val <= 16'b0100111110010000;
            14'h1b55 	:	o_val <= 16'b0100111110010010;
            14'h1b56 	:	o_val <= 16'b0100111110010101;
            14'h1b57 	:	o_val <= 16'b0100111110010111;
            14'h1b58 	:	o_val <= 16'b0100111110011010;
            14'h1b59 	:	o_val <= 16'b0100111110011100;
            14'h1b5a 	:	o_val <= 16'b0100111110011111;
            14'h1b5b 	:	o_val <= 16'b0100111110100001;
            14'h1b5c 	:	o_val <= 16'b0100111110100100;
            14'h1b5d 	:	o_val <= 16'b0100111110100110;
            14'h1b5e 	:	o_val <= 16'b0100111110101001;
            14'h1b5f 	:	o_val <= 16'b0100111110101011;
            14'h1b60 	:	o_val <= 16'b0100111110101110;
            14'h1b61 	:	o_val <= 16'b0100111110110000;
            14'h1b62 	:	o_val <= 16'b0100111110110010;
            14'h1b63 	:	o_val <= 16'b0100111110110101;
            14'h1b64 	:	o_val <= 16'b0100111110110111;
            14'h1b65 	:	o_val <= 16'b0100111110111010;
            14'h1b66 	:	o_val <= 16'b0100111110111100;
            14'h1b67 	:	o_val <= 16'b0100111110111111;
            14'h1b68 	:	o_val <= 16'b0100111111000001;
            14'h1b69 	:	o_val <= 16'b0100111111000100;
            14'h1b6a 	:	o_val <= 16'b0100111111000110;
            14'h1b6b 	:	o_val <= 16'b0100111111001001;
            14'h1b6c 	:	o_val <= 16'b0100111111001011;
            14'h1b6d 	:	o_val <= 16'b0100111111001101;
            14'h1b6e 	:	o_val <= 16'b0100111111010000;
            14'h1b6f 	:	o_val <= 16'b0100111111010010;
            14'h1b70 	:	o_val <= 16'b0100111111010101;
            14'h1b71 	:	o_val <= 16'b0100111111010111;
            14'h1b72 	:	o_val <= 16'b0100111111011010;
            14'h1b73 	:	o_val <= 16'b0100111111011100;
            14'h1b74 	:	o_val <= 16'b0100111111011111;
            14'h1b75 	:	o_val <= 16'b0100111111100001;
            14'h1b76 	:	o_val <= 16'b0100111111100100;
            14'h1b77 	:	o_val <= 16'b0100111111100110;
            14'h1b78 	:	o_val <= 16'b0100111111101000;
            14'h1b79 	:	o_val <= 16'b0100111111101011;
            14'h1b7a 	:	o_val <= 16'b0100111111101101;
            14'h1b7b 	:	o_val <= 16'b0100111111110000;
            14'h1b7c 	:	o_val <= 16'b0100111111110010;
            14'h1b7d 	:	o_val <= 16'b0100111111110101;
            14'h1b7e 	:	o_val <= 16'b0100111111110111;
            14'h1b7f 	:	o_val <= 16'b0100111111111010;
            14'h1b80 	:	o_val <= 16'b0100111111111100;
            14'h1b81 	:	o_val <= 16'b0100111111111111;
            14'h1b82 	:	o_val <= 16'b0101000000000001;
            14'h1b83 	:	o_val <= 16'b0101000000000011;
            14'h1b84 	:	o_val <= 16'b0101000000000110;
            14'h1b85 	:	o_val <= 16'b0101000000001000;
            14'h1b86 	:	o_val <= 16'b0101000000001011;
            14'h1b87 	:	o_val <= 16'b0101000000001101;
            14'h1b88 	:	o_val <= 16'b0101000000010000;
            14'h1b89 	:	o_val <= 16'b0101000000010010;
            14'h1b8a 	:	o_val <= 16'b0101000000010101;
            14'h1b8b 	:	o_val <= 16'b0101000000010111;
            14'h1b8c 	:	o_val <= 16'b0101000000011010;
            14'h1b8d 	:	o_val <= 16'b0101000000011100;
            14'h1b8e 	:	o_val <= 16'b0101000000011110;
            14'h1b8f 	:	o_val <= 16'b0101000000100001;
            14'h1b90 	:	o_val <= 16'b0101000000100011;
            14'h1b91 	:	o_val <= 16'b0101000000100110;
            14'h1b92 	:	o_val <= 16'b0101000000101000;
            14'h1b93 	:	o_val <= 16'b0101000000101011;
            14'h1b94 	:	o_val <= 16'b0101000000101101;
            14'h1b95 	:	o_val <= 16'b0101000000110000;
            14'h1b96 	:	o_val <= 16'b0101000000110010;
            14'h1b97 	:	o_val <= 16'b0101000000110100;
            14'h1b98 	:	o_val <= 16'b0101000000110111;
            14'h1b99 	:	o_val <= 16'b0101000000111001;
            14'h1b9a 	:	o_val <= 16'b0101000000111100;
            14'h1b9b 	:	o_val <= 16'b0101000000111110;
            14'h1b9c 	:	o_val <= 16'b0101000001000001;
            14'h1b9d 	:	o_val <= 16'b0101000001000011;
            14'h1b9e 	:	o_val <= 16'b0101000001000110;
            14'h1b9f 	:	o_val <= 16'b0101000001001000;
            14'h1ba0 	:	o_val <= 16'b0101000001001011;
            14'h1ba1 	:	o_val <= 16'b0101000001001101;
            14'h1ba2 	:	o_val <= 16'b0101000001001111;
            14'h1ba3 	:	o_val <= 16'b0101000001010010;
            14'h1ba4 	:	o_val <= 16'b0101000001010100;
            14'h1ba5 	:	o_val <= 16'b0101000001010111;
            14'h1ba6 	:	o_val <= 16'b0101000001011001;
            14'h1ba7 	:	o_val <= 16'b0101000001011100;
            14'h1ba8 	:	o_val <= 16'b0101000001011110;
            14'h1ba9 	:	o_val <= 16'b0101000001100001;
            14'h1baa 	:	o_val <= 16'b0101000001100011;
            14'h1bab 	:	o_val <= 16'b0101000001100101;
            14'h1bac 	:	o_val <= 16'b0101000001101000;
            14'h1bad 	:	o_val <= 16'b0101000001101010;
            14'h1bae 	:	o_val <= 16'b0101000001101101;
            14'h1baf 	:	o_val <= 16'b0101000001101111;
            14'h1bb0 	:	o_val <= 16'b0101000001110010;
            14'h1bb1 	:	o_val <= 16'b0101000001110100;
            14'h1bb2 	:	o_val <= 16'b0101000001110111;
            14'h1bb3 	:	o_val <= 16'b0101000001111001;
            14'h1bb4 	:	o_val <= 16'b0101000001111011;
            14'h1bb5 	:	o_val <= 16'b0101000001111110;
            14'h1bb6 	:	o_val <= 16'b0101000010000000;
            14'h1bb7 	:	o_val <= 16'b0101000010000011;
            14'h1bb8 	:	o_val <= 16'b0101000010000101;
            14'h1bb9 	:	o_val <= 16'b0101000010001000;
            14'h1bba 	:	o_val <= 16'b0101000010001010;
            14'h1bbb 	:	o_val <= 16'b0101000010001101;
            14'h1bbc 	:	o_val <= 16'b0101000010001111;
            14'h1bbd 	:	o_val <= 16'b0101000010010001;
            14'h1bbe 	:	o_val <= 16'b0101000010010100;
            14'h1bbf 	:	o_val <= 16'b0101000010010110;
            14'h1bc0 	:	o_val <= 16'b0101000010011001;
            14'h1bc1 	:	o_val <= 16'b0101000010011011;
            14'h1bc2 	:	o_val <= 16'b0101000010011110;
            14'h1bc3 	:	o_val <= 16'b0101000010100000;
            14'h1bc4 	:	o_val <= 16'b0101000010100010;
            14'h1bc5 	:	o_val <= 16'b0101000010100101;
            14'h1bc6 	:	o_val <= 16'b0101000010100111;
            14'h1bc7 	:	o_val <= 16'b0101000010101010;
            14'h1bc8 	:	o_val <= 16'b0101000010101100;
            14'h1bc9 	:	o_val <= 16'b0101000010101111;
            14'h1bca 	:	o_val <= 16'b0101000010110001;
            14'h1bcb 	:	o_val <= 16'b0101000010110100;
            14'h1bcc 	:	o_val <= 16'b0101000010110110;
            14'h1bcd 	:	o_val <= 16'b0101000010111000;
            14'h1bce 	:	o_val <= 16'b0101000010111011;
            14'h1bcf 	:	o_val <= 16'b0101000010111101;
            14'h1bd0 	:	o_val <= 16'b0101000011000000;
            14'h1bd1 	:	o_val <= 16'b0101000011000010;
            14'h1bd2 	:	o_val <= 16'b0101000011000101;
            14'h1bd3 	:	o_val <= 16'b0101000011000111;
            14'h1bd4 	:	o_val <= 16'b0101000011001001;
            14'h1bd5 	:	o_val <= 16'b0101000011001100;
            14'h1bd6 	:	o_val <= 16'b0101000011001110;
            14'h1bd7 	:	o_val <= 16'b0101000011010001;
            14'h1bd8 	:	o_val <= 16'b0101000011010011;
            14'h1bd9 	:	o_val <= 16'b0101000011010110;
            14'h1bda 	:	o_val <= 16'b0101000011011000;
            14'h1bdb 	:	o_val <= 16'b0101000011011011;
            14'h1bdc 	:	o_val <= 16'b0101000011011101;
            14'h1bdd 	:	o_val <= 16'b0101000011011111;
            14'h1bde 	:	o_val <= 16'b0101000011100010;
            14'h1bdf 	:	o_val <= 16'b0101000011100100;
            14'h1be0 	:	o_val <= 16'b0101000011100111;
            14'h1be1 	:	o_val <= 16'b0101000011101001;
            14'h1be2 	:	o_val <= 16'b0101000011101100;
            14'h1be3 	:	o_val <= 16'b0101000011101110;
            14'h1be4 	:	o_val <= 16'b0101000011110000;
            14'h1be5 	:	o_val <= 16'b0101000011110011;
            14'h1be6 	:	o_val <= 16'b0101000011110101;
            14'h1be7 	:	o_val <= 16'b0101000011111000;
            14'h1be8 	:	o_val <= 16'b0101000011111010;
            14'h1be9 	:	o_val <= 16'b0101000011111101;
            14'h1bea 	:	o_val <= 16'b0101000011111111;
            14'h1beb 	:	o_val <= 16'b0101000100000001;
            14'h1bec 	:	o_val <= 16'b0101000100000100;
            14'h1bed 	:	o_val <= 16'b0101000100000110;
            14'h1bee 	:	o_val <= 16'b0101000100001001;
            14'h1bef 	:	o_val <= 16'b0101000100001011;
            14'h1bf0 	:	o_val <= 16'b0101000100001110;
            14'h1bf1 	:	o_val <= 16'b0101000100010000;
            14'h1bf2 	:	o_val <= 16'b0101000100010010;
            14'h1bf3 	:	o_val <= 16'b0101000100010101;
            14'h1bf4 	:	o_val <= 16'b0101000100010111;
            14'h1bf5 	:	o_val <= 16'b0101000100011010;
            14'h1bf6 	:	o_val <= 16'b0101000100011100;
            14'h1bf7 	:	o_val <= 16'b0101000100011111;
            14'h1bf8 	:	o_val <= 16'b0101000100100001;
            14'h1bf9 	:	o_val <= 16'b0101000100100100;
            14'h1bfa 	:	o_val <= 16'b0101000100100110;
            14'h1bfb 	:	o_val <= 16'b0101000100101000;
            14'h1bfc 	:	o_val <= 16'b0101000100101011;
            14'h1bfd 	:	o_val <= 16'b0101000100101101;
            14'h1bfe 	:	o_val <= 16'b0101000100110000;
            14'h1bff 	:	o_val <= 16'b0101000100110010;
            14'h1c00 	:	o_val <= 16'b0101000100110101;
            14'h1c01 	:	o_val <= 16'b0101000100110111;
            14'h1c02 	:	o_val <= 16'b0101000100111001;
            14'h1c03 	:	o_val <= 16'b0101000100111100;
            14'h1c04 	:	o_val <= 16'b0101000100111110;
            14'h1c05 	:	o_val <= 16'b0101000101000001;
            14'h1c06 	:	o_val <= 16'b0101000101000011;
            14'h1c07 	:	o_val <= 16'b0101000101000110;
            14'h1c08 	:	o_val <= 16'b0101000101001000;
            14'h1c09 	:	o_val <= 16'b0101000101001010;
            14'h1c0a 	:	o_val <= 16'b0101000101001101;
            14'h1c0b 	:	o_val <= 16'b0101000101001111;
            14'h1c0c 	:	o_val <= 16'b0101000101010010;
            14'h1c0d 	:	o_val <= 16'b0101000101010100;
            14'h1c0e 	:	o_val <= 16'b0101000101010110;
            14'h1c0f 	:	o_val <= 16'b0101000101011001;
            14'h1c10 	:	o_val <= 16'b0101000101011011;
            14'h1c11 	:	o_val <= 16'b0101000101011110;
            14'h1c12 	:	o_val <= 16'b0101000101100000;
            14'h1c13 	:	o_val <= 16'b0101000101100011;
            14'h1c14 	:	o_val <= 16'b0101000101100101;
            14'h1c15 	:	o_val <= 16'b0101000101100111;
            14'h1c16 	:	o_val <= 16'b0101000101101010;
            14'h1c17 	:	o_val <= 16'b0101000101101100;
            14'h1c18 	:	o_val <= 16'b0101000101101111;
            14'h1c19 	:	o_val <= 16'b0101000101110001;
            14'h1c1a 	:	o_val <= 16'b0101000101110100;
            14'h1c1b 	:	o_val <= 16'b0101000101110110;
            14'h1c1c 	:	o_val <= 16'b0101000101111000;
            14'h1c1d 	:	o_val <= 16'b0101000101111011;
            14'h1c1e 	:	o_val <= 16'b0101000101111101;
            14'h1c1f 	:	o_val <= 16'b0101000110000000;
            14'h1c20 	:	o_val <= 16'b0101000110000010;
            14'h1c21 	:	o_val <= 16'b0101000110000101;
            14'h1c22 	:	o_val <= 16'b0101000110000111;
            14'h1c23 	:	o_val <= 16'b0101000110001001;
            14'h1c24 	:	o_val <= 16'b0101000110001100;
            14'h1c25 	:	o_val <= 16'b0101000110001110;
            14'h1c26 	:	o_val <= 16'b0101000110010001;
            14'h1c27 	:	o_val <= 16'b0101000110010011;
            14'h1c28 	:	o_val <= 16'b0101000110010101;
            14'h1c29 	:	o_val <= 16'b0101000110011000;
            14'h1c2a 	:	o_val <= 16'b0101000110011010;
            14'h1c2b 	:	o_val <= 16'b0101000110011101;
            14'h1c2c 	:	o_val <= 16'b0101000110011111;
            14'h1c2d 	:	o_val <= 16'b0101000110100010;
            14'h1c2e 	:	o_val <= 16'b0101000110100100;
            14'h1c2f 	:	o_val <= 16'b0101000110100110;
            14'h1c30 	:	o_val <= 16'b0101000110101001;
            14'h1c31 	:	o_val <= 16'b0101000110101011;
            14'h1c32 	:	o_val <= 16'b0101000110101110;
            14'h1c33 	:	o_val <= 16'b0101000110110000;
            14'h1c34 	:	o_val <= 16'b0101000110110011;
            14'h1c35 	:	o_val <= 16'b0101000110110101;
            14'h1c36 	:	o_val <= 16'b0101000110110111;
            14'h1c37 	:	o_val <= 16'b0101000110111010;
            14'h1c38 	:	o_val <= 16'b0101000110111100;
            14'h1c39 	:	o_val <= 16'b0101000110111111;
            14'h1c3a 	:	o_val <= 16'b0101000111000001;
            14'h1c3b 	:	o_val <= 16'b0101000111000011;
            14'h1c3c 	:	o_val <= 16'b0101000111000110;
            14'h1c3d 	:	o_val <= 16'b0101000111001000;
            14'h1c3e 	:	o_val <= 16'b0101000111001011;
            14'h1c3f 	:	o_val <= 16'b0101000111001101;
            14'h1c40 	:	o_val <= 16'b0101000111010000;
            14'h1c41 	:	o_val <= 16'b0101000111010010;
            14'h1c42 	:	o_val <= 16'b0101000111010100;
            14'h1c43 	:	o_val <= 16'b0101000111010111;
            14'h1c44 	:	o_val <= 16'b0101000111011001;
            14'h1c45 	:	o_val <= 16'b0101000111011100;
            14'h1c46 	:	o_val <= 16'b0101000111011110;
            14'h1c47 	:	o_val <= 16'b0101000111100000;
            14'h1c48 	:	o_val <= 16'b0101000111100011;
            14'h1c49 	:	o_val <= 16'b0101000111100101;
            14'h1c4a 	:	o_val <= 16'b0101000111101000;
            14'h1c4b 	:	o_val <= 16'b0101000111101010;
            14'h1c4c 	:	o_val <= 16'b0101000111101101;
            14'h1c4d 	:	o_val <= 16'b0101000111101111;
            14'h1c4e 	:	o_val <= 16'b0101000111110001;
            14'h1c4f 	:	o_val <= 16'b0101000111110100;
            14'h1c50 	:	o_val <= 16'b0101000111110110;
            14'h1c51 	:	o_val <= 16'b0101000111111001;
            14'h1c52 	:	o_val <= 16'b0101000111111011;
            14'h1c53 	:	o_val <= 16'b0101000111111101;
            14'h1c54 	:	o_val <= 16'b0101001000000000;
            14'h1c55 	:	o_val <= 16'b0101001000000010;
            14'h1c56 	:	o_val <= 16'b0101001000000101;
            14'h1c57 	:	o_val <= 16'b0101001000000111;
            14'h1c58 	:	o_val <= 16'b0101001000001001;
            14'h1c59 	:	o_val <= 16'b0101001000001100;
            14'h1c5a 	:	o_val <= 16'b0101001000001110;
            14'h1c5b 	:	o_val <= 16'b0101001000010001;
            14'h1c5c 	:	o_val <= 16'b0101001000010011;
            14'h1c5d 	:	o_val <= 16'b0101001000010110;
            14'h1c5e 	:	o_val <= 16'b0101001000011000;
            14'h1c5f 	:	o_val <= 16'b0101001000011010;
            14'h1c60 	:	o_val <= 16'b0101001000011101;
            14'h1c61 	:	o_val <= 16'b0101001000011111;
            14'h1c62 	:	o_val <= 16'b0101001000100010;
            14'h1c63 	:	o_val <= 16'b0101001000100100;
            14'h1c64 	:	o_val <= 16'b0101001000100110;
            14'h1c65 	:	o_val <= 16'b0101001000101001;
            14'h1c66 	:	o_val <= 16'b0101001000101011;
            14'h1c67 	:	o_val <= 16'b0101001000101110;
            14'h1c68 	:	o_val <= 16'b0101001000110000;
            14'h1c69 	:	o_val <= 16'b0101001000110010;
            14'h1c6a 	:	o_val <= 16'b0101001000110101;
            14'h1c6b 	:	o_val <= 16'b0101001000110111;
            14'h1c6c 	:	o_val <= 16'b0101001000111010;
            14'h1c6d 	:	o_val <= 16'b0101001000111100;
            14'h1c6e 	:	o_val <= 16'b0101001000111110;
            14'h1c6f 	:	o_val <= 16'b0101001001000001;
            14'h1c70 	:	o_val <= 16'b0101001001000011;
            14'h1c71 	:	o_val <= 16'b0101001001000110;
            14'h1c72 	:	o_val <= 16'b0101001001001000;
            14'h1c73 	:	o_val <= 16'b0101001001001011;
            14'h1c74 	:	o_val <= 16'b0101001001001101;
            14'h1c75 	:	o_val <= 16'b0101001001001111;
            14'h1c76 	:	o_val <= 16'b0101001001010010;
            14'h1c77 	:	o_val <= 16'b0101001001010100;
            14'h1c78 	:	o_val <= 16'b0101001001010111;
            14'h1c79 	:	o_val <= 16'b0101001001011001;
            14'h1c7a 	:	o_val <= 16'b0101001001011011;
            14'h1c7b 	:	o_val <= 16'b0101001001011110;
            14'h1c7c 	:	o_val <= 16'b0101001001100000;
            14'h1c7d 	:	o_val <= 16'b0101001001100011;
            14'h1c7e 	:	o_val <= 16'b0101001001100101;
            14'h1c7f 	:	o_val <= 16'b0101001001100111;
            14'h1c80 	:	o_val <= 16'b0101001001101010;
            14'h1c81 	:	o_val <= 16'b0101001001101100;
            14'h1c82 	:	o_val <= 16'b0101001001101111;
            14'h1c83 	:	o_val <= 16'b0101001001110001;
            14'h1c84 	:	o_val <= 16'b0101001001110011;
            14'h1c85 	:	o_val <= 16'b0101001001110110;
            14'h1c86 	:	o_val <= 16'b0101001001111000;
            14'h1c87 	:	o_val <= 16'b0101001001111011;
            14'h1c88 	:	o_val <= 16'b0101001001111101;
            14'h1c89 	:	o_val <= 16'b0101001001111111;
            14'h1c8a 	:	o_val <= 16'b0101001010000010;
            14'h1c8b 	:	o_val <= 16'b0101001010000100;
            14'h1c8c 	:	o_val <= 16'b0101001010000111;
            14'h1c8d 	:	o_val <= 16'b0101001010001001;
            14'h1c8e 	:	o_val <= 16'b0101001010001011;
            14'h1c8f 	:	o_val <= 16'b0101001010001110;
            14'h1c90 	:	o_val <= 16'b0101001010010000;
            14'h1c91 	:	o_val <= 16'b0101001010010011;
            14'h1c92 	:	o_val <= 16'b0101001010010101;
            14'h1c93 	:	o_val <= 16'b0101001010010111;
            14'h1c94 	:	o_val <= 16'b0101001010011010;
            14'h1c95 	:	o_val <= 16'b0101001010011100;
            14'h1c96 	:	o_val <= 16'b0101001010011111;
            14'h1c97 	:	o_val <= 16'b0101001010100001;
            14'h1c98 	:	o_val <= 16'b0101001010100011;
            14'h1c99 	:	o_val <= 16'b0101001010100110;
            14'h1c9a 	:	o_val <= 16'b0101001010101000;
            14'h1c9b 	:	o_val <= 16'b0101001010101011;
            14'h1c9c 	:	o_val <= 16'b0101001010101101;
            14'h1c9d 	:	o_val <= 16'b0101001010101111;
            14'h1c9e 	:	o_val <= 16'b0101001010110010;
            14'h1c9f 	:	o_val <= 16'b0101001010110100;
            14'h1ca0 	:	o_val <= 16'b0101001010110111;
            14'h1ca1 	:	o_val <= 16'b0101001010111001;
            14'h1ca2 	:	o_val <= 16'b0101001010111011;
            14'h1ca3 	:	o_val <= 16'b0101001010111110;
            14'h1ca4 	:	o_val <= 16'b0101001011000000;
            14'h1ca5 	:	o_val <= 16'b0101001011000011;
            14'h1ca6 	:	o_val <= 16'b0101001011000101;
            14'h1ca7 	:	o_val <= 16'b0101001011000111;
            14'h1ca8 	:	o_val <= 16'b0101001011001010;
            14'h1ca9 	:	o_val <= 16'b0101001011001100;
            14'h1caa 	:	o_val <= 16'b0101001011001111;
            14'h1cab 	:	o_val <= 16'b0101001011010001;
            14'h1cac 	:	o_val <= 16'b0101001011010011;
            14'h1cad 	:	o_val <= 16'b0101001011010110;
            14'h1cae 	:	o_val <= 16'b0101001011011000;
            14'h1caf 	:	o_val <= 16'b0101001011011011;
            14'h1cb0 	:	o_val <= 16'b0101001011011101;
            14'h1cb1 	:	o_val <= 16'b0101001011011111;
            14'h1cb2 	:	o_val <= 16'b0101001011100010;
            14'h1cb3 	:	o_val <= 16'b0101001011100100;
            14'h1cb4 	:	o_val <= 16'b0101001011100111;
            14'h1cb5 	:	o_val <= 16'b0101001011101001;
            14'h1cb6 	:	o_val <= 16'b0101001011101011;
            14'h1cb7 	:	o_val <= 16'b0101001011101110;
            14'h1cb8 	:	o_val <= 16'b0101001011110000;
            14'h1cb9 	:	o_val <= 16'b0101001011110010;
            14'h1cba 	:	o_val <= 16'b0101001011110101;
            14'h1cbb 	:	o_val <= 16'b0101001011110111;
            14'h1cbc 	:	o_val <= 16'b0101001011111010;
            14'h1cbd 	:	o_val <= 16'b0101001011111100;
            14'h1cbe 	:	o_val <= 16'b0101001011111110;
            14'h1cbf 	:	o_val <= 16'b0101001100000001;
            14'h1cc0 	:	o_val <= 16'b0101001100000011;
            14'h1cc1 	:	o_val <= 16'b0101001100000110;
            14'h1cc2 	:	o_val <= 16'b0101001100001000;
            14'h1cc3 	:	o_val <= 16'b0101001100001010;
            14'h1cc4 	:	o_val <= 16'b0101001100001101;
            14'h1cc5 	:	o_val <= 16'b0101001100001111;
            14'h1cc6 	:	o_val <= 16'b0101001100010010;
            14'h1cc7 	:	o_val <= 16'b0101001100010100;
            14'h1cc8 	:	o_val <= 16'b0101001100010110;
            14'h1cc9 	:	o_val <= 16'b0101001100011001;
            14'h1cca 	:	o_val <= 16'b0101001100011011;
            14'h1ccb 	:	o_val <= 16'b0101001100011110;
            14'h1ccc 	:	o_val <= 16'b0101001100100000;
            14'h1ccd 	:	o_val <= 16'b0101001100100010;
            14'h1cce 	:	o_val <= 16'b0101001100100101;
            14'h1ccf 	:	o_val <= 16'b0101001100100111;
            14'h1cd0 	:	o_val <= 16'b0101001100101001;
            14'h1cd1 	:	o_val <= 16'b0101001100101100;
            14'h1cd2 	:	o_val <= 16'b0101001100101110;
            14'h1cd3 	:	o_val <= 16'b0101001100110001;
            14'h1cd4 	:	o_val <= 16'b0101001100110011;
            14'h1cd5 	:	o_val <= 16'b0101001100110101;
            14'h1cd6 	:	o_val <= 16'b0101001100111000;
            14'h1cd7 	:	o_val <= 16'b0101001100111010;
            14'h1cd8 	:	o_val <= 16'b0101001100111101;
            14'h1cd9 	:	o_val <= 16'b0101001100111111;
            14'h1cda 	:	o_val <= 16'b0101001101000001;
            14'h1cdb 	:	o_val <= 16'b0101001101000100;
            14'h1cdc 	:	o_val <= 16'b0101001101000110;
            14'h1cdd 	:	o_val <= 16'b0101001101001000;
            14'h1cde 	:	o_val <= 16'b0101001101001011;
            14'h1cdf 	:	o_val <= 16'b0101001101001101;
            14'h1ce0 	:	o_val <= 16'b0101001101010000;
            14'h1ce1 	:	o_val <= 16'b0101001101010010;
            14'h1ce2 	:	o_val <= 16'b0101001101010100;
            14'h1ce3 	:	o_val <= 16'b0101001101010111;
            14'h1ce4 	:	o_val <= 16'b0101001101011001;
            14'h1ce5 	:	o_val <= 16'b0101001101011100;
            14'h1ce6 	:	o_val <= 16'b0101001101011110;
            14'h1ce7 	:	o_val <= 16'b0101001101100000;
            14'h1ce8 	:	o_val <= 16'b0101001101100011;
            14'h1ce9 	:	o_val <= 16'b0101001101100101;
            14'h1cea 	:	o_val <= 16'b0101001101100111;
            14'h1ceb 	:	o_val <= 16'b0101001101101010;
            14'h1cec 	:	o_val <= 16'b0101001101101100;
            14'h1ced 	:	o_val <= 16'b0101001101101111;
            14'h1cee 	:	o_val <= 16'b0101001101110001;
            14'h1cef 	:	o_val <= 16'b0101001101110011;
            14'h1cf0 	:	o_val <= 16'b0101001101110110;
            14'h1cf1 	:	o_val <= 16'b0101001101111000;
            14'h1cf2 	:	o_val <= 16'b0101001101111011;
            14'h1cf3 	:	o_val <= 16'b0101001101111101;
            14'h1cf4 	:	o_val <= 16'b0101001101111111;
            14'h1cf5 	:	o_val <= 16'b0101001110000010;
            14'h1cf6 	:	o_val <= 16'b0101001110000100;
            14'h1cf7 	:	o_val <= 16'b0101001110000110;
            14'h1cf8 	:	o_val <= 16'b0101001110001001;
            14'h1cf9 	:	o_val <= 16'b0101001110001011;
            14'h1cfa 	:	o_val <= 16'b0101001110001110;
            14'h1cfb 	:	o_val <= 16'b0101001110010000;
            14'h1cfc 	:	o_val <= 16'b0101001110010010;
            14'h1cfd 	:	o_val <= 16'b0101001110010101;
            14'h1cfe 	:	o_val <= 16'b0101001110010111;
            14'h1cff 	:	o_val <= 16'b0101001110011001;
            14'h1d00 	:	o_val <= 16'b0101001110011100;
            14'h1d01 	:	o_val <= 16'b0101001110011110;
            14'h1d02 	:	o_val <= 16'b0101001110100001;
            14'h1d03 	:	o_val <= 16'b0101001110100011;
            14'h1d04 	:	o_val <= 16'b0101001110100101;
            14'h1d05 	:	o_val <= 16'b0101001110101000;
            14'h1d06 	:	o_val <= 16'b0101001110101010;
            14'h1d07 	:	o_val <= 16'b0101001110101101;
            14'h1d08 	:	o_val <= 16'b0101001110101111;
            14'h1d09 	:	o_val <= 16'b0101001110110001;
            14'h1d0a 	:	o_val <= 16'b0101001110110100;
            14'h1d0b 	:	o_val <= 16'b0101001110110110;
            14'h1d0c 	:	o_val <= 16'b0101001110111000;
            14'h1d0d 	:	o_val <= 16'b0101001110111011;
            14'h1d0e 	:	o_val <= 16'b0101001110111101;
            14'h1d0f 	:	o_val <= 16'b0101001111000000;
            14'h1d10 	:	o_val <= 16'b0101001111000010;
            14'h1d11 	:	o_val <= 16'b0101001111000100;
            14'h1d12 	:	o_val <= 16'b0101001111000111;
            14'h1d13 	:	o_val <= 16'b0101001111001001;
            14'h1d14 	:	o_val <= 16'b0101001111001011;
            14'h1d15 	:	o_val <= 16'b0101001111001110;
            14'h1d16 	:	o_val <= 16'b0101001111010000;
            14'h1d17 	:	o_val <= 16'b0101001111010011;
            14'h1d18 	:	o_val <= 16'b0101001111010101;
            14'h1d19 	:	o_val <= 16'b0101001111010111;
            14'h1d1a 	:	o_val <= 16'b0101001111011010;
            14'h1d1b 	:	o_val <= 16'b0101001111011100;
            14'h1d1c 	:	o_val <= 16'b0101001111011110;
            14'h1d1d 	:	o_val <= 16'b0101001111100001;
            14'h1d1e 	:	o_val <= 16'b0101001111100011;
            14'h1d1f 	:	o_val <= 16'b0101001111100110;
            14'h1d20 	:	o_val <= 16'b0101001111101000;
            14'h1d21 	:	o_val <= 16'b0101001111101010;
            14'h1d22 	:	o_val <= 16'b0101001111101101;
            14'h1d23 	:	o_val <= 16'b0101001111101111;
            14'h1d24 	:	o_val <= 16'b0101001111110001;
            14'h1d25 	:	o_val <= 16'b0101001111110100;
            14'h1d26 	:	o_val <= 16'b0101001111110110;
            14'h1d27 	:	o_val <= 16'b0101001111111000;
            14'h1d28 	:	o_val <= 16'b0101001111111011;
            14'h1d29 	:	o_val <= 16'b0101001111111101;
            14'h1d2a 	:	o_val <= 16'b0101010000000000;
            14'h1d2b 	:	o_val <= 16'b0101010000000010;
            14'h1d2c 	:	o_val <= 16'b0101010000000100;
            14'h1d2d 	:	o_val <= 16'b0101010000000111;
            14'h1d2e 	:	o_val <= 16'b0101010000001001;
            14'h1d2f 	:	o_val <= 16'b0101010000001011;
            14'h1d30 	:	o_val <= 16'b0101010000001110;
            14'h1d31 	:	o_val <= 16'b0101010000010000;
            14'h1d32 	:	o_val <= 16'b0101010000010011;
            14'h1d33 	:	o_val <= 16'b0101010000010101;
            14'h1d34 	:	o_val <= 16'b0101010000010111;
            14'h1d35 	:	o_val <= 16'b0101010000011010;
            14'h1d36 	:	o_val <= 16'b0101010000011100;
            14'h1d37 	:	o_val <= 16'b0101010000011110;
            14'h1d38 	:	o_val <= 16'b0101010000100001;
            14'h1d39 	:	o_val <= 16'b0101010000100011;
            14'h1d3a 	:	o_val <= 16'b0101010000100101;
            14'h1d3b 	:	o_val <= 16'b0101010000101000;
            14'h1d3c 	:	o_val <= 16'b0101010000101010;
            14'h1d3d 	:	o_val <= 16'b0101010000101101;
            14'h1d3e 	:	o_val <= 16'b0101010000101111;
            14'h1d3f 	:	o_val <= 16'b0101010000110001;
            14'h1d40 	:	o_val <= 16'b0101010000110100;
            14'h1d41 	:	o_val <= 16'b0101010000110110;
            14'h1d42 	:	o_val <= 16'b0101010000111000;
            14'h1d43 	:	o_val <= 16'b0101010000111011;
            14'h1d44 	:	o_val <= 16'b0101010000111101;
            14'h1d45 	:	o_val <= 16'b0101010001000000;
            14'h1d46 	:	o_val <= 16'b0101010001000010;
            14'h1d47 	:	o_val <= 16'b0101010001000100;
            14'h1d48 	:	o_val <= 16'b0101010001000111;
            14'h1d49 	:	o_val <= 16'b0101010001001001;
            14'h1d4a 	:	o_val <= 16'b0101010001001011;
            14'h1d4b 	:	o_val <= 16'b0101010001001110;
            14'h1d4c 	:	o_val <= 16'b0101010001010000;
            14'h1d4d 	:	o_val <= 16'b0101010001010010;
            14'h1d4e 	:	o_val <= 16'b0101010001010101;
            14'h1d4f 	:	o_val <= 16'b0101010001010111;
            14'h1d50 	:	o_val <= 16'b0101010001011010;
            14'h1d51 	:	o_val <= 16'b0101010001011100;
            14'h1d52 	:	o_val <= 16'b0101010001011110;
            14'h1d53 	:	o_val <= 16'b0101010001100001;
            14'h1d54 	:	o_val <= 16'b0101010001100011;
            14'h1d55 	:	o_val <= 16'b0101010001100101;
            14'h1d56 	:	o_val <= 16'b0101010001101000;
            14'h1d57 	:	o_val <= 16'b0101010001101010;
            14'h1d58 	:	o_val <= 16'b0101010001101100;
            14'h1d59 	:	o_val <= 16'b0101010001101111;
            14'h1d5a 	:	o_val <= 16'b0101010001110001;
            14'h1d5b 	:	o_val <= 16'b0101010001110100;
            14'h1d5c 	:	o_val <= 16'b0101010001110110;
            14'h1d5d 	:	o_val <= 16'b0101010001111000;
            14'h1d5e 	:	o_val <= 16'b0101010001111011;
            14'h1d5f 	:	o_val <= 16'b0101010001111101;
            14'h1d60 	:	o_val <= 16'b0101010001111111;
            14'h1d61 	:	o_val <= 16'b0101010010000010;
            14'h1d62 	:	o_val <= 16'b0101010010000100;
            14'h1d63 	:	o_val <= 16'b0101010010000110;
            14'h1d64 	:	o_val <= 16'b0101010010001001;
            14'h1d65 	:	o_val <= 16'b0101010010001011;
            14'h1d66 	:	o_val <= 16'b0101010010001101;
            14'h1d67 	:	o_val <= 16'b0101010010010000;
            14'h1d68 	:	o_val <= 16'b0101010010010010;
            14'h1d69 	:	o_val <= 16'b0101010010010101;
            14'h1d6a 	:	o_val <= 16'b0101010010010111;
            14'h1d6b 	:	o_val <= 16'b0101010010011001;
            14'h1d6c 	:	o_val <= 16'b0101010010011100;
            14'h1d6d 	:	o_val <= 16'b0101010010011110;
            14'h1d6e 	:	o_val <= 16'b0101010010100000;
            14'h1d6f 	:	o_val <= 16'b0101010010100011;
            14'h1d70 	:	o_val <= 16'b0101010010100101;
            14'h1d71 	:	o_val <= 16'b0101010010100111;
            14'h1d72 	:	o_val <= 16'b0101010010101010;
            14'h1d73 	:	o_val <= 16'b0101010010101100;
            14'h1d74 	:	o_val <= 16'b0101010010101110;
            14'h1d75 	:	o_val <= 16'b0101010010110001;
            14'h1d76 	:	o_val <= 16'b0101010010110011;
            14'h1d77 	:	o_val <= 16'b0101010010110110;
            14'h1d78 	:	o_val <= 16'b0101010010111000;
            14'h1d79 	:	o_val <= 16'b0101010010111010;
            14'h1d7a 	:	o_val <= 16'b0101010010111101;
            14'h1d7b 	:	o_val <= 16'b0101010010111111;
            14'h1d7c 	:	o_val <= 16'b0101010011000001;
            14'h1d7d 	:	o_val <= 16'b0101010011000100;
            14'h1d7e 	:	o_val <= 16'b0101010011000110;
            14'h1d7f 	:	o_val <= 16'b0101010011001000;
            14'h1d80 	:	o_val <= 16'b0101010011001011;
            14'h1d81 	:	o_val <= 16'b0101010011001101;
            14'h1d82 	:	o_val <= 16'b0101010011001111;
            14'h1d83 	:	o_val <= 16'b0101010011010010;
            14'h1d84 	:	o_val <= 16'b0101010011010100;
            14'h1d85 	:	o_val <= 16'b0101010011010110;
            14'h1d86 	:	o_val <= 16'b0101010011011001;
            14'h1d87 	:	o_val <= 16'b0101010011011011;
            14'h1d88 	:	o_val <= 16'b0101010011011110;
            14'h1d89 	:	o_val <= 16'b0101010011100000;
            14'h1d8a 	:	o_val <= 16'b0101010011100010;
            14'h1d8b 	:	o_val <= 16'b0101010011100101;
            14'h1d8c 	:	o_val <= 16'b0101010011100111;
            14'h1d8d 	:	o_val <= 16'b0101010011101001;
            14'h1d8e 	:	o_val <= 16'b0101010011101100;
            14'h1d8f 	:	o_val <= 16'b0101010011101110;
            14'h1d90 	:	o_val <= 16'b0101010011110000;
            14'h1d91 	:	o_val <= 16'b0101010011110011;
            14'h1d92 	:	o_val <= 16'b0101010011110101;
            14'h1d93 	:	o_val <= 16'b0101010011110111;
            14'h1d94 	:	o_val <= 16'b0101010011111010;
            14'h1d95 	:	o_val <= 16'b0101010011111100;
            14'h1d96 	:	o_val <= 16'b0101010011111110;
            14'h1d97 	:	o_val <= 16'b0101010100000001;
            14'h1d98 	:	o_val <= 16'b0101010100000011;
            14'h1d99 	:	o_val <= 16'b0101010100000101;
            14'h1d9a 	:	o_val <= 16'b0101010100001000;
            14'h1d9b 	:	o_val <= 16'b0101010100001010;
            14'h1d9c 	:	o_val <= 16'b0101010100001101;
            14'h1d9d 	:	o_val <= 16'b0101010100001111;
            14'h1d9e 	:	o_val <= 16'b0101010100010001;
            14'h1d9f 	:	o_val <= 16'b0101010100010100;
            14'h1da0 	:	o_val <= 16'b0101010100010110;
            14'h1da1 	:	o_val <= 16'b0101010100011000;
            14'h1da2 	:	o_val <= 16'b0101010100011011;
            14'h1da3 	:	o_val <= 16'b0101010100011101;
            14'h1da4 	:	o_val <= 16'b0101010100011111;
            14'h1da5 	:	o_val <= 16'b0101010100100010;
            14'h1da6 	:	o_val <= 16'b0101010100100100;
            14'h1da7 	:	o_val <= 16'b0101010100100110;
            14'h1da8 	:	o_val <= 16'b0101010100101001;
            14'h1da9 	:	o_val <= 16'b0101010100101011;
            14'h1daa 	:	o_val <= 16'b0101010100101101;
            14'h1dab 	:	o_val <= 16'b0101010100110000;
            14'h1dac 	:	o_val <= 16'b0101010100110010;
            14'h1dad 	:	o_val <= 16'b0101010100110100;
            14'h1dae 	:	o_val <= 16'b0101010100110111;
            14'h1daf 	:	o_val <= 16'b0101010100111001;
            14'h1db0 	:	o_val <= 16'b0101010100111011;
            14'h1db1 	:	o_val <= 16'b0101010100111110;
            14'h1db2 	:	o_val <= 16'b0101010101000000;
            14'h1db3 	:	o_val <= 16'b0101010101000010;
            14'h1db4 	:	o_val <= 16'b0101010101000101;
            14'h1db5 	:	o_val <= 16'b0101010101000111;
            14'h1db6 	:	o_val <= 16'b0101010101001010;
            14'h1db7 	:	o_val <= 16'b0101010101001100;
            14'h1db8 	:	o_val <= 16'b0101010101001110;
            14'h1db9 	:	o_val <= 16'b0101010101010001;
            14'h1dba 	:	o_val <= 16'b0101010101010011;
            14'h1dbb 	:	o_val <= 16'b0101010101010101;
            14'h1dbc 	:	o_val <= 16'b0101010101011000;
            14'h1dbd 	:	o_val <= 16'b0101010101011010;
            14'h1dbe 	:	o_val <= 16'b0101010101011100;
            14'h1dbf 	:	o_val <= 16'b0101010101011111;
            14'h1dc0 	:	o_val <= 16'b0101010101100001;
            14'h1dc1 	:	o_val <= 16'b0101010101100011;
            14'h1dc2 	:	o_val <= 16'b0101010101100110;
            14'h1dc3 	:	o_val <= 16'b0101010101101000;
            14'h1dc4 	:	o_val <= 16'b0101010101101010;
            14'h1dc5 	:	o_val <= 16'b0101010101101101;
            14'h1dc6 	:	o_val <= 16'b0101010101101111;
            14'h1dc7 	:	o_val <= 16'b0101010101110001;
            14'h1dc8 	:	o_val <= 16'b0101010101110100;
            14'h1dc9 	:	o_val <= 16'b0101010101110110;
            14'h1dca 	:	o_val <= 16'b0101010101111000;
            14'h1dcb 	:	o_val <= 16'b0101010101111011;
            14'h1dcc 	:	o_val <= 16'b0101010101111101;
            14'h1dcd 	:	o_val <= 16'b0101010101111111;
            14'h1dce 	:	o_val <= 16'b0101010110000010;
            14'h1dcf 	:	o_val <= 16'b0101010110000100;
            14'h1dd0 	:	o_val <= 16'b0101010110000110;
            14'h1dd1 	:	o_val <= 16'b0101010110001001;
            14'h1dd2 	:	o_val <= 16'b0101010110001011;
            14'h1dd3 	:	o_val <= 16'b0101010110001101;
            14'h1dd4 	:	o_val <= 16'b0101010110010000;
            14'h1dd5 	:	o_val <= 16'b0101010110010010;
            14'h1dd6 	:	o_val <= 16'b0101010110010100;
            14'h1dd7 	:	o_val <= 16'b0101010110010111;
            14'h1dd8 	:	o_val <= 16'b0101010110011001;
            14'h1dd9 	:	o_val <= 16'b0101010110011011;
            14'h1dda 	:	o_val <= 16'b0101010110011110;
            14'h1ddb 	:	o_val <= 16'b0101010110100000;
            14'h1ddc 	:	o_val <= 16'b0101010110100010;
            14'h1ddd 	:	o_val <= 16'b0101010110100101;
            14'h1dde 	:	o_val <= 16'b0101010110100111;
            14'h1ddf 	:	o_val <= 16'b0101010110101001;
            14'h1de0 	:	o_val <= 16'b0101010110101100;
            14'h1de1 	:	o_val <= 16'b0101010110101110;
            14'h1de2 	:	o_val <= 16'b0101010110110000;
            14'h1de3 	:	o_val <= 16'b0101010110110011;
            14'h1de4 	:	o_val <= 16'b0101010110110101;
            14'h1de5 	:	o_val <= 16'b0101010110110111;
            14'h1de6 	:	o_val <= 16'b0101010110111010;
            14'h1de7 	:	o_val <= 16'b0101010110111100;
            14'h1de8 	:	o_val <= 16'b0101010110111110;
            14'h1de9 	:	o_val <= 16'b0101010111000001;
            14'h1dea 	:	o_val <= 16'b0101010111000011;
            14'h1deb 	:	o_val <= 16'b0101010111000101;
            14'h1dec 	:	o_val <= 16'b0101010111001000;
            14'h1ded 	:	o_val <= 16'b0101010111001010;
            14'h1dee 	:	o_val <= 16'b0101010111001100;
            14'h1def 	:	o_val <= 16'b0101010111001111;
            14'h1df0 	:	o_val <= 16'b0101010111010001;
            14'h1df1 	:	o_val <= 16'b0101010111010011;
            14'h1df2 	:	o_val <= 16'b0101010111010110;
            14'h1df3 	:	o_val <= 16'b0101010111011000;
            14'h1df4 	:	o_val <= 16'b0101010111011010;
            14'h1df5 	:	o_val <= 16'b0101010111011101;
            14'h1df6 	:	o_val <= 16'b0101010111011111;
            14'h1df7 	:	o_val <= 16'b0101010111100001;
            14'h1df8 	:	o_val <= 16'b0101010111100100;
            14'h1df9 	:	o_val <= 16'b0101010111100110;
            14'h1dfa 	:	o_val <= 16'b0101010111101000;
            14'h1dfb 	:	o_val <= 16'b0101010111101011;
            14'h1dfc 	:	o_val <= 16'b0101010111101101;
            14'h1dfd 	:	o_val <= 16'b0101010111101111;
            14'h1dfe 	:	o_val <= 16'b0101010111110010;
            14'h1dff 	:	o_val <= 16'b0101010111110100;
            14'h1e00 	:	o_val <= 16'b0101010111110110;
            14'h1e01 	:	o_val <= 16'b0101010111111001;
            14'h1e02 	:	o_val <= 16'b0101010111111011;
            14'h1e03 	:	o_val <= 16'b0101010111111101;
            14'h1e04 	:	o_val <= 16'b0101011000000000;
            14'h1e05 	:	o_val <= 16'b0101011000000010;
            14'h1e06 	:	o_val <= 16'b0101011000000100;
            14'h1e07 	:	o_val <= 16'b0101011000000111;
            14'h1e08 	:	o_val <= 16'b0101011000001001;
            14'h1e09 	:	o_val <= 16'b0101011000001011;
            14'h1e0a 	:	o_val <= 16'b0101011000001110;
            14'h1e0b 	:	o_val <= 16'b0101011000010000;
            14'h1e0c 	:	o_val <= 16'b0101011000010010;
            14'h1e0d 	:	o_val <= 16'b0101011000010101;
            14'h1e0e 	:	o_val <= 16'b0101011000010111;
            14'h1e0f 	:	o_val <= 16'b0101011000011001;
            14'h1e10 	:	o_val <= 16'b0101011000011100;
            14'h1e11 	:	o_val <= 16'b0101011000011110;
            14'h1e12 	:	o_val <= 16'b0101011000100000;
            14'h1e13 	:	o_val <= 16'b0101011000100010;
            14'h1e14 	:	o_val <= 16'b0101011000100101;
            14'h1e15 	:	o_val <= 16'b0101011000100111;
            14'h1e16 	:	o_val <= 16'b0101011000101001;
            14'h1e17 	:	o_val <= 16'b0101011000101100;
            14'h1e18 	:	o_val <= 16'b0101011000101110;
            14'h1e19 	:	o_val <= 16'b0101011000110000;
            14'h1e1a 	:	o_val <= 16'b0101011000110011;
            14'h1e1b 	:	o_val <= 16'b0101011000110101;
            14'h1e1c 	:	o_val <= 16'b0101011000110111;
            14'h1e1d 	:	o_val <= 16'b0101011000111010;
            14'h1e1e 	:	o_val <= 16'b0101011000111100;
            14'h1e1f 	:	o_val <= 16'b0101011000111110;
            14'h1e20 	:	o_val <= 16'b0101011001000001;
            14'h1e21 	:	o_val <= 16'b0101011001000011;
            14'h1e22 	:	o_val <= 16'b0101011001000101;
            14'h1e23 	:	o_val <= 16'b0101011001001000;
            14'h1e24 	:	o_val <= 16'b0101011001001010;
            14'h1e25 	:	o_val <= 16'b0101011001001100;
            14'h1e26 	:	o_val <= 16'b0101011001001111;
            14'h1e27 	:	o_val <= 16'b0101011001010001;
            14'h1e28 	:	o_val <= 16'b0101011001010011;
            14'h1e29 	:	o_val <= 16'b0101011001010110;
            14'h1e2a 	:	o_val <= 16'b0101011001011000;
            14'h1e2b 	:	o_val <= 16'b0101011001011010;
            14'h1e2c 	:	o_val <= 16'b0101011001011101;
            14'h1e2d 	:	o_val <= 16'b0101011001011111;
            14'h1e2e 	:	o_val <= 16'b0101011001100001;
            14'h1e2f 	:	o_val <= 16'b0101011001100011;
            14'h1e30 	:	o_val <= 16'b0101011001100110;
            14'h1e31 	:	o_val <= 16'b0101011001101000;
            14'h1e32 	:	o_val <= 16'b0101011001101010;
            14'h1e33 	:	o_val <= 16'b0101011001101101;
            14'h1e34 	:	o_val <= 16'b0101011001101111;
            14'h1e35 	:	o_val <= 16'b0101011001110001;
            14'h1e36 	:	o_val <= 16'b0101011001110100;
            14'h1e37 	:	o_val <= 16'b0101011001110110;
            14'h1e38 	:	o_val <= 16'b0101011001111000;
            14'h1e39 	:	o_val <= 16'b0101011001111011;
            14'h1e3a 	:	o_val <= 16'b0101011001111101;
            14'h1e3b 	:	o_val <= 16'b0101011001111111;
            14'h1e3c 	:	o_val <= 16'b0101011010000010;
            14'h1e3d 	:	o_val <= 16'b0101011010000100;
            14'h1e3e 	:	o_val <= 16'b0101011010000110;
            14'h1e3f 	:	o_val <= 16'b0101011010001001;
            14'h1e40 	:	o_val <= 16'b0101011010001011;
            14'h1e41 	:	o_val <= 16'b0101011010001101;
            14'h1e42 	:	o_val <= 16'b0101011010001111;
            14'h1e43 	:	o_val <= 16'b0101011010010010;
            14'h1e44 	:	o_val <= 16'b0101011010010100;
            14'h1e45 	:	o_val <= 16'b0101011010010110;
            14'h1e46 	:	o_val <= 16'b0101011010011001;
            14'h1e47 	:	o_val <= 16'b0101011010011011;
            14'h1e48 	:	o_val <= 16'b0101011010011101;
            14'h1e49 	:	o_val <= 16'b0101011010100000;
            14'h1e4a 	:	o_val <= 16'b0101011010100010;
            14'h1e4b 	:	o_val <= 16'b0101011010100100;
            14'h1e4c 	:	o_val <= 16'b0101011010100111;
            14'h1e4d 	:	o_val <= 16'b0101011010101001;
            14'h1e4e 	:	o_val <= 16'b0101011010101011;
            14'h1e4f 	:	o_val <= 16'b0101011010101110;
            14'h1e50 	:	o_val <= 16'b0101011010110000;
            14'h1e51 	:	o_val <= 16'b0101011010110010;
            14'h1e52 	:	o_val <= 16'b0101011010110100;
            14'h1e53 	:	o_val <= 16'b0101011010110111;
            14'h1e54 	:	o_val <= 16'b0101011010111001;
            14'h1e55 	:	o_val <= 16'b0101011010111011;
            14'h1e56 	:	o_val <= 16'b0101011010111110;
            14'h1e57 	:	o_val <= 16'b0101011011000000;
            14'h1e58 	:	o_val <= 16'b0101011011000010;
            14'h1e59 	:	o_val <= 16'b0101011011000101;
            14'h1e5a 	:	o_val <= 16'b0101011011000111;
            14'h1e5b 	:	o_val <= 16'b0101011011001001;
            14'h1e5c 	:	o_val <= 16'b0101011011001100;
            14'h1e5d 	:	o_val <= 16'b0101011011001110;
            14'h1e5e 	:	o_val <= 16'b0101011011010000;
            14'h1e5f 	:	o_val <= 16'b0101011011010011;
            14'h1e60 	:	o_val <= 16'b0101011011010101;
            14'h1e61 	:	o_val <= 16'b0101011011010111;
            14'h1e62 	:	o_val <= 16'b0101011011011001;
            14'h1e63 	:	o_val <= 16'b0101011011011100;
            14'h1e64 	:	o_val <= 16'b0101011011011110;
            14'h1e65 	:	o_val <= 16'b0101011011100000;
            14'h1e66 	:	o_val <= 16'b0101011011100011;
            14'h1e67 	:	o_val <= 16'b0101011011100101;
            14'h1e68 	:	o_val <= 16'b0101011011100111;
            14'h1e69 	:	o_val <= 16'b0101011011101010;
            14'h1e6a 	:	o_val <= 16'b0101011011101100;
            14'h1e6b 	:	o_val <= 16'b0101011011101110;
            14'h1e6c 	:	o_val <= 16'b0101011011110001;
            14'h1e6d 	:	o_val <= 16'b0101011011110011;
            14'h1e6e 	:	o_val <= 16'b0101011011110101;
            14'h1e6f 	:	o_val <= 16'b0101011011110111;
            14'h1e70 	:	o_val <= 16'b0101011011111010;
            14'h1e71 	:	o_val <= 16'b0101011011111100;
            14'h1e72 	:	o_val <= 16'b0101011011111110;
            14'h1e73 	:	o_val <= 16'b0101011100000001;
            14'h1e74 	:	o_val <= 16'b0101011100000011;
            14'h1e75 	:	o_val <= 16'b0101011100000101;
            14'h1e76 	:	o_val <= 16'b0101011100001000;
            14'h1e77 	:	o_val <= 16'b0101011100001010;
            14'h1e78 	:	o_val <= 16'b0101011100001100;
            14'h1e79 	:	o_val <= 16'b0101011100001110;
            14'h1e7a 	:	o_val <= 16'b0101011100010001;
            14'h1e7b 	:	o_val <= 16'b0101011100010011;
            14'h1e7c 	:	o_val <= 16'b0101011100010101;
            14'h1e7d 	:	o_val <= 16'b0101011100011000;
            14'h1e7e 	:	o_val <= 16'b0101011100011010;
            14'h1e7f 	:	o_val <= 16'b0101011100011100;
            14'h1e80 	:	o_val <= 16'b0101011100011111;
            14'h1e81 	:	o_val <= 16'b0101011100100001;
            14'h1e82 	:	o_val <= 16'b0101011100100011;
            14'h1e83 	:	o_val <= 16'b0101011100100101;
            14'h1e84 	:	o_val <= 16'b0101011100101000;
            14'h1e85 	:	o_val <= 16'b0101011100101010;
            14'h1e86 	:	o_val <= 16'b0101011100101100;
            14'h1e87 	:	o_val <= 16'b0101011100101111;
            14'h1e88 	:	o_val <= 16'b0101011100110001;
            14'h1e89 	:	o_val <= 16'b0101011100110011;
            14'h1e8a 	:	o_val <= 16'b0101011100110110;
            14'h1e8b 	:	o_val <= 16'b0101011100111000;
            14'h1e8c 	:	o_val <= 16'b0101011100111010;
            14'h1e8d 	:	o_val <= 16'b0101011100111100;
            14'h1e8e 	:	o_val <= 16'b0101011100111111;
            14'h1e8f 	:	o_val <= 16'b0101011101000001;
            14'h1e90 	:	o_val <= 16'b0101011101000011;
            14'h1e91 	:	o_val <= 16'b0101011101000110;
            14'h1e92 	:	o_val <= 16'b0101011101001000;
            14'h1e93 	:	o_val <= 16'b0101011101001010;
            14'h1e94 	:	o_val <= 16'b0101011101001101;
            14'h1e95 	:	o_val <= 16'b0101011101001111;
            14'h1e96 	:	o_val <= 16'b0101011101010001;
            14'h1e97 	:	o_val <= 16'b0101011101010011;
            14'h1e98 	:	o_val <= 16'b0101011101010110;
            14'h1e99 	:	o_val <= 16'b0101011101011000;
            14'h1e9a 	:	o_val <= 16'b0101011101011010;
            14'h1e9b 	:	o_val <= 16'b0101011101011101;
            14'h1e9c 	:	o_val <= 16'b0101011101011111;
            14'h1e9d 	:	o_val <= 16'b0101011101100001;
            14'h1e9e 	:	o_val <= 16'b0101011101100100;
            14'h1e9f 	:	o_val <= 16'b0101011101100110;
            14'h1ea0 	:	o_val <= 16'b0101011101101000;
            14'h1ea1 	:	o_val <= 16'b0101011101101010;
            14'h1ea2 	:	o_val <= 16'b0101011101101101;
            14'h1ea3 	:	o_val <= 16'b0101011101101111;
            14'h1ea4 	:	o_val <= 16'b0101011101110001;
            14'h1ea5 	:	o_val <= 16'b0101011101110100;
            14'h1ea6 	:	o_val <= 16'b0101011101110110;
            14'h1ea7 	:	o_val <= 16'b0101011101111000;
            14'h1ea8 	:	o_val <= 16'b0101011101111010;
            14'h1ea9 	:	o_val <= 16'b0101011101111101;
            14'h1eaa 	:	o_val <= 16'b0101011101111111;
            14'h1eab 	:	o_val <= 16'b0101011110000001;
            14'h1eac 	:	o_val <= 16'b0101011110000100;
            14'h1ead 	:	o_val <= 16'b0101011110000110;
            14'h1eae 	:	o_val <= 16'b0101011110001000;
            14'h1eaf 	:	o_val <= 16'b0101011110001011;
            14'h1eb0 	:	o_val <= 16'b0101011110001101;
            14'h1eb1 	:	o_val <= 16'b0101011110001111;
            14'h1eb2 	:	o_val <= 16'b0101011110010001;
            14'h1eb3 	:	o_val <= 16'b0101011110010100;
            14'h1eb4 	:	o_val <= 16'b0101011110010110;
            14'h1eb5 	:	o_val <= 16'b0101011110011000;
            14'h1eb6 	:	o_val <= 16'b0101011110011011;
            14'h1eb7 	:	o_val <= 16'b0101011110011101;
            14'h1eb8 	:	o_val <= 16'b0101011110011111;
            14'h1eb9 	:	o_val <= 16'b0101011110100001;
            14'h1eba 	:	o_val <= 16'b0101011110100100;
            14'h1ebb 	:	o_val <= 16'b0101011110100110;
            14'h1ebc 	:	o_val <= 16'b0101011110101000;
            14'h1ebd 	:	o_val <= 16'b0101011110101011;
            14'h1ebe 	:	o_val <= 16'b0101011110101101;
            14'h1ebf 	:	o_val <= 16'b0101011110101111;
            14'h1ec0 	:	o_val <= 16'b0101011110110001;
            14'h1ec1 	:	o_val <= 16'b0101011110110100;
            14'h1ec2 	:	o_val <= 16'b0101011110110110;
            14'h1ec3 	:	o_val <= 16'b0101011110111000;
            14'h1ec4 	:	o_val <= 16'b0101011110111011;
            14'h1ec5 	:	o_val <= 16'b0101011110111101;
            14'h1ec6 	:	o_val <= 16'b0101011110111111;
            14'h1ec7 	:	o_val <= 16'b0101011111000001;
            14'h1ec8 	:	o_val <= 16'b0101011111000100;
            14'h1ec9 	:	o_val <= 16'b0101011111000110;
            14'h1eca 	:	o_val <= 16'b0101011111001000;
            14'h1ecb 	:	o_val <= 16'b0101011111001011;
            14'h1ecc 	:	o_val <= 16'b0101011111001101;
            14'h1ecd 	:	o_val <= 16'b0101011111001111;
            14'h1ece 	:	o_val <= 16'b0101011111010001;
            14'h1ecf 	:	o_val <= 16'b0101011111010100;
            14'h1ed0 	:	o_val <= 16'b0101011111010110;
            14'h1ed1 	:	o_val <= 16'b0101011111011000;
            14'h1ed2 	:	o_val <= 16'b0101011111011011;
            14'h1ed3 	:	o_val <= 16'b0101011111011101;
            14'h1ed4 	:	o_val <= 16'b0101011111011111;
            14'h1ed5 	:	o_val <= 16'b0101011111100001;
            14'h1ed6 	:	o_val <= 16'b0101011111100100;
            14'h1ed7 	:	o_val <= 16'b0101011111100110;
            14'h1ed8 	:	o_val <= 16'b0101011111101000;
            14'h1ed9 	:	o_val <= 16'b0101011111101011;
            14'h1eda 	:	o_val <= 16'b0101011111101101;
            14'h1edb 	:	o_val <= 16'b0101011111101111;
            14'h1edc 	:	o_val <= 16'b0101011111110001;
            14'h1edd 	:	o_val <= 16'b0101011111110100;
            14'h1ede 	:	o_val <= 16'b0101011111110110;
            14'h1edf 	:	o_val <= 16'b0101011111111000;
            14'h1ee0 	:	o_val <= 16'b0101011111111011;
            14'h1ee1 	:	o_val <= 16'b0101011111111101;
            14'h1ee2 	:	o_val <= 16'b0101011111111111;
            14'h1ee3 	:	o_val <= 16'b0101100000000001;
            14'h1ee4 	:	o_val <= 16'b0101100000000100;
            14'h1ee5 	:	o_val <= 16'b0101100000000110;
            14'h1ee6 	:	o_val <= 16'b0101100000001000;
            14'h1ee7 	:	o_val <= 16'b0101100000001011;
            14'h1ee8 	:	o_val <= 16'b0101100000001101;
            14'h1ee9 	:	o_val <= 16'b0101100000001111;
            14'h1eea 	:	o_val <= 16'b0101100000010001;
            14'h1eeb 	:	o_val <= 16'b0101100000010100;
            14'h1eec 	:	o_val <= 16'b0101100000010110;
            14'h1eed 	:	o_val <= 16'b0101100000011000;
            14'h1eee 	:	o_val <= 16'b0101100000011011;
            14'h1eef 	:	o_val <= 16'b0101100000011101;
            14'h1ef0 	:	o_val <= 16'b0101100000011111;
            14'h1ef1 	:	o_val <= 16'b0101100000100001;
            14'h1ef2 	:	o_val <= 16'b0101100000100100;
            14'h1ef3 	:	o_val <= 16'b0101100000100110;
            14'h1ef4 	:	o_val <= 16'b0101100000101000;
            14'h1ef5 	:	o_val <= 16'b0101100000101010;
            14'h1ef6 	:	o_val <= 16'b0101100000101101;
            14'h1ef7 	:	o_val <= 16'b0101100000101111;
            14'h1ef8 	:	o_val <= 16'b0101100000110001;
            14'h1ef9 	:	o_val <= 16'b0101100000110100;
            14'h1efa 	:	o_val <= 16'b0101100000110110;
            14'h1efb 	:	o_val <= 16'b0101100000111000;
            14'h1efc 	:	o_val <= 16'b0101100000111010;
            14'h1efd 	:	o_val <= 16'b0101100000111101;
            14'h1efe 	:	o_val <= 16'b0101100000111111;
            14'h1eff 	:	o_val <= 16'b0101100001000001;
            14'h1f00 	:	o_val <= 16'b0101100001000100;
            14'h1f01 	:	o_val <= 16'b0101100001000110;
            14'h1f02 	:	o_val <= 16'b0101100001001000;
            14'h1f03 	:	o_val <= 16'b0101100001001010;
            14'h1f04 	:	o_val <= 16'b0101100001001101;
            14'h1f05 	:	o_val <= 16'b0101100001001111;
            14'h1f06 	:	o_val <= 16'b0101100001010001;
            14'h1f07 	:	o_val <= 16'b0101100001010011;
            14'h1f08 	:	o_val <= 16'b0101100001010110;
            14'h1f09 	:	o_val <= 16'b0101100001011000;
            14'h1f0a 	:	o_val <= 16'b0101100001011010;
            14'h1f0b 	:	o_val <= 16'b0101100001011101;
            14'h1f0c 	:	o_val <= 16'b0101100001011111;
            14'h1f0d 	:	o_val <= 16'b0101100001100001;
            14'h1f0e 	:	o_val <= 16'b0101100001100011;
            14'h1f0f 	:	o_val <= 16'b0101100001100110;
            14'h1f10 	:	o_val <= 16'b0101100001101000;
            14'h1f11 	:	o_val <= 16'b0101100001101010;
            14'h1f12 	:	o_val <= 16'b0101100001101100;
            14'h1f13 	:	o_val <= 16'b0101100001101111;
            14'h1f14 	:	o_val <= 16'b0101100001110001;
            14'h1f15 	:	o_val <= 16'b0101100001110011;
            14'h1f16 	:	o_val <= 16'b0101100001110110;
            14'h1f17 	:	o_val <= 16'b0101100001111000;
            14'h1f18 	:	o_val <= 16'b0101100001111010;
            14'h1f19 	:	o_val <= 16'b0101100001111100;
            14'h1f1a 	:	o_val <= 16'b0101100001111111;
            14'h1f1b 	:	o_val <= 16'b0101100010000001;
            14'h1f1c 	:	o_val <= 16'b0101100010000011;
            14'h1f1d 	:	o_val <= 16'b0101100010000101;
            14'h1f1e 	:	o_val <= 16'b0101100010001000;
            14'h1f1f 	:	o_val <= 16'b0101100010001010;
            14'h1f20 	:	o_val <= 16'b0101100010001100;
            14'h1f21 	:	o_val <= 16'b0101100010001110;
            14'h1f22 	:	o_val <= 16'b0101100010010001;
            14'h1f23 	:	o_val <= 16'b0101100010010011;
            14'h1f24 	:	o_val <= 16'b0101100010010101;
            14'h1f25 	:	o_val <= 16'b0101100010011000;
            14'h1f26 	:	o_val <= 16'b0101100010011010;
            14'h1f27 	:	o_val <= 16'b0101100010011100;
            14'h1f28 	:	o_val <= 16'b0101100010011110;
            14'h1f29 	:	o_val <= 16'b0101100010100001;
            14'h1f2a 	:	o_val <= 16'b0101100010100011;
            14'h1f2b 	:	o_val <= 16'b0101100010100101;
            14'h1f2c 	:	o_val <= 16'b0101100010100111;
            14'h1f2d 	:	o_val <= 16'b0101100010101010;
            14'h1f2e 	:	o_val <= 16'b0101100010101100;
            14'h1f2f 	:	o_val <= 16'b0101100010101110;
            14'h1f30 	:	o_val <= 16'b0101100010110000;
            14'h1f31 	:	o_val <= 16'b0101100010110011;
            14'h1f32 	:	o_val <= 16'b0101100010110101;
            14'h1f33 	:	o_val <= 16'b0101100010110111;
            14'h1f34 	:	o_val <= 16'b0101100010111010;
            14'h1f35 	:	o_val <= 16'b0101100010111100;
            14'h1f36 	:	o_val <= 16'b0101100010111110;
            14'h1f37 	:	o_val <= 16'b0101100011000000;
            14'h1f38 	:	o_val <= 16'b0101100011000011;
            14'h1f39 	:	o_val <= 16'b0101100011000101;
            14'h1f3a 	:	o_val <= 16'b0101100011000111;
            14'h1f3b 	:	o_val <= 16'b0101100011001001;
            14'h1f3c 	:	o_val <= 16'b0101100011001100;
            14'h1f3d 	:	o_val <= 16'b0101100011001110;
            14'h1f3e 	:	o_val <= 16'b0101100011010000;
            14'h1f3f 	:	o_val <= 16'b0101100011010010;
            14'h1f40 	:	o_val <= 16'b0101100011010101;
            14'h1f41 	:	o_val <= 16'b0101100011010111;
            14'h1f42 	:	o_val <= 16'b0101100011011001;
            14'h1f43 	:	o_val <= 16'b0101100011011011;
            14'h1f44 	:	o_val <= 16'b0101100011011110;
            14'h1f45 	:	o_val <= 16'b0101100011100000;
            14'h1f46 	:	o_val <= 16'b0101100011100010;
            14'h1f47 	:	o_val <= 16'b0101100011100101;
            14'h1f48 	:	o_val <= 16'b0101100011100111;
            14'h1f49 	:	o_val <= 16'b0101100011101001;
            14'h1f4a 	:	o_val <= 16'b0101100011101011;
            14'h1f4b 	:	o_val <= 16'b0101100011101110;
            14'h1f4c 	:	o_val <= 16'b0101100011110000;
            14'h1f4d 	:	o_val <= 16'b0101100011110010;
            14'h1f4e 	:	o_val <= 16'b0101100011110100;
            14'h1f4f 	:	o_val <= 16'b0101100011110111;
            14'h1f50 	:	o_val <= 16'b0101100011111001;
            14'h1f51 	:	o_val <= 16'b0101100011111011;
            14'h1f52 	:	o_val <= 16'b0101100011111101;
            14'h1f53 	:	o_val <= 16'b0101100100000000;
            14'h1f54 	:	o_val <= 16'b0101100100000010;
            14'h1f55 	:	o_val <= 16'b0101100100000100;
            14'h1f56 	:	o_val <= 16'b0101100100000110;
            14'h1f57 	:	o_val <= 16'b0101100100001001;
            14'h1f58 	:	o_val <= 16'b0101100100001011;
            14'h1f59 	:	o_val <= 16'b0101100100001101;
            14'h1f5a 	:	o_val <= 16'b0101100100001111;
            14'h1f5b 	:	o_val <= 16'b0101100100010010;
            14'h1f5c 	:	o_val <= 16'b0101100100010100;
            14'h1f5d 	:	o_val <= 16'b0101100100010110;
            14'h1f5e 	:	o_val <= 16'b0101100100011000;
            14'h1f5f 	:	o_val <= 16'b0101100100011011;
            14'h1f60 	:	o_val <= 16'b0101100100011101;
            14'h1f61 	:	o_val <= 16'b0101100100011111;
            14'h1f62 	:	o_val <= 16'b0101100100100001;
            14'h1f63 	:	o_val <= 16'b0101100100100100;
            14'h1f64 	:	o_val <= 16'b0101100100100110;
            14'h1f65 	:	o_val <= 16'b0101100100101000;
            14'h1f66 	:	o_val <= 16'b0101100100101010;
            14'h1f67 	:	o_val <= 16'b0101100100101101;
            14'h1f68 	:	o_val <= 16'b0101100100101111;
            14'h1f69 	:	o_val <= 16'b0101100100110001;
            14'h1f6a 	:	o_val <= 16'b0101100100110100;
            14'h1f6b 	:	o_val <= 16'b0101100100110110;
            14'h1f6c 	:	o_val <= 16'b0101100100111000;
            14'h1f6d 	:	o_val <= 16'b0101100100111010;
            14'h1f6e 	:	o_val <= 16'b0101100100111101;
            14'h1f6f 	:	o_val <= 16'b0101100100111111;
            14'h1f70 	:	o_val <= 16'b0101100101000001;
            14'h1f71 	:	o_val <= 16'b0101100101000011;
            14'h1f72 	:	o_val <= 16'b0101100101000110;
            14'h1f73 	:	o_val <= 16'b0101100101001000;
            14'h1f74 	:	o_val <= 16'b0101100101001010;
            14'h1f75 	:	o_val <= 16'b0101100101001100;
            14'h1f76 	:	o_val <= 16'b0101100101001111;
            14'h1f77 	:	o_val <= 16'b0101100101010001;
            14'h1f78 	:	o_val <= 16'b0101100101010011;
            14'h1f79 	:	o_val <= 16'b0101100101010101;
            14'h1f7a 	:	o_val <= 16'b0101100101011000;
            14'h1f7b 	:	o_val <= 16'b0101100101011010;
            14'h1f7c 	:	o_val <= 16'b0101100101011100;
            14'h1f7d 	:	o_val <= 16'b0101100101011110;
            14'h1f7e 	:	o_val <= 16'b0101100101100001;
            14'h1f7f 	:	o_val <= 16'b0101100101100011;
            14'h1f80 	:	o_val <= 16'b0101100101100101;
            14'h1f81 	:	o_val <= 16'b0101100101100111;
            14'h1f82 	:	o_val <= 16'b0101100101101010;
            14'h1f83 	:	o_val <= 16'b0101100101101100;
            14'h1f84 	:	o_val <= 16'b0101100101101110;
            14'h1f85 	:	o_val <= 16'b0101100101110000;
            14'h1f86 	:	o_val <= 16'b0101100101110011;
            14'h1f87 	:	o_val <= 16'b0101100101110101;
            14'h1f88 	:	o_val <= 16'b0101100101110111;
            14'h1f89 	:	o_val <= 16'b0101100101111001;
            14'h1f8a 	:	o_val <= 16'b0101100101111011;
            14'h1f8b 	:	o_val <= 16'b0101100101111110;
            14'h1f8c 	:	o_val <= 16'b0101100110000000;
            14'h1f8d 	:	o_val <= 16'b0101100110000010;
            14'h1f8e 	:	o_val <= 16'b0101100110000100;
            14'h1f8f 	:	o_val <= 16'b0101100110000111;
            14'h1f90 	:	o_val <= 16'b0101100110001001;
            14'h1f91 	:	o_val <= 16'b0101100110001011;
            14'h1f92 	:	o_val <= 16'b0101100110001101;
            14'h1f93 	:	o_val <= 16'b0101100110010000;
            14'h1f94 	:	o_val <= 16'b0101100110010010;
            14'h1f95 	:	o_val <= 16'b0101100110010100;
            14'h1f96 	:	o_val <= 16'b0101100110010110;
            14'h1f97 	:	o_val <= 16'b0101100110011001;
            14'h1f98 	:	o_val <= 16'b0101100110011011;
            14'h1f99 	:	o_val <= 16'b0101100110011101;
            14'h1f9a 	:	o_val <= 16'b0101100110011111;
            14'h1f9b 	:	o_val <= 16'b0101100110100010;
            14'h1f9c 	:	o_val <= 16'b0101100110100100;
            14'h1f9d 	:	o_val <= 16'b0101100110100110;
            14'h1f9e 	:	o_val <= 16'b0101100110101000;
            14'h1f9f 	:	o_val <= 16'b0101100110101011;
            14'h1fa0 	:	o_val <= 16'b0101100110101101;
            14'h1fa1 	:	o_val <= 16'b0101100110101111;
            14'h1fa2 	:	o_val <= 16'b0101100110110001;
            14'h1fa3 	:	o_val <= 16'b0101100110110100;
            14'h1fa4 	:	o_val <= 16'b0101100110110110;
            14'h1fa5 	:	o_val <= 16'b0101100110111000;
            14'h1fa6 	:	o_val <= 16'b0101100110111010;
            14'h1fa7 	:	o_val <= 16'b0101100110111101;
            14'h1fa8 	:	o_val <= 16'b0101100110111111;
            14'h1fa9 	:	o_val <= 16'b0101100111000001;
            14'h1faa 	:	o_val <= 16'b0101100111000011;
            14'h1fab 	:	o_val <= 16'b0101100111000110;
            14'h1fac 	:	o_val <= 16'b0101100111001000;
            14'h1fad 	:	o_val <= 16'b0101100111001010;
            14'h1fae 	:	o_val <= 16'b0101100111001100;
            14'h1faf 	:	o_val <= 16'b0101100111001110;
            14'h1fb0 	:	o_val <= 16'b0101100111010001;
            14'h1fb1 	:	o_val <= 16'b0101100111010011;
            14'h1fb2 	:	o_val <= 16'b0101100111010101;
            14'h1fb3 	:	o_val <= 16'b0101100111010111;
            14'h1fb4 	:	o_val <= 16'b0101100111011010;
            14'h1fb5 	:	o_val <= 16'b0101100111011100;
            14'h1fb6 	:	o_val <= 16'b0101100111011110;
            14'h1fb7 	:	o_val <= 16'b0101100111100000;
            14'h1fb8 	:	o_val <= 16'b0101100111100011;
            14'h1fb9 	:	o_val <= 16'b0101100111100101;
            14'h1fba 	:	o_val <= 16'b0101100111100111;
            14'h1fbb 	:	o_val <= 16'b0101100111101001;
            14'h1fbc 	:	o_val <= 16'b0101100111101100;
            14'h1fbd 	:	o_val <= 16'b0101100111101110;
            14'h1fbe 	:	o_val <= 16'b0101100111110000;
            14'h1fbf 	:	o_val <= 16'b0101100111110010;
            14'h1fc0 	:	o_val <= 16'b0101100111110100;
            14'h1fc1 	:	o_val <= 16'b0101100111110111;
            14'h1fc2 	:	o_val <= 16'b0101100111111001;
            14'h1fc3 	:	o_val <= 16'b0101100111111011;
            14'h1fc4 	:	o_val <= 16'b0101100111111101;
            14'h1fc5 	:	o_val <= 16'b0101101000000000;
            14'h1fc6 	:	o_val <= 16'b0101101000000010;
            14'h1fc7 	:	o_val <= 16'b0101101000000100;
            14'h1fc8 	:	o_val <= 16'b0101101000000110;
            14'h1fc9 	:	o_val <= 16'b0101101000001001;
            14'h1fca 	:	o_val <= 16'b0101101000001011;
            14'h1fcb 	:	o_val <= 16'b0101101000001101;
            14'h1fcc 	:	o_val <= 16'b0101101000001111;
            14'h1fcd 	:	o_val <= 16'b0101101000010010;
            14'h1fce 	:	o_val <= 16'b0101101000010100;
            14'h1fcf 	:	o_val <= 16'b0101101000010110;
            14'h1fd0 	:	o_val <= 16'b0101101000011000;
            14'h1fd1 	:	o_val <= 16'b0101101000011010;
            14'h1fd2 	:	o_val <= 16'b0101101000011101;
            14'h1fd3 	:	o_val <= 16'b0101101000011111;
            14'h1fd4 	:	o_val <= 16'b0101101000100001;
            14'h1fd5 	:	o_val <= 16'b0101101000100011;
            14'h1fd6 	:	o_val <= 16'b0101101000100110;
            14'h1fd7 	:	o_val <= 16'b0101101000101000;
            14'h1fd8 	:	o_val <= 16'b0101101000101010;
            14'h1fd9 	:	o_val <= 16'b0101101000101100;
            14'h1fda 	:	o_val <= 16'b0101101000101111;
            14'h1fdb 	:	o_val <= 16'b0101101000110001;
            14'h1fdc 	:	o_val <= 16'b0101101000110011;
            14'h1fdd 	:	o_val <= 16'b0101101000110101;
            14'h1fde 	:	o_val <= 16'b0101101000110111;
            14'h1fdf 	:	o_val <= 16'b0101101000111010;
            14'h1fe0 	:	o_val <= 16'b0101101000111100;
            14'h1fe1 	:	o_val <= 16'b0101101000111110;
            14'h1fe2 	:	o_val <= 16'b0101101001000000;
            14'h1fe3 	:	o_val <= 16'b0101101001000011;
            14'h1fe4 	:	o_val <= 16'b0101101001000101;
            14'h1fe5 	:	o_val <= 16'b0101101001000111;
            14'h1fe6 	:	o_val <= 16'b0101101001001001;
            14'h1fe7 	:	o_val <= 16'b0101101001001011;
            14'h1fe8 	:	o_val <= 16'b0101101001001110;
            14'h1fe9 	:	o_val <= 16'b0101101001010000;
            14'h1fea 	:	o_val <= 16'b0101101001010010;
            14'h1feb 	:	o_val <= 16'b0101101001010100;
            14'h1fec 	:	o_val <= 16'b0101101001010111;
            14'h1fed 	:	o_val <= 16'b0101101001011001;
            14'h1fee 	:	o_val <= 16'b0101101001011011;
            14'h1fef 	:	o_val <= 16'b0101101001011101;
            14'h1ff0 	:	o_val <= 16'b0101101001100000;
            14'h1ff1 	:	o_val <= 16'b0101101001100010;
            14'h1ff2 	:	o_val <= 16'b0101101001100100;
            14'h1ff3 	:	o_val <= 16'b0101101001100110;
            14'h1ff4 	:	o_val <= 16'b0101101001101000;
            14'h1ff5 	:	o_val <= 16'b0101101001101011;
            14'h1ff6 	:	o_val <= 16'b0101101001101101;
            14'h1ff7 	:	o_val <= 16'b0101101001101111;
            14'h1ff8 	:	o_val <= 16'b0101101001110001;
            14'h1ff9 	:	o_val <= 16'b0101101001110100;
            14'h1ffa 	:	o_val <= 16'b0101101001110110;
            14'h1ffb 	:	o_val <= 16'b0101101001111000;
            14'h1ffc 	:	o_val <= 16'b0101101001111010;
            14'h1ffd 	:	o_val <= 16'b0101101001111100;
            14'h1ffe 	:	o_val <= 16'b0101101001111111;
            14'h1fff 	:	o_val <= 16'b0101101010000001;
            14'h2000 	:	o_val <= 16'b0101101010000011;
            14'h2001 	:	o_val <= 16'b0101101010000101;
            14'h2002 	:	o_val <= 16'b0101101010001000;
            14'h2003 	:	o_val <= 16'b0101101010001010;
            14'h2004 	:	o_val <= 16'b0101101010001100;
            14'h2005 	:	o_val <= 16'b0101101010001110;
            14'h2006 	:	o_val <= 16'b0101101010010000;
            14'h2007 	:	o_val <= 16'b0101101010010011;
            14'h2008 	:	o_val <= 16'b0101101010010101;
            14'h2009 	:	o_val <= 16'b0101101010010111;
            14'h200a 	:	o_val <= 16'b0101101010011001;
            14'h200b 	:	o_val <= 16'b0101101010011100;
            14'h200c 	:	o_val <= 16'b0101101010011110;
            14'h200d 	:	o_val <= 16'b0101101010100000;
            14'h200e 	:	o_val <= 16'b0101101010100010;
            14'h200f 	:	o_val <= 16'b0101101010100100;
            14'h2010 	:	o_val <= 16'b0101101010100111;
            14'h2011 	:	o_val <= 16'b0101101010101001;
            14'h2012 	:	o_val <= 16'b0101101010101011;
            14'h2013 	:	o_val <= 16'b0101101010101101;
            14'h2014 	:	o_val <= 16'b0101101010101111;
            14'h2015 	:	o_val <= 16'b0101101010110010;
            14'h2016 	:	o_val <= 16'b0101101010110100;
            14'h2017 	:	o_val <= 16'b0101101010110110;
            14'h2018 	:	o_val <= 16'b0101101010111000;
            14'h2019 	:	o_val <= 16'b0101101010111011;
            14'h201a 	:	o_val <= 16'b0101101010111101;
            14'h201b 	:	o_val <= 16'b0101101010111111;
            14'h201c 	:	o_val <= 16'b0101101011000001;
            14'h201d 	:	o_val <= 16'b0101101011000011;
            14'h201e 	:	o_val <= 16'b0101101011000110;
            14'h201f 	:	o_val <= 16'b0101101011001000;
            14'h2020 	:	o_val <= 16'b0101101011001010;
            14'h2021 	:	o_val <= 16'b0101101011001100;
            14'h2022 	:	o_val <= 16'b0101101011001110;
            14'h2023 	:	o_val <= 16'b0101101011010001;
            14'h2024 	:	o_val <= 16'b0101101011010011;
            14'h2025 	:	o_val <= 16'b0101101011010101;
            14'h2026 	:	o_val <= 16'b0101101011010111;
            14'h2027 	:	o_val <= 16'b0101101011011010;
            14'h2028 	:	o_val <= 16'b0101101011011100;
            14'h2029 	:	o_val <= 16'b0101101011011110;
            14'h202a 	:	o_val <= 16'b0101101011100000;
            14'h202b 	:	o_val <= 16'b0101101011100010;
            14'h202c 	:	o_val <= 16'b0101101011100101;
            14'h202d 	:	o_val <= 16'b0101101011100111;
            14'h202e 	:	o_val <= 16'b0101101011101001;
            14'h202f 	:	o_val <= 16'b0101101011101011;
            14'h2030 	:	o_val <= 16'b0101101011101101;
            14'h2031 	:	o_val <= 16'b0101101011110000;
            14'h2032 	:	o_val <= 16'b0101101011110010;
            14'h2033 	:	o_val <= 16'b0101101011110100;
            14'h2034 	:	o_val <= 16'b0101101011110110;
            14'h2035 	:	o_val <= 16'b0101101011111001;
            14'h2036 	:	o_val <= 16'b0101101011111011;
            14'h2037 	:	o_val <= 16'b0101101011111101;
            14'h2038 	:	o_val <= 16'b0101101011111111;
            14'h2039 	:	o_val <= 16'b0101101100000001;
            14'h203a 	:	o_val <= 16'b0101101100000100;
            14'h203b 	:	o_val <= 16'b0101101100000110;
            14'h203c 	:	o_val <= 16'b0101101100001000;
            14'h203d 	:	o_val <= 16'b0101101100001010;
            14'h203e 	:	o_val <= 16'b0101101100001100;
            14'h203f 	:	o_val <= 16'b0101101100001111;
            14'h2040 	:	o_val <= 16'b0101101100010001;
            14'h2041 	:	o_val <= 16'b0101101100010011;
            14'h2042 	:	o_val <= 16'b0101101100010101;
            14'h2043 	:	o_val <= 16'b0101101100010111;
            14'h2044 	:	o_val <= 16'b0101101100011010;
            14'h2045 	:	o_val <= 16'b0101101100011100;
            14'h2046 	:	o_val <= 16'b0101101100011110;
            14'h2047 	:	o_val <= 16'b0101101100100000;
            14'h2048 	:	o_val <= 16'b0101101100100010;
            14'h2049 	:	o_val <= 16'b0101101100100101;
            14'h204a 	:	o_val <= 16'b0101101100100111;
            14'h204b 	:	o_val <= 16'b0101101100101001;
            14'h204c 	:	o_val <= 16'b0101101100101011;
            14'h204d 	:	o_val <= 16'b0101101100101101;
            14'h204e 	:	o_val <= 16'b0101101100110000;
            14'h204f 	:	o_val <= 16'b0101101100110010;
            14'h2050 	:	o_val <= 16'b0101101100110100;
            14'h2051 	:	o_val <= 16'b0101101100110110;
            14'h2052 	:	o_val <= 16'b0101101100111001;
            14'h2053 	:	o_val <= 16'b0101101100111011;
            14'h2054 	:	o_val <= 16'b0101101100111101;
            14'h2055 	:	o_val <= 16'b0101101100111111;
            14'h2056 	:	o_val <= 16'b0101101101000001;
            14'h2057 	:	o_val <= 16'b0101101101000100;
            14'h2058 	:	o_val <= 16'b0101101101000110;
            14'h2059 	:	o_val <= 16'b0101101101001000;
            14'h205a 	:	o_val <= 16'b0101101101001010;
            14'h205b 	:	o_val <= 16'b0101101101001100;
            14'h205c 	:	o_val <= 16'b0101101101001111;
            14'h205d 	:	o_val <= 16'b0101101101010001;
            14'h205e 	:	o_val <= 16'b0101101101010011;
            14'h205f 	:	o_val <= 16'b0101101101010101;
            14'h2060 	:	o_val <= 16'b0101101101010111;
            14'h2061 	:	o_val <= 16'b0101101101011010;
            14'h2062 	:	o_val <= 16'b0101101101011100;
            14'h2063 	:	o_val <= 16'b0101101101011110;
            14'h2064 	:	o_val <= 16'b0101101101100000;
            14'h2065 	:	o_val <= 16'b0101101101100010;
            14'h2066 	:	o_val <= 16'b0101101101100101;
            14'h2067 	:	o_val <= 16'b0101101101100111;
            14'h2068 	:	o_val <= 16'b0101101101101001;
            14'h2069 	:	o_val <= 16'b0101101101101011;
            14'h206a 	:	o_val <= 16'b0101101101101101;
            14'h206b 	:	o_val <= 16'b0101101101110000;
            14'h206c 	:	o_val <= 16'b0101101101110010;
            14'h206d 	:	o_val <= 16'b0101101101110100;
            14'h206e 	:	o_val <= 16'b0101101101110110;
            14'h206f 	:	o_val <= 16'b0101101101111000;
            14'h2070 	:	o_val <= 16'b0101101101111011;
            14'h2071 	:	o_val <= 16'b0101101101111101;
            14'h2072 	:	o_val <= 16'b0101101101111111;
            14'h2073 	:	o_val <= 16'b0101101110000001;
            14'h2074 	:	o_val <= 16'b0101101110000011;
            14'h2075 	:	o_val <= 16'b0101101110000110;
            14'h2076 	:	o_val <= 16'b0101101110001000;
            14'h2077 	:	o_val <= 16'b0101101110001010;
            14'h2078 	:	o_val <= 16'b0101101110001100;
            14'h2079 	:	o_val <= 16'b0101101110001110;
            14'h207a 	:	o_val <= 16'b0101101110010000;
            14'h207b 	:	o_val <= 16'b0101101110010011;
            14'h207c 	:	o_val <= 16'b0101101110010101;
            14'h207d 	:	o_val <= 16'b0101101110010111;
            14'h207e 	:	o_val <= 16'b0101101110011001;
            14'h207f 	:	o_val <= 16'b0101101110011011;
            14'h2080 	:	o_val <= 16'b0101101110011110;
            14'h2081 	:	o_val <= 16'b0101101110100000;
            14'h2082 	:	o_val <= 16'b0101101110100010;
            14'h2083 	:	o_val <= 16'b0101101110100100;
            14'h2084 	:	o_val <= 16'b0101101110100110;
            14'h2085 	:	o_val <= 16'b0101101110101001;
            14'h2086 	:	o_val <= 16'b0101101110101011;
            14'h2087 	:	o_val <= 16'b0101101110101101;
            14'h2088 	:	o_val <= 16'b0101101110101111;
            14'h2089 	:	o_val <= 16'b0101101110110001;
            14'h208a 	:	o_val <= 16'b0101101110110100;
            14'h208b 	:	o_val <= 16'b0101101110110110;
            14'h208c 	:	o_val <= 16'b0101101110111000;
            14'h208d 	:	o_val <= 16'b0101101110111010;
            14'h208e 	:	o_val <= 16'b0101101110111100;
            14'h208f 	:	o_val <= 16'b0101101110111111;
            14'h2090 	:	o_val <= 16'b0101101111000001;
            14'h2091 	:	o_val <= 16'b0101101111000011;
            14'h2092 	:	o_val <= 16'b0101101111000101;
            14'h2093 	:	o_val <= 16'b0101101111000111;
            14'h2094 	:	o_val <= 16'b0101101111001001;
            14'h2095 	:	o_val <= 16'b0101101111001100;
            14'h2096 	:	o_val <= 16'b0101101111001110;
            14'h2097 	:	o_val <= 16'b0101101111010000;
            14'h2098 	:	o_val <= 16'b0101101111010010;
            14'h2099 	:	o_val <= 16'b0101101111010100;
            14'h209a 	:	o_val <= 16'b0101101111010111;
            14'h209b 	:	o_val <= 16'b0101101111011001;
            14'h209c 	:	o_val <= 16'b0101101111011011;
            14'h209d 	:	o_val <= 16'b0101101111011101;
            14'h209e 	:	o_val <= 16'b0101101111011111;
            14'h209f 	:	o_val <= 16'b0101101111100010;
            14'h20a0 	:	o_val <= 16'b0101101111100100;
            14'h20a1 	:	o_val <= 16'b0101101111100110;
            14'h20a2 	:	o_val <= 16'b0101101111101000;
            14'h20a3 	:	o_val <= 16'b0101101111101010;
            14'h20a4 	:	o_val <= 16'b0101101111101101;
            14'h20a5 	:	o_val <= 16'b0101101111101111;
            14'h20a6 	:	o_val <= 16'b0101101111110001;
            14'h20a7 	:	o_val <= 16'b0101101111110011;
            14'h20a8 	:	o_val <= 16'b0101101111110101;
            14'h20a9 	:	o_val <= 16'b0101101111110111;
            14'h20aa 	:	o_val <= 16'b0101101111111010;
            14'h20ab 	:	o_val <= 16'b0101101111111100;
            14'h20ac 	:	o_val <= 16'b0101101111111110;
            14'h20ad 	:	o_val <= 16'b0101110000000000;
            14'h20ae 	:	o_val <= 16'b0101110000000010;
            14'h20af 	:	o_val <= 16'b0101110000000101;
            14'h20b0 	:	o_val <= 16'b0101110000000111;
            14'h20b1 	:	o_val <= 16'b0101110000001001;
            14'h20b2 	:	o_val <= 16'b0101110000001011;
            14'h20b3 	:	o_val <= 16'b0101110000001101;
            14'h20b4 	:	o_val <= 16'b0101110000001111;
            14'h20b5 	:	o_val <= 16'b0101110000010010;
            14'h20b6 	:	o_val <= 16'b0101110000010100;
            14'h20b7 	:	o_val <= 16'b0101110000010110;
            14'h20b8 	:	o_val <= 16'b0101110000011000;
            14'h20b9 	:	o_val <= 16'b0101110000011010;
            14'h20ba 	:	o_val <= 16'b0101110000011101;
            14'h20bb 	:	o_val <= 16'b0101110000011111;
            14'h20bc 	:	o_val <= 16'b0101110000100001;
            14'h20bd 	:	o_val <= 16'b0101110000100011;
            14'h20be 	:	o_val <= 16'b0101110000100101;
            14'h20bf 	:	o_val <= 16'b0101110000100111;
            14'h20c0 	:	o_val <= 16'b0101110000101010;
            14'h20c1 	:	o_val <= 16'b0101110000101100;
            14'h20c2 	:	o_val <= 16'b0101110000101110;
            14'h20c3 	:	o_val <= 16'b0101110000110000;
            14'h20c4 	:	o_val <= 16'b0101110000110010;
            14'h20c5 	:	o_val <= 16'b0101110000110101;
            14'h20c6 	:	o_val <= 16'b0101110000110111;
            14'h20c7 	:	o_val <= 16'b0101110000111001;
            14'h20c8 	:	o_val <= 16'b0101110000111011;
            14'h20c9 	:	o_val <= 16'b0101110000111101;
            14'h20ca 	:	o_val <= 16'b0101110000111111;
            14'h20cb 	:	o_val <= 16'b0101110001000010;
            14'h20cc 	:	o_val <= 16'b0101110001000100;
            14'h20cd 	:	o_val <= 16'b0101110001000110;
            14'h20ce 	:	o_val <= 16'b0101110001001000;
            14'h20cf 	:	o_val <= 16'b0101110001001010;
            14'h20d0 	:	o_val <= 16'b0101110001001100;
            14'h20d1 	:	o_val <= 16'b0101110001001111;
            14'h20d2 	:	o_val <= 16'b0101110001010001;
            14'h20d3 	:	o_val <= 16'b0101110001010011;
            14'h20d4 	:	o_val <= 16'b0101110001010101;
            14'h20d5 	:	o_val <= 16'b0101110001010111;
            14'h20d6 	:	o_val <= 16'b0101110001011010;
            14'h20d7 	:	o_val <= 16'b0101110001011100;
            14'h20d8 	:	o_val <= 16'b0101110001011110;
            14'h20d9 	:	o_val <= 16'b0101110001100000;
            14'h20da 	:	o_val <= 16'b0101110001100010;
            14'h20db 	:	o_val <= 16'b0101110001100100;
            14'h20dc 	:	o_val <= 16'b0101110001100111;
            14'h20dd 	:	o_val <= 16'b0101110001101001;
            14'h20de 	:	o_val <= 16'b0101110001101011;
            14'h20df 	:	o_val <= 16'b0101110001101101;
            14'h20e0 	:	o_val <= 16'b0101110001101111;
            14'h20e1 	:	o_val <= 16'b0101110001110001;
            14'h20e2 	:	o_val <= 16'b0101110001110100;
            14'h20e3 	:	o_val <= 16'b0101110001110110;
            14'h20e4 	:	o_val <= 16'b0101110001111000;
            14'h20e5 	:	o_val <= 16'b0101110001111010;
            14'h20e6 	:	o_val <= 16'b0101110001111100;
            14'h20e7 	:	o_val <= 16'b0101110001111110;
            14'h20e8 	:	o_val <= 16'b0101110010000001;
            14'h20e9 	:	o_val <= 16'b0101110010000011;
            14'h20ea 	:	o_val <= 16'b0101110010000101;
            14'h20eb 	:	o_val <= 16'b0101110010000111;
            14'h20ec 	:	o_val <= 16'b0101110010001001;
            14'h20ed 	:	o_val <= 16'b0101110010001100;
            14'h20ee 	:	o_val <= 16'b0101110010001110;
            14'h20ef 	:	o_val <= 16'b0101110010010000;
            14'h20f0 	:	o_val <= 16'b0101110010010010;
            14'h20f1 	:	o_val <= 16'b0101110010010100;
            14'h20f2 	:	o_val <= 16'b0101110010010110;
            14'h20f3 	:	o_val <= 16'b0101110010011001;
            14'h20f4 	:	o_val <= 16'b0101110010011011;
            14'h20f5 	:	o_val <= 16'b0101110010011101;
            14'h20f6 	:	o_val <= 16'b0101110010011111;
            14'h20f7 	:	o_val <= 16'b0101110010100001;
            14'h20f8 	:	o_val <= 16'b0101110010100011;
            14'h20f9 	:	o_val <= 16'b0101110010100110;
            14'h20fa 	:	o_val <= 16'b0101110010101000;
            14'h20fb 	:	o_val <= 16'b0101110010101010;
            14'h20fc 	:	o_val <= 16'b0101110010101100;
            14'h20fd 	:	o_val <= 16'b0101110010101110;
            14'h20fe 	:	o_val <= 16'b0101110010110000;
            14'h20ff 	:	o_val <= 16'b0101110010110011;
            14'h2100 	:	o_val <= 16'b0101110010110101;
            14'h2101 	:	o_val <= 16'b0101110010110111;
            14'h2102 	:	o_val <= 16'b0101110010111001;
            14'h2103 	:	o_val <= 16'b0101110010111011;
            14'h2104 	:	o_val <= 16'b0101110010111101;
            14'h2105 	:	o_val <= 16'b0101110011000000;
            14'h2106 	:	o_val <= 16'b0101110011000010;
            14'h2107 	:	o_val <= 16'b0101110011000100;
            14'h2108 	:	o_val <= 16'b0101110011000110;
            14'h2109 	:	o_val <= 16'b0101110011001000;
            14'h210a 	:	o_val <= 16'b0101110011001010;
            14'h210b 	:	o_val <= 16'b0101110011001101;
            14'h210c 	:	o_val <= 16'b0101110011001111;
            14'h210d 	:	o_val <= 16'b0101110011010001;
            14'h210e 	:	o_val <= 16'b0101110011010011;
            14'h210f 	:	o_val <= 16'b0101110011010101;
            14'h2110 	:	o_val <= 16'b0101110011010111;
            14'h2111 	:	o_val <= 16'b0101110011011010;
            14'h2112 	:	o_val <= 16'b0101110011011100;
            14'h2113 	:	o_val <= 16'b0101110011011110;
            14'h2114 	:	o_val <= 16'b0101110011100000;
            14'h2115 	:	o_val <= 16'b0101110011100010;
            14'h2116 	:	o_val <= 16'b0101110011100100;
            14'h2117 	:	o_val <= 16'b0101110011100110;
            14'h2118 	:	o_val <= 16'b0101110011101001;
            14'h2119 	:	o_val <= 16'b0101110011101011;
            14'h211a 	:	o_val <= 16'b0101110011101101;
            14'h211b 	:	o_val <= 16'b0101110011101111;
            14'h211c 	:	o_val <= 16'b0101110011110001;
            14'h211d 	:	o_val <= 16'b0101110011110011;
            14'h211e 	:	o_val <= 16'b0101110011110110;
            14'h211f 	:	o_val <= 16'b0101110011111000;
            14'h2120 	:	o_val <= 16'b0101110011111010;
            14'h2121 	:	o_val <= 16'b0101110011111100;
            14'h2122 	:	o_val <= 16'b0101110011111110;
            14'h2123 	:	o_val <= 16'b0101110100000000;
            14'h2124 	:	o_val <= 16'b0101110100000011;
            14'h2125 	:	o_val <= 16'b0101110100000101;
            14'h2126 	:	o_val <= 16'b0101110100000111;
            14'h2127 	:	o_val <= 16'b0101110100001001;
            14'h2128 	:	o_val <= 16'b0101110100001011;
            14'h2129 	:	o_val <= 16'b0101110100001101;
            14'h212a 	:	o_val <= 16'b0101110100001111;
            14'h212b 	:	o_val <= 16'b0101110100010010;
            14'h212c 	:	o_val <= 16'b0101110100010100;
            14'h212d 	:	o_val <= 16'b0101110100010110;
            14'h212e 	:	o_val <= 16'b0101110100011000;
            14'h212f 	:	o_val <= 16'b0101110100011010;
            14'h2130 	:	o_val <= 16'b0101110100011100;
            14'h2131 	:	o_val <= 16'b0101110100011111;
            14'h2132 	:	o_val <= 16'b0101110100100001;
            14'h2133 	:	o_val <= 16'b0101110100100011;
            14'h2134 	:	o_val <= 16'b0101110100100101;
            14'h2135 	:	o_val <= 16'b0101110100100111;
            14'h2136 	:	o_val <= 16'b0101110100101001;
            14'h2137 	:	o_val <= 16'b0101110100101100;
            14'h2138 	:	o_val <= 16'b0101110100101110;
            14'h2139 	:	o_val <= 16'b0101110100110000;
            14'h213a 	:	o_val <= 16'b0101110100110010;
            14'h213b 	:	o_val <= 16'b0101110100110100;
            14'h213c 	:	o_val <= 16'b0101110100110110;
            14'h213d 	:	o_val <= 16'b0101110100111000;
            14'h213e 	:	o_val <= 16'b0101110100111011;
            14'h213f 	:	o_val <= 16'b0101110100111101;
            14'h2140 	:	o_val <= 16'b0101110100111111;
            14'h2141 	:	o_val <= 16'b0101110101000001;
            14'h2142 	:	o_val <= 16'b0101110101000011;
            14'h2143 	:	o_val <= 16'b0101110101000101;
            14'h2144 	:	o_val <= 16'b0101110101001000;
            14'h2145 	:	o_val <= 16'b0101110101001010;
            14'h2146 	:	o_val <= 16'b0101110101001100;
            14'h2147 	:	o_val <= 16'b0101110101001110;
            14'h2148 	:	o_val <= 16'b0101110101010000;
            14'h2149 	:	o_val <= 16'b0101110101010010;
            14'h214a 	:	o_val <= 16'b0101110101010100;
            14'h214b 	:	o_val <= 16'b0101110101010111;
            14'h214c 	:	o_val <= 16'b0101110101011001;
            14'h214d 	:	o_val <= 16'b0101110101011011;
            14'h214e 	:	o_val <= 16'b0101110101011101;
            14'h214f 	:	o_val <= 16'b0101110101011111;
            14'h2150 	:	o_val <= 16'b0101110101100001;
            14'h2151 	:	o_val <= 16'b0101110101100011;
            14'h2152 	:	o_val <= 16'b0101110101100110;
            14'h2153 	:	o_val <= 16'b0101110101101000;
            14'h2154 	:	o_val <= 16'b0101110101101010;
            14'h2155 	:	o_val <= 16'b0101110101101100;
            14'h2156 	:	o_val <= 16'b0101110101101110;
            14'h2157 	:	o_val <= 16'b0101110101110000;
            14'h2158 	:	o_val <= 16'b0101110101110010;
            14'h2159 	:	o_val <= 16'b0101110101110101;
            14'h215a 	:	o_val <= 16'b0101110101110111;
            14'h215b 	:	o_val <= 16'b0101110101111001;
            14'h215c 	:	o_val <= 16'b0101110101111011;
            14'h215d 	:	o_val <= 16'b0101110101111101;
            14'h215e 	:	o_val <= 16'b0101110101111111;
            14'h215f 	:	o_val <= 16'b0101110110000010;
            14'h2160 	:	o_val <= 16'b0101110110000100;
            14'h2161 	:	o_val <= 16'b0101110110000110;
            14'h2162 	:	o_val <= 16'b0101110110001000;
            14'h2163 	:	o_val <= 16'b0101110110001010;
            14'h2164 	:	o_val <= 16'b0101110110001100;
            14'h2165 	:	o_val <= 16'b0101110110001110;
            14'h2166 	:	o_val <= 16'b0101110110010001;
            14'h2167 	:	o_val <= 16'b0101110110010011;
            14'h2168 	:	o_val <= 16'b0101110110010101;
            14'h2169 	:	o_val <= 16'b0101110110010111;
            14'h216a 	:	o_val <= 16'b0101110110011001;
            14'h216b 	:	o_val <= 16'b0101110110011011;
            14'h216c 	:	o_val <= 16'b0101110110011101;
            14'h216d 	:	o_val <= 16'b0101110110100000;
            14'h216e 	:	o_val <= 16'b0101110110100010;
            14'h216f 	:	o_val <= 16'b0101110110100100;
            14'h2170 	:	o_val <= 16'b0101110110100110;
            14'h2171 	:	o_val <= 16'b0101110110101000;
            14'h2172 	:	o_val <= 16'b0101110110101010;
            14'h2173 	:	o_val <= 16'b0101110110101100;
            14'h2174 	:	o_val <= 16'b0101110110101111;
            14'h2175 	:	o_val <= 16'b0101110110110001;
            14'h2176 	:	o_val <= 16'b0101110110110011;
            14'h2177 	:	o_val <= 16'b0101110110110101;
            14'h2178 	:	o_val <= 16'b0101110110110111;
            14'h2179 	:	o_val <= 16'b0101110110111001;
            14'h217a 	:	o_val <= 16'b0101110110111011;
            14'h217b 	:	o_val <= 16'b0101110110111101;
            14'h217c 	:	o_val <= 16'b0101110111000000;
            14'h217d 	:	o_val <= 16'b0101110111000010;
            14'h217e 	:	o_val <= 16'b0101110111000100;
            14'h217f 	:	o_val <= 16'b0101110111000110;
            14'h2180 	:	o_val <= 16'b0101110111001000;
            14'h2181 	:	o_val <= 16'b0101110111001010;
            14'h2182 	:	o_val <= 16'b0101110111001100;
            14'h2183 	:	o_val <= 16'b0101110111001111;
            14'h2184 	:	o_val <= 16'b0101110111010001;
            14'h2185 	:	o_val <= 16'b0101110111010011;
            14'h2186 	:	o_val <= 16'b0101110111010101;
            14'h2187 	:	o_val <= 16'b0101110111010111;
            14'h2188 	:	o_val <= 16'b0101110111011001;
            14'h2189 	:	o_val <= 16'b0101110111011011;
            14'h218a 	:	o_val <= 16'b0101110111011110;
            14'h218b 	:	o_val <= 16'b0101110111100000;
            14'h218c 	:	o_val <= 16'b0101110111100010;
            14'h218d 	:	o_val <= 16'b0101110111100100;
            14'h218e 	:	o_val <= 16'b0101110111100110;
            14'h218f 	:	o_val <= 16'b0101110111101000;
            14'h2190 	:	o_val <= 16'b0101110111101010;
            14'h2191 	:	o_val <= 16'b0101110111101100;
            14'h2192 	:	o_val <= 16'b0101110111101111;
            14'h2193 	:	o_val <= 16'b0101110111110001;
            14'h2194 	:	o_val <= 16'b0101110111110011;
            14'h2195 	:	o_val <= 16'b0101110111110101;
            14'h2196 	:	o_val <= 16'b0101110111110111;
            14'h2197 	:	o_val <= 16'b0101110111111001;
            14'h2198 	:	o_val <= 16'b0101110111111011;
            14'h2199 	:	o_val <= 16'b0101110111111110;
            14'h219a 	:	o_val <= 16'b0101111000000000;
            14'h219b 	:	o_val <= 16'b0101111000000010;
            14'h219c 	:	o_val <= 16'b0101111000000100;
            14'h219d 	:	o_val <= 16'b0101111000000110;
            14'h219e 	:	o_val <= 16'b0101111000001000;
            14'h219f 	:	o_val <= 16'b0101111000001010;
            14'h21a0 	:	o_val <= 16'b0101111000001100;
            14'h21a1 	:	o_val <= 16'b0101111000001111;
            14'h21a2 	:	o_val <= 16'b0101111000010001;
            14'h21a3 	:	o_val <= 16'b0101111000010011;
            14'h21a4 	:	o_val <= 16'b0101111000010101;
            14'h21a5 	:	o_val <= 16'b0101111000010111;
            14'h21a6 	:	o_val <= 16'b0101111000011001;
            14'h21a7 	:	o_val <= 16'b0101111000011011;
            14'h21a8 	:	o_val <= 16'b0101111000011110;
            14'h21a9 	:	o_val <= 16'b0101111000100000;
            14'h21aa 	:	o_val <= 16'b0101111000100010;
            14'h21ab 	:	o_val <= 16'b0101111000100100;
            14'h21ac 	:	o_val <= 16'b0101111000100110;
            14'h21ad 	:	o_val <= 16'b0101111000101000;
            14'h21ae 	:	o_val <= 16'b0101111000101010;
            14'h21af 	:	o_val <= 16'b0101111000101100;
            14'h21b0 	:	o_val <= 16'b0101111000101111;
            14'h21b1 	:	o_val <= 16'b0101111000110001;
            14'h21b2 	:	o_val <= 16'b0101111000110011;
            14'h21b3 	:	o_val <= 16'b0101111000110101;
            14'h21b4 	:	o_val <= 16'b0101111000110111;
            14'h21b5 	:	o_val <= 16'b0101111000111001;
            14'h21b6 	:	o_val <= 16'b0101111000111011;
            14'h21b7 	:	o_val <= 16'b0101111000111101;
            14'h21b8 	:	o_val <= 16'b0101111001000000;
            14'h21b9 	:	o_val <= 16'b0101111001000010;
            14'h21ba 	:	o_val <= 16'b0101111001000100;
            14'h21bb 	:	o_val <= 16'b0101111001000110;
            14'h21bc 	:	o_val <= 16'b0101111001001000;
            14'h21bd 	:	o_val <= 16'b0101111001001010;
            14'h21be 	:	o_val <= 16'b0101111001001100;
            14'h21bf 	:	o_val <= 16'b0101111001001110;
            14'h21c0 	:	o_val <= 16'b0101111001010001;
            14'h21c1 	:	o_val <= 16'b0101111001010011;
            14'h21c2 	:	o_val <= 16'b0101111001010101;
            14'h21c3 	:	o_val <= 16'b0101111001010111;
            14'h21c4 	:	o_val <= 16'b0101111001011001;
            14'h21c5 	:	o_val <= 16'b0101111001011011;
            14'h21c6 	:	o_val <= 16'b0101111001011101;
            14'h21c7 	:	o_val <= 16'b0101111001011111;
            14'h21c8 	:	o_val <= 16'b0101111001100010;
            14'h21c9 	:	o_val <= 16'b0101111001100100;
            14'h21ca 	:	o_val <= 16'b0101111001100110;
            14'h21cb 	:	o_val <= 16'b0101111001101000;
            14'h21cc 	:	o_val <= 16'b0101111001101010;
            14'h21cd 	:	o_val <= 16'b0101111001101100;
            14'h21ce 	:	o_val <= 16'b0101111001101110;
            14'h21cf 	:	o_val <= 16'b0101111001110000;
            14'h21d0 	:	o_val <= 16'b0101111001110011;
            14'h21d1 	:	o_val <= 16'b0101111001110101;
            14'h21d2 	:	o_val <= 16'b0101111001110111;
            14'h21d3 	:	o_val <= 16'b0101111001111001;
            14'h21d4 	:	o_val <= 16'b0101111001111011;
            14'h21d5 	:	o_val <= 16'b0101111001111101;
            14'h21d6 	:	o_val <= 16'b0101111001111111;
            14'h21d7 	:	o_val <= 16'b0101111010000001;
            14'h21d8 	:	o_val <= 16'b0101111010000011;
            14'h21d9 	:	o_val <= 16'b0101111010000110;
            14'h21da 	:	o_val <= 16'b0101111010001000;
            14'h21db 	:	o_val <= 16'b0101111010001010;
            14'h21dc 	:	o_val <= 16'b0101111010001100;
            14'h21dd 	:	o_val <= 16'b0101111010001110;
            14'h21de 	:	o_val <= 16'b0101111010010000;
            14'h21df 	:	o_val <= 16'b0101111010010010;
            14'h21e0 	:	o_val <= 16'b0101111010010100;
            14'h21e1 	:	o_val <= 16'b0101111010010111;
            14'h21e2 	:	o_val <= 16'b0101111010011001;
            14'h21e3 	:	o_val <= 16'b0101111010011011;
            14'h21e4 	:	o_val <= 16'b0101111010011101;
            14'h21e5 	:	o_val <= 16'b0101111010011111;
            14'h21e6 	:	o_val <= 16'b0101111010100001;
            14'h21e7 	:	o_val <= 16'b0101111010100011;
            14'h21e8 	:	o_val <= 16'b0101111010100101;
            14'h21e9 	:	o_val <= 16'b0101111010100111;
            14'h21ea 	:	o_val <= 16'b0101111010101010;
            14'h21eb 	:	o_val <= 16'b0101111010101100;
            14'h21ec 	:	o_val <= 16'b0101111010101110;
            14'h21ed 	:	o_val <= 16'b0101111010110000;
            14'h21ee 	:	o_val <= 16'b0101111010110010;
            14'h21ef 	:	o_val <= 16'b0101111010110100;
            14'h21f0 	:	o_val <= 16'b0101111010110110;
            14'h21f1 	:	o_val <= 16'b0101111010111000;
            14'h21f2 	:	o_val <= 16'b0101111010111010;
            14'h21f3 	:	o_val <= 16'b0101111010111101;
            14'h21f4 	:	o_val <= 16'b0101111010111111;
            14'h21f5 	:	o_val <= 16'b0101111011000001;
            14'h21f6 	:	o_val <= 16'b0101111011000011;
            14'h21f7 	:	o_val <= 16'b0101111011000101;
            14'h21f8 	:	o_val <= 16'b0101111011000111;
            14'h21f9 	:	o_val <= 16'b0101111011001001;
            14'h21fa 	:	o_val <= 16'b0101111011001011;
            14'h21fb 	:	o_val <= 16'b0101111011001101;
            14'h21fc 	:	o_val <= 16'b0101111011010000;
            14'h21fd 	:	o_val <= 16'b0101111011010010;
            14'h21fe 	:	o_val <= 16'b0101111011010100;
            14'h21ff 	:	o_val <= 16'b0101111011010110;
            14'h2200 	:	o_val <= 16'b0101111011011000;
            14'h2201 	:	o_val <= 16'b0101111011011010;
            14'h2202 	:	o_val <= 16'b0101111011011100;
            14'h2203 	:	o_val <= 16'b0101111011011110;
            14'h2204 	:	o_val <= 16'b0101111011100000;
            14'h2205 	:	o_val <= 16'b0101111011100011;
            14'h2206 	:	o_val <= 16'b0101111011100101;
            14'h2207 	:	o_val <= 16'b0101111011100111;
            14'h2208 	:	o_val <= 16'b0101111011101001;
            14'h2209 	:	o_val <= 16'b0101111011101011;
            14'h220a 	:	o_val <= 16'b0101111011101101;
            14'h220b 	:	o_val <= 16'b0101111011101111;
            14'h220c 	:	o_val <= 16'b0101111011110001;
            14'h220d 	:	o_val <= 16'b0101111011110011;
            14'h220e 	:	o_val <= 16'b0101111011110110;
            14'h220f 	:	o_val <= 16'b0101111011111000;
            14'h2210 	:	o_val <= 16'b0101111011111010;
            14'h2211 	:	o_val <= 16'b0101111011111100;
            14'h2212 	:	o_val <= 16'b0101111011111110;
            14'h2213 	:	o_val <= 16'b0101111100000000;
            14'h2214 	:	o_val <= 16'b0101111100000010;
            14'h2215 	:	o_val <= 16'b0101111100000100;
            14'h2216 	:	o_val <= 16'b0101111100000110;
            14'h2217 	:	o_val <= 16'b0101111100001001;
            14'h2218 	:	o_val <= 16'b0101111100001011;
            14'h2219 	:	o_val <= 16'b0101111100001101;
            14'h221a 	:	o_val <= 16'b0101111100001111;
            14'h221b 	:	o_val <= 16'b0101111100010001;
            14'h221c 	:	o_val <= 16'b0101111100010011;
            14'h221d 	:	o_val <= 16'b0101111100010101;
            14'h221e 	:	o_val <= 16'b0101111100010111;
            14'h221f 	:	o_val <= 16'b0101111100011001;
            14'h2220 	:	o_val <= 16'b0101111100011011;
            14'h2221 	:	o_val <= 16'b0101111100011110;
            14'h2222 	:	o_val <= 16'b0101111100100000;
            14'h2223 	:	o_val <= 16'b0101111100100010;
            14'h2224 	:	o_val <= 16'b0101111100100100;
            14'h2225 	:	o_val <= 16'b0101111100100110;
            14'h2226 	:	o_val <= 16'b0101111100101000;
            14'h2227 	:	o_val <= 16'b0101111100101010;
            14'h2228 	:	o_val <= 16'b0101111100101100;
            14'h2229 	:	o_val <= 16'b0101111100101110;
            14'h222a 	:	o_val <= 16'b0101111100110000;
            14'h222b 	:	o_val <= 16'b0101111100110011;
            14'h222c 	:	o_val <= 16'b0101111100110101;
            14'h222d 	:	o_val <= 16'b0101111100110111;
            14'h222e 	:	o_val <= 16'b0101111100111001;
            14'h222f 	:	o_val <= 16'b0101111100111011;
            14'h2230 	:	o_val <= 16'b0101111100111101;
            14'h2231 	:	o_val <= 16'b0101111100111111;
            14'h2232 	:	o_val <= 16'b0101111101000001;
            14'h2233 	:	o_val <= 16'b0101111101000011;
            14'h2234 	:	o_val <= 16'b0101111101000101;
            14'h2235 	:	o_val <= 16'b0101111101001000;
            14'h2236 	:	o_val <= 16'b0101111101001010;
            14'h2237 	:	o_val <= 16'b0101111101001100;
            14'h2238 	:	o_val <= 16'b0101111101001110;
            14'h2239 	:	o_val <= 16'b0101111101010000;
            14'h223a 	:	o_val <= 16'b0101111101010010;
            14'h223b 	:	o_val <= 16'b0101111101010100;
            14'h223c 	:	o_val <= 16'b0101111101010110;
            14'h223d 	:	o_val <= 16'b0101111101011000;
            14'h223e 	:	o_val <= 16'b0101111101011010;
            14'h223f 	:	o_val <= 16'b0101111101011101;
            14'h2240 	:	o_val <= 16'b0101111101011111;
            14'h2241 	:	o_val <= 16'b0101111101100001;
            14'h2242 	:	o_val <= 16'b0101111101100011;
            14'h2243 	:	o_val <= 16'b0101111101100101;
            14'h2244 	:	o_val <= 16'b0101111101100111;
            14'h2245 	:	o_val <= 16'b0101111101101001;
            14'h2246 	:	o_val <= 16'b0101111101101011;
            14'h2247 	:	o_val <= 16'b0101111101101101;
            14'h2248 	:	o_val <= 16'b0101111101101111;
            14'h2249 	:	o_val <= 16'b0101111101110001;
            14'h224a 	:	o_val <= 16'b0101111101110100;
            14'h224b 	:	o_val <= 16'b0101111101110110;
            14'h224c 	:	o_val <= 16'b0101111101111000;
            14'h224d 	:	o_val <= 16'b0101111101111010;
            14'h224e 	:	o_val <= 16'b0101111101111100;
            14'h224f 	:	o_val <= 16'b0101111101111110;
            14'h2250 	:	o_val <= 16'b0101111110000000;
            14'h2251 	:	o_val <= 16'b0101111110000010;
            14'h2252 	:	o_val <= 16'b0101111110000100;
            14'h2253 	:	o_val <= 16'b0101111110000110;
            14'h2254 	:	o_val <= 16'b0101111110001000;
            14'h2255 	:	o_val <= 16'b0101111110001011;
            14'h2256 	:	o_val <= 16'b0101111110001101;
            14'h2257 	:	o_val <= 16'b0101111110001111;
            14'h2258 	:	o_val <= 16'b0101111110010001;
            14'h2259 	:	o_val <= 16'b0101111110010011;
            14'h225a 	:	o_val <= 16'b0101111110010101;
            14'h225b 	:	o_val <= 16'b0101111110010111;
            14'h225c 	:	o_val <= 16'b0101111110011001;
            14'h225d 	:	o_val <= 16'b0101111110011011;
            14'h225e 	:	o_val <= 16'b0101111110011101;
            14'h225f 	:	o_val <= 16'b0101111110011111;
            14'h2260 	:	o_val <= 16'b0101111110100010;
            14'h2261 	:	o_val <= 16'b0101111110100100;
            14'h2262 	:	o_val <= 16'b0101111110100110;
            14'h2263 	:	o_val <= 16'b0101111110101000;
            14'h2264 	:	o_val <= 16'b0101111110101010;
            14'h2265 	:	o_val <= 16'b0101111110101100;
            14'h2266 	:	o_val <= 16'b0101111110101110;
            14'h2267 	:	o_val <= 16'b0101111110110000;
            14'h2268 	:	o_val <= 16'b0101111110110010;
            14'h2269 	:	o_val <= 16'b0101111110110100;
            14'h226a 	:	o_val <= 16'b0101111110110110;
            14'h226b 	:	o_val <= 16'b0101111110111000;
            14'h226c 	:	o_val <= 16'b0101111110111011;
            14'h226d 	:	o_val <= 16'b0101111110111101;
            14'h226e 	:	o_val <= 16'b0101111110111111;
            14'h226f 	:	o_val <= 16'b0101111111000001;
            14'h2270 	:	o_val <= 16'b0101111111000011;
            14'h2271 	:	o_val <= 16'b0101111111000101;
            14'h2272 	:	o_val <= 16'b0101111111000111;
            14'h2273 	:	o_val <= 16'b0101111111001001;
            14'h2274 	:	o_val <= 16'b0101111111001011;
            14'h2275 	:	o_val <= 16'b0101111111001101;
            14'h2276 	:	o_val <= 16'b0101111111001111;
            14'h2277 	:	o_val <= 16'b0101111111010010;
            14'h2278 	:	o_val <= 16'b0101111111010100;
            14'h2279 	:	o_val <= 16'b0101111111010110;
            14'h227a 	:	o_val <= 16'b0101111111011000;
            14'h227b 	:	o_val <= 16'b0101111111011010;
            14'h227c 	:	o_val <= 16'b0101111111011100;
            14'h227d 	:	o_val <= 16'b0101111111011110;
            14'h227e 	:	o_val <= 16'b0101111111100000;
            14'h227f 	:	o_val <= 16'b0101111111100010;
            14'h2280 	:	o_val <= 16'b0101111111100100;
            14'h2281 	:	o_val <= 16'b0101111111100110;
            14'h2282 	:	o_val <= 16'b0101111111101000;
            14'h2283 	:	o_val <= 16'b0101111111101010;
            14'h2284 	:	o_val <= 16'b0101111111101101;
            14'h2285 	:	o_val <= 16'b0101111111101111;
            14'h2286 	:	o_val <= 16'b0101111111110001;
            14'h2287 	:	o_val <= 16'b0101111111110011;
            14'h2288 	:	o_val <= 16'b0101111111110101;
            14'h2289 	:	o_val <= 16'b0101111111110111;
            14'h228a 	:	o_val <= 16'b0101111111111001;
            14'h228b 	:	o_val <= 16'b0101111111111011;
            14'h228c 	:	o_val <= 16'b0101111111111101;
            14'h228d 	:	o_val <= 16'b0101111111111111;
            14'h228e 	:	o_val <= 16'b0110000000000001;
            14'h228f 	:	o_val <= 16'b0110000000000011;
            14'h2290 	:	o_val <= 16'b0110000000000110;
            14'h2291 	:	o_val <= 16'b0110000000001000;
            14'h2292 	:	o_val <= 16'b0110000000001010;
            14'h2293 	:	o_val <= 16'b0110000000001100;
            14'h2294 	:	o_val <= 16'b0110000000001110;
            14'h2295 	:	o_val <= 16'b0110000000010000;
            14'h2296 	:	o_val <= 16'b0110000000010010;
            14'h2297 	:	o_val <= 16'b0110000000010100;
            14'h2298 	:	o_val <= 16'b0110000000010110;
            14'h2299 	:	o_val <= 16'b0110000000011000;
            14'h229a 	:	o_val <= 16'b0110000000011010;
            14'h229b 	:	o_val <= 16'b0110000000011100;
            14'h229c 	:	o_val <= 16'b0110000000011110;
            14'h229d 	:	o_val <= 16'b0110000000100000;
            14'h229e 	:	o_val <= 16'b0110000000100011;
            14'h229f 	:	o_val <= 16'b0110000000100101;
            14'h22a0 	:	o_val <= 16'b0110000000100111;
            14'h22a1 	:	o_val <= 16'b0110000000101001;
            14'h22a2 	:	o_val <= 16'b0110000000101011;
            14'h22a3 	:	o_val <= 16'b0110000000101101;
            14'h22a4 	:	o_val <= 16'b0110000000101111;
            14'h22a5 	:	o_val <= 16'b0110000000110001;
            14'h22a6 	:	o_val <= 16'b0110000000110011;
            14'h22a7 	:	o_val <= 16'b0110000000110101;
            14'h22a8 	:	o_val <= 16'b0110000000110111;
            14'h22a9 	:	o_val <= 16'b0110000000111001;
            14'h22aa 	:	o_val <= 16'b0110000000111011;
            14'h22ab 	:	o_val <= 16'b0110000000111110;
            14'h22ac 	:	o_val <= 16'b0110000001000000;
            14'h22ad 	:	o_val <= 16'b0110000001000010;
            14'h22ae 	:	o_val <= 16'b0110000001000100;
            14'h22af 	:	o_val <= 16'b0110000001000110;
            14'h22b0 	:	o_val <= 16'b0110000001001000;
            14'h22b1 	:	o_val <= 16'b0110000001001010;
            14'h22b2 	:	o_val <= 16'b0110000001001100;
            14'h22b3 	:	o_val <= 16'b0110000001001110;
            14'h22b4 	:	o_val <= 16'b0110000001010000;
            14'h22b5 	:	o_val <= 16'b0110000001010010;
            14'h22b6 	:	o_val <= 16'b0110000001010100;
            14'h22b7 	:	o_val <= 16'b0110000001010110;
            14'h22b8 	:	o_val <= 16'b0110000001011000;
            14'h22b9 	:	o_val <= 16'b0110000001011010;
            14'h22ba 	:	o_val <= 16'b0110000001011101;
            14'h22bb 	:	o_val <= 16'b0110000001011111;
            14'h22bc 	:	o_val <= 16'b0110000001100001;
            14'h22bd 	:	o_val <= 16'b0110000001100011;
            14'h22be 	:	o_val <= 16'b0110000001100101;
            14'h22bf 	:	o_val <= 16'b0110000001100111;
            14'h22c0 	:	o_val <= 16'b0110000001101001;
            14'h22c1 	:	o_val <= 16'b0110000001101011;
            14'h22c2 	:	o_val <= 16'b0110000001101101;
            14'h22c3 	:	o_val <= 16'b0110000001101111;
            14'h22c4 	:	o_val <= 16'b0110000001110001;
            14'h22c5 	:	o_val <= 16'b0110000001110011;
            14'h22c6 	:	o_val <= 16'b0110000001110101;
            14'h22c7 	:	o_val <= 16'b0110000001110111;
            14'h22c8 	:	o_val <= 16'b0110000001111001;
            14'h22c9 	:	o_val <= 16'b0110000001111100;
            14'h22ca 	:	o_val <= 16'b0110000001111110;
            14'h22cb 	:	o_val <= 16'b0110000010000000;
            14'h22cc 	:	o_val <= 16'b0110000010000010;
            14'h22cd 	:	o_val <= 16'b0110000010000100;
            14'h22ce 	:	o_val <= 16'b0110000010000110;
            14'h22cf 	:	o_val <= 16'b0110000010001000;
            14'h22d0 	:	o_val <= 16'b0110000010001010;
            14'h22d1 	:	o_val <= 16'b0110000010001100;
            14'h22d2 	:	o_val <= 16'b0110000010001110;
            14'h22d3 	:	o_val <= 16'b0110000010010000;
            14'h22d4 	:	o_val <= 16'b0110000010010010;
            14'h22d5 	:	o_val <= 16'b0110000010010100;
            14'h22d6 	:	o_val <= 16'b0110000010010110;
            14'h22d7 	:	o_val <= 16'b0110000010011000;
            14'h22d8 	:	o_val <= 16'b0110000010011010;
            14'h22d9 	:	o_val <= 16'b0110000010011101;
            14'h22da 	:	o_val <= 16'b0110000010011111;
            14'h22db 	:	o_val <= 16'b0110000010100001;
            14'h22dc 	:	o_val <= 16'b0110000010100011;
            14'h22dd 	:	o_val <= 16'b0110000010100101;
            14'h22de 	:	o_val <= 16'b0110000010100111;
            14'h22df 	:	o_val <= 16'b0110000010101001;
            14'h22e0 	:	o_val <= 16'b0110000010101011;
            14'h22e1 	:	o_val <= 16'b0110000010101101;
            14'h22e2 	:	o_val <= 16'b0110000010101111;
            14'h22e3 	:	o_val <= 16'b0110000010110001;
            14'h22e4 	:	o_val <= 16'b0110000010110011;
            14'h22e5 	:	o_val <= 16'b0110000010110101;
            14'h22e6 	:	o_val <= 16'b0110000010110111;
            14'h22e7 	:	o_val <= 16'b0110000010111001;
            14'h22e8 	:	o_val <= 16'b0110000010111011;
            14'h22e9 	:	o_val <= 16'b0110000010111101;
            14'h22ea 	:	o_val <= 16'b0110000011000000;
            14'h22eb 	:	o_val <= 16'b0110000011000010;
            14'h22ec 	:	o_val <= 16'b0110000011000100;
            14'h22ed 	:	o_val <= 16'b0110000011000110;
            14'h22ee 	:	o_val <= 16'b0110000011001000;
            14'h22ef 	:	o_val <= 16'b0110000011001010;
            14'h22f0 	:	o_val <= 16'b0110000011001100;
            14'h22f1 	:	o_val <= 16'b0110000011001110;
            14'h22f2 	:	o_val <= 16'b0110000011010000;
            14'h22f3 	:	o_val <= 16'b0110000011010010;
            14'h22f4 	:	o_val <= 16'b0110000011010100;
            14'h22f5 	:	o_val <= 16'b0110000011010110;
            14'h22f6 	:	o_val <= 16'b0110000011011000;
            14'h22f7 	:	o_val <= 16'b0110000011011010;
            14'h22f8 	:	o_val <= 16'b0110000011011100;
            14'h22f9 	:	o_val <= 16'b0110000011011110;
            14'h22fa 	:	o_val <= 16'b0110000011100000;
            14'h22fb 	:	o_val <= 16'b0110000011100010;
            14'h22fc 	:	o_val <= 16'b0110000011100101;
            14'h22fd 	:	o_val <= 16'b0110000011100111;
            14'h22fe 	:	o_val <= 16'b0110000011101001;
            14'h22ff 	:	o_val <= 16'b0110000011101011;
            14'h2300 	:	o_val <= 16'b0110000011101101;
            14'h2301 	:	o_val <= 16'b0110000011101111;
            14'h2302 	:	o_val <= 16'b0110000011110001;
            14'h2303 	:	o_val <= 16'b0110000011110011;
            14'h2304 	:	o_val <= 16'b0110000011110101;
            14'h2305 	:	o_val <= 16'b0110000011110111;
            14'h2306 	:	o_val <= 16'b0110000011111001;
            14'h2307 	:	o_val <= 16'b0110000011111011;
            14'h2308 	:	o_val <= 16'b0110000011111101;
            14'h2309 	:	o_val <= 16'b0110000011111111;
            14'h230a 	:	o_val <= 16'b0110000100000001;
            14'h230b 	:	o_val <= 16'b0110000100000011;
            14'h230c 	:	o_val <= 16'b0110000100000101;
            14'h230d 	:	o_val <= 16'b0110000100000111;
            14'h230e 	:	o_val <= 16'b0110000100001001;
            14'h230f 	:	o_val <= 16'b0110000100001011;
            14'h2310 	:	o_val <= 16'b0110000100001110;
            14'h2311 	:	o_val <= 16'b0110000100010000;
            14'h2312 	:	o_val <= 16'b0110000100010010;
            14'h2313 	:	o_val <= 16'b0110000100010100;
            14'h2314 	:	o_val <= 16'b0110000100010110;
            14'h2315 	:	o_val <= 16'b0110000100011000;
            14'h2316 	:	o_val <= 16'b0110000100011010;
            14'h2317 	:	o_val <= 16'b0110000100011100;
            14'h2318 	:	o_val <= 16'b0110000100011110;
            14'h2319 	:	o_val <= 16'b0110000100100000;
            14'h231a 	:	o_val <= 16'b0110000100100010;
            14'h231b 	:	o_val <= 16'b0110000100100100;
            14'h231c 	:	o_val <= 16'b0110000100100110;
            14'h231d 	:	o_val <= 16'b0110000100101000;
            14'h231e 	:	o_val <= 16'b0110000100101010;
            14'h231f 	:	o_val <= 16'b0110000100101100;
            14'h2320 	:	o_val <= 16'b0110000100101110;
            14'h2321 	:	o_val <= 16'b0110000100110000;
            14'h2322 	:	o_val <= 16'b0110000100110010;
            14'h2323 	:	o_val <= 16'b0110000100110100;
            14'h2324 	:	o_val <= 16'b0110000100110110;
            14'h2325 	:	o_val <= 16'b0110000100111001;
            14'h2326 	:	o_val <= 16'b0110000100111011;
            14'h2327 	:	o_val <= 16'b0110000100111101;
            14'h2328 	:	o_val <= 16'b0110000100111111;
            14'h2329 	:	o_val <= 16'b0110000101000001;
            14'h232a 	:	o_val <= 16'b0110000101000011;
            14'h232b 	:	o_val <= 16'b0110000101000101;
            14'h232c 	:	o_val <= 16'b0110000101000111;
            14'h232d 	:	o_val <= 16'b0110000101001001;
            14'h232e 	:	o_val <= 16'b0110000101001011;
            14'h232f 	:	o_val <= 16'b0110000101001101;
            14'h2330 	:	o_val <= 16'b0110000101001111;
            14'h2331 	:	o_val <= 16'b0110000101010001;
            14'h2332 	:	o_val <= 16'b0110000101010011;
            14'h2333 	:	o_val <= 16'b0110000101010101;
            14'h2334 	:	o_val <= 16'b0110000101010111;
            14'h2335 	:	o_val <= 16'b0110000101011001;
            14'h2336 	:	o_val <= 16'b0110000101011011;
            14'h2337 	:	o_val <= 16'b0110000101011101;
            14'h2338 	:	o_val <= 16'b0110000101011111;
            14'h2339 	:	o_val <= 16'b0110000101100001;
            14'h233a 	:	o_val <= 16'b0110000101100011;
            14'h233b 	:	o_val <= 16'b0110000101100101;
            14'h233c 	:	o_val <= 16'b0110000101100111;
            14'h233d 	:	o_val <= 16'b0110000101101001;
            14'h233e 	:	o_val <= 16'b0110000101101100;
            14'h233f 	:	o_val <= 16'b0110000101101110;
            14'h2340 	:	o_val <= 16'b0110000101110000;
            14'h2341 	:	o_val <= 16'b0110000101110010;
            14'h2342 	:	o_val <= 16'b0110000101110100;
            14'h2343 	:	o_val <= 16'b0110000101110110;
            14'h2344 	:	o_val <= 16'b0110000101111000;
            14'h2345 	:	o_val <= 16'b0110000101111010;
            14'h2346 	:	o_val <= 16'b0110000101111100;
            14'h2347 	:	o_val <= 16'b0110000101111110;
            14'h2348 	:	o_val <= 16'b0110000110000000;
            14'h2349 	:	o_val <= 16'b0110000110000010;
            14'h234a 	:	o_val <= 16'b0110000110000100;
            14'h234b 	:	o_val <= 16'b0110000110000110;
            14'h234c 	:	o_val <= 16'b0110000110001000;
            14'h234d 	:	o_val <= 16'b0110000110001010;
            14'h234e 	:	o_val <= 16'b0110000110001100;
            14'h234f 	:	o_val <= 16'b0110000110001110;
            14'h2350 	:	o_val <= 16'b0110000110010000;
            14'h2351 	:	o_val <= 16'b0110000110010010;
            14'h2352 	:	o_val <= 16'b0110000110010100;
            14'h2353 	:	o_val <= 16'b0110000110010110;
            14'h2354 	:	o_val <= 16'b0110000110011000;
            14'h2355 	:	o_val <= 16'b0110000110011010;
            14'h2356 	:	o_val <= 16'b0110000110011100;
            14'h2357 	:	o_val <= 16'b0110000110011110;
            14'h2358 	:	o_val <= 16'b0110000110100000;
            14'h2359 	:	o_val <= 16'b0110000110100010;
            14'h235a 	:	o_val <= 16'b0110000110100100;
            14'h235b 	:	o_val <= 16'b0110000110100111;
            14'h235c 	:	o_val <= 16'b0110000110101001;
            14'h235d 	:	o_val <= 16'b0110000110101011;
            14'h235e 	:	o_val <= 16'b0110000110101101;
            14'h235f 	:	o_val <= 16'b0110000110101111;
            14'h2360 	:	o_val <= 16'b0110000110110001;
            14'h2361 	:	o_val <= 16'b0110000110110011;
            14'h2362 	:	o_val <= 16'b0110000110110101;
            14'h2363 	:	o_val <= 16'b0110000110110111;
            14'h2364 	:	o_val <= 16'b0110000110111001;
            14'h2365 	:	o_val <= 16'b0110000110111011;
            14'h2366 	:	o_val <= 16'b0110000110111101;
            14'h2367 	:	o_val <= 16'b0110000110111111;
            14'h2368 	:	o_val <= 16'b0110000111000001;
            14'h2369 	:	o_val <= 16'b0110000111000011;
            14'h236a 	:	o_val <= 16'b0110000111000101;
            14'h236b 	:	o_val <= 16'b0110000111000111;
            14'h236c 	:	o_val <= 16'b0110000111001001;
            14'h236d 	:	o_val <= 16'b0110000111001011;
            14'h236e 	:	o_val <= 16'b0110000111001101;
            14'h236f 	:	o_val <= 16'b0110000111001111;
            14'h2370 	:	o_val <= 16'b0110000111010001;
            14'h2371 	:	o_val <= 16'b0110000111010011;
            14'h2372 	:	o_val <= 16'b0110000111010101;
            14'h2373 	:	o_val <= 16'b0110000111010111;
            14'h2374 	:	o_val <= 16'b0110000111011001;
            14'h2375 	:	o_val <= 16'b0110000111011011;
            14'h2376 	:	o_val <= 16'b0110000111011101;
            14'h2377 	:	o_val <= 16'b0110000111011111;
            14'h2378 	:	o_val <= 16'b0110000111100001;
            14'h2379 	:	o_val <= 16'b0110000111100011;
            14'h237a 	:	o_val <= 16'b0110000111100101;
            14'h237b 	:	o_val <= 16'b0110000111100111;
            14'h237c 	:	o_val <= 16'b0110000111101001;
            14'h237d 	:	o_val <= 16'b0110000111101011;
            14'h237e 	:	o_val <= 16'b0110000111101101;
            14'h237f 	:	o_val <= 16'b0110000111101111;
            14'h2380 	:	o_val <= 16'b0110000111110010;
            14'h2381 	:	o_val <= 16'b0110000111110100;
            14'h2382 	:	o_val <= 16'b0110000111110110;
            14'h2383 	:	o_val <= 16'b0110000111111000;
            14'h2384 	:	o_val <= 16'b0110000111111010;
            14'h2385 	:	o_val <= 16'b0110000111111100;
            14'h2386 	:	o_val <= 16'b0110000111111110;
            14'h2387 	:	o_val <= 16'b0110001000000000;
            14'h2388 	:	o_val <= 16'b0110001000000010;
            14'h2389 	:	o_val <= 16'b0110001000000100;
            14'h238a 	:	o_val <= 16'b0110001000000110;
            14'h238b 	:	o_val <= 16'b0110001000001000;
            14'h238c 	:	o_val <= 16'b0110001000001010;
            14'h238d 	:	o_val <= 16'b0110001000001100;
            14'h238e 	:	o_val <= 16'b0110001000001110;
            14'h238f 	:	o_val <= 16'b0110001000010000;
            14'h2390 	:	o_val <= 16'b0110001000010010;
            14'h2391 	:	o_val <= 16'b0110001000010100;
            14'h2392 	:	o_val <= 16'b0110001000010110;
            14'h2393 	:	o_val <= 16'b0110001000011000;
            14'h2394 	:	o_val <= 16'b0110001000011010;
            14'h2395 	:	o_val <= 16'b0110001000011100;
            14'h2396 	:	o_val <= 16'b0110001000011110;
            14'h2397 	:	o_val <= 16'b0110001000100000;
            14'h2398 	:	o_val <= 16'b0110001000100010;
            14'h2399 	:	o_val <= 16'b0110001000100100;
            14'h239a 	:	o_val <= 16'b0110001000100110;
            14'h239b 	:	o_val <= 16'b0110001000101000;
            14'h239c 	:	o_val <= 16'b0110001000101010;
            14'h239d 	:	o_val <= 16'b0110001000101100;
            14'h239e 	:	o_val <= 16'b0110001000101110;
            14'h239f 	:	o_val <= 16'b0110001000110000;
            14'h23a0 	:	o_val <= 16'b0110001000110010;
            14'h23a1 	:	o_val <= 16'b0110001000110100;
            14'h23a2 	:	o_val <= 16'b0110001000110110;
            14'h23a3 	:	o_val <= 16'b0110001000111000;
            14'h23a4 	:	o_val <= 16'b0110001000111010;
            14'h23a5 	:	o_val <= 16'b0110001000111100;
            14'h23a6 	:	o_val <= 16'b0110001000111110;
            14'h23a7 	:	o_val <= 16'b0110001001000000;
            14'h23a8 	:	o_val <= 16'b0110001001000010;
            14'h23a9 	:	o_val <= 16'b0110001001000100;
            14'h23aa 	:	o_val <= 16'b0110001001000110;
            14'h23ab 	:	o_val <= 16'b0110001001001000;
            14'h23ac 	:	o_val <= 16'b0110001001001010;
            14'h23ad 	:	o_val <= 16'b0110001001001100;
            14'h23ae 	:	o_val <= 16'b0110001001001110;
            14'h23af 	:	o_val <= 16'b0110001001010000;
            14'h23b0 	:	o_val <= 16'b0110001001010010;
            14'h23b1 	:	o_val <= 16'b0110001001010100;
            14'h23b2 	:	o_val <= 16'b0110001001010110;
            14'h23b3 	:	o_val <= 16'b0110001001011000;
            14'h23b4 	:	o_val <= 16'b0110001001011010;
            14'h23b5 	:	o_val <= 16'b0110001001011100;
            14'h23b6 	:	o_val <= 16'b0110001001011110;
            14'h23b7 	:	o_val <= 16'b0110001001100000;
            14'h23b8 	:	o_val <= 16'b0110001001100010;
            14'h23b9 	:	o_val <= 16'b0110001001100100;
            14'h23ba 	:	o_val <= 16'b0110001001100110;
            14'h23bb 	:	o_val <= 16'b0110001001101000;
            14'h23bc 	:	o_val <= 16'b0110001001101010;
            14'h23bd 	:	o_val <= 16'b0110001001101100;
            14'h23be 	:	o_val <= 16'b0110001001101110;
            14'h23bf 	:	o_val <= 16'b0110001001110000;
            14'h23c0 	:	o_val <= 16'b0110001001110010;
            14'h23c1 	:	o_val <= 16'b0110001001110100;
            14'h23c2 	:	o_val <= 16'b0110001001110110;
            14'h23c3 	:	o_val <= 16'b0110001001111001;
            14'h23c4 	:	o_val <= 16'b0110001001111011;
            14'h23c5 	:	o_val <= 16'b0110001001111101;
            14'h23c6 	:	o_val <= 16'b0110001001111111;
            14'h23c7 	:	o_val <= 16'b0110001010000001;
            14'h23c8 	:	o_val <= 16'b0110001010000011;
            14'h23c9 	:	o_val <= 16'b0110001010000101;
            14'h23ca 	:	o_val <= 16'b0110001010000111;
            14'h23cb 	:	o_val <= 16'b0110001010001001;
            14'h23cc 	:	o_val <= 16'b0110001010001011;
            14'h23cd 	:	o_val <= 16'b0110001010001101;
            14'h23ce 	:	o_val <= 16'b0110001010001111;
            14'h23cf 	:	o_val <= 16'b0110001010010001;
            14'h23d0 	:	o_val <= 16'b0110001010010011;
            14'h23d1 	:	o_val <= 16'b0110001010010101;
            14'h23d2 	:	o_val <= 16'b0110001010010111;
            14'h23d3 	:	o_val <= 16'b0110001010011001;
            14'h23d4 	:	o_val <= 16'b0110001010011011;
            14'h23d5 	:	o_val <= 16'b0110001010011101;
            14'h23d6 	:	o_val <= 16'b0110001010011111;
            14'h23d7 	:	o_val <= 16'b0110001010100001;
            14'h23d8 	:	o_val <= 16'b0110001010100011;
            14'h23d9 	:	o_val <= 16'b0110001010100101;
            14'h23da 	:	o_val <= 16'b0110001010100111;
            14'h23db 	:	o_val <= 16'b0110001010101001;
            14'h23dc 	:	o_val <= 16'b0110001010101011;
            14'h23dd 	:	o_val <= 16'b0110001010101101;
            14'h23de 	:	o_val <= 16'b0110001010101111;
            14'h23df 	:	o_val <= 16'b0110001010110001;
            14'h23e0 	:	o_val <= 16'b0110001010110011;
            14'h23e1 	:	o_val <= 16'b0110001010110101;
            14'h23e2 	:	o_val <= 16'b0110001010110111;
            14'h23e3 	:	o_val <= 16'b0110001010111001;
            14'h23e4 	:	o_val <= 16'b0110001010111011;
            14'h23e5 	:	o_val <= 16'b0110001010111101;
            14'h23e6 	:	o_val <= 16'b0110001010111111;
            14'h23e7 	:	o_val <= 16'b0110001011000001;
            14'h23e8 	:	o_val <= 16'b0110001011000011;
            14'h23e9 	:	o_val <= 16'b0110001011000101;
            14'h23ea 	:	o_val <= 16'b0110001011000111;
            14'h23eb 	:	o_val <= 16'b0110001011001001;
            14'h23ec 	:	o_val <= 16'b0110001011001011;
            14'h23ed 	:	o_val <= 16'b0110001011001101;
            14'h23ee 	:	o_val <= 16'b0110001011001111;
            14'h23ef 	:	o_val <= 16'b0110001011010001;
            14'h23f0 	:	o_val <= 16'b0110001011010011;
            14'h23f1 	:	o_val <= 16'b0110001011010101;
            14'h23f2 	:	o_val <= 16'b0110001011010111;
            14'h23f3 	:	o_val <= 16'b0110001011011001;
            14'h23f4 	:	o_val <= 16'b0110001011011011;
            14'h23f5 	:	o_val <= 16'b0110001011011101;
            14'h23f6 	:	o_val <= 16'b0110001011011111;
            14'h23f7 	:	o_val <= 16'b0110001011100001;
            14'h23f8 	:	o_val <= 16'b0110001011100011;
            14'h23f9 	:	o_val <= 16'b0110001011100101;
            14'h23fa 	:	o_val <= 16'b0110001011100111;
            14'h23fb 	:	o_val <= 16'b0110001011101001;
            14'h23fc 	:	o_val <= 16'b0110001011101011;
            14'h23fd 	:	o_val <= 16'b0110001011101101;
            14'h23fe 	:	o_val <= 16'b0110001011101111;
            14'h23ff 	:	o_val <= 16'b0110001011110001;
            14'h2400 	:	o_val <= 16'b0110001011110011;
            14'h2401 	:	o_val <= 16'b0110001011110100;
            14'h2402 	:	o_val <= 16'b0110001011110110;
            14'h2403 	:	o_val <= 16'b0110001011111000;
            14'h2404 	:	o_val <= 16'b0110001011111010;
            14'h2405 	:	o_val <= 16'b0110001011111100;
            14'h2406 	:	o_val <= 16'b0110001011111110;
            14'h2407 	:	o_val <= 16'b0110001100000000;
            14'h2408 	:	o_val <= 16'b0110001100000010;
            14'h2409 	:	o_val <= 16'b0110001100000100;
            14'h240a 	:	o_val <= 16'b0110001100000110;
            14'h240b 	:	o_val <= 16'b0110001100001000;
            14'h240c 	:	o_val <= 16'b0110001100001010;
            14'h240d 	:	o_val <= 16'b0110001100001100;
            14'h240e 	:	o_val <= 16'b0110001100001110;
            14'h240f 	:	o_val <= 16'b0110001100010000;
            14'h2410 	:	o_val <= 16'b0110001100010010;
            14'h2411 	:	o_val <= 16'b0110001100010100;
            14'h2412 	:	o_val <= 16'b0110001100010110;
            14'h2413 	:	o_val <= 16'b0110001100011000;
            14'h2414 	:	o_val <= 16'b0110001100011010;
            14'h2415 	:	o_val <= 16'b0110001100011100;
            14'h2416 	:	o_val <= 16'b0110001100011110;
            14'h2417 	:	o_val <= 16'b0110001100100000;
            14'h2418 	:	o_val <= 16'b0110001100100010;
            14'h2419 	:	o_val <= 16'b0110001100100100;
            14'h241a 	:	o_val <= 16'b0110001100100110;
            14'h241b 	:	o_val <= 16'b0110001100101000;
            14'h241c 	:	o_val <= 16'b0110001100101010;
            14'h241d 	:	o_val <= 16'b0110001100101100;
            14'h241e 	:	o_val <= 16'b0110001100101110;
            14'h241f 	:	o_val <= 16'b0110001100110000;
            14'h2420 	:	o_val <= 16'b0110001100110010;
            14'h2421 	:	o_val <= 16'b0110001100110100;
            14'h2422 	:	o_val <= 16'b0110001100110110;
            14'h2423 	:	o_val <= 16'b0110001100111000;
            14'h2424 	:	o_val <= 16'b0110001100111010;
            14'h2425 	:	o_val <= 16'b0110001100111100;
            14'h2426 	:	o_val <= 16'b0110001100111110;
            14'h2427 	:	o_val <= 16'b0110001101000000;
            14'h2428 	:	o_val <= 16'b0110001101000010;
            14'h2429 	:	o_val <= 16'b0110001101000100;
            14'h242a 	:	o_val <= 16'b0110001101000110;
            14'h242b 	:	o_val <= 16'b0110001101001000;
            14'h242c 	:	o_val <= 16'b0110001101001010;
            14'h242d 	:	o_val <= 16'b0110001101001100;
            14'h242e 	:	o_val <= 16'b0110001101001110;
            14'h242f 	:	o_val <= 16'b0110001101010000;
            14'h2430 	:	o_val <= 16'b0110001101010010;
            14'h2431 	:	o_val <= 16'b0110001101010100;
            14'h2432 	:	o_val <= 16'b0110001101010110;
            14'h2433 	:	o_val <= 16'b0110001101011000;
            14'h2434 	:	o_val <= 16'b0110001101011010;
            14'h2435 	:	o_val <= 16'b0110001101011100;
            14'h2436 	:	o_val <= 16'b0110001101011110;
            14'h2437 	:	o_val <= 16'b0110001101100000;
            14'h2438 	:	o_val <= 16'b0110001101100010;
            14'h2439 	:	o_val <= 16'b0110001101100100;
            14'h243a 	:	o_val <= 16'b0110001101100110;
            14'h243b 	:	o_val <= 16'b0110001101101000;
            14'h243c 	:	o_val <= 16'b0110001101101010;
            14'h243d 	:	o_val <= 16'b0110001101101100;
            14'h243e 	:	o_val <= 16'b0110001101101110;
            14'h243f 	:	o_val <= 16'b0110001101110000;
            14'h2440 	:	o_val <= 16'b0110001101110010;
            14'h2441 	:	o_val <= 16'b0110001101110100;
            14'h2442 	:	o_val <= 16'b0110001101110110;
            14'h2443 	:	o_val <= 16'b0110001101111000;
            14'h2444 	:	o_val <= 16'b0110001101111001;
            14'h2445 	:	o_val <= 16'b0110001101111011;
            14'h2446 	:	o_val <= 16'b0110001101111101;
            14'h2447 	:	o_val <= 16'b0110001101111111;
            14'h2448 	:	o_val <= 16'b0110001110000001;
            14'h2449 	:	o_val <= 16'b0110001110000011;
            14'h244a 	:	o_val <= 16'b0110001110000101;
            14'h244b 	:	o_val <= 16'b0110001110000111;
            14'h244c 	:	o_val <= 16'b0110001110001001;
            14'h244d 	:	o_val <= 16'b0110001110001011;
            14'h244e 	:	o_val <= 16'b0110001110001101;
            14'h244f 	:	o_val <= 16'b0110001110001111;
            14'h2450 	:	o_val <= 16'b0110001110010001;
            14'h2451 	:	o_val <= 16'b0110001110010011;
            14'h2452 	:	o_val <= 16'b0110001110010101;
            14'h2453 	:	o_val <= 16'b0110001110010111;
            14'h2454 	:	o_val <= 16'b0110001110011001;
            14'h2455 	:	o_val <= 16'b0110001110011011;
            14'h2456 	:	o_val <= 16'b0110001110011101;
            14'h2457 	:	o_val <= 16'b0110001110011111;
            14'h2458 	:	o_val <= 16'b0110001110100001;
            14'h2459 	:	o_val <= 16'b0110001110100011;
            14'h245a 	:	o_val <= 16'b0110001110100101;
            14'h245b 	:	o_val <= 16'b0110001110100111;
            14'h245c 	:	o_val <= 16'b0110001110101001;
            14'h245d 	:	o_val <= 16'b0110001110101011;
            14'h245e 	:	o_val <= 16'b0110001110101101;
            14'h245f 	:	o_val <= 16'b0110001110101111;
            14'h2460 	:	o_val <= 16'b0110001110110001;
            14'h2461 	:	o_val <= 16'b0110001110110011;
            14'h2462 	:	o_val <= 16'b0110001110110101;
            14'h2463 	:	o_val <= 16'b0110001110110111;
            14'h2464 	:	o_val <= 16'b0110001110111001;
            14'h2465 	:	o_val <= 16'b0110001110111011;
            14'h2466 	:	o_val <= 16'b0110001110111101;
            14'h2467 	:	o_val <= 16'b0110001110111111;
            14'h2468 	:	o_val <= 16'b0110001111000001;
            14'h2469 	:	o_val <= 16'b0110001111000010;
            14'h246a 	:	o_val <= 16'b0110001111000100;
            14'h246b 	:	o_val <= 16'b0110001111000110;
            14'h246c 	:	o_val <= 16'b0110001111001000;
            14'h246d 	:	o_val <= 16'b0110001111001010;
            14'h246e 	:	o_val <= 16'b0110001111001100;
            14'h246f 	:	o_val <= 16'b0110001111001110;
            14'h2470 	:	o_val <= 16'b0110001111010000;
            14'h2471 	:	o_val <= 16'b0110001111010010;
            14'h2472 	:	o_val <= 16'b0110001111010100;
            14'h2473 	:	o_val <= 16'b0110001111010110;
            14'h2474 	:	o_val <= 16'b0110001111011000;
            14'h2475 	:	o_val <= 16'b0110001111011010;
            14'h2476 	:	o_val <= 16'b0110001111011100;
            14'h2477 	:	o_val <= 16'b0110001111011110;
            14'h2478 	:	o_val <= 16'b0110001111100000;
            14'h2479 	:	o_val <= 16'b0110001111100010;
            14'h247a 	:	o_val <= 16'b0110001111100100;
            14'h247b 	:	o_val <= 16'b0110001111100110;
            14'h247c 	:	o_val <= 16'b0110001111101000;
            14'h247d 	:	o_val <= 16'b0110001111101010;
            14'h247e 	:	o_val <= 16'b0110001111101100;
            14'h247f 	:	o_val <= 16'b0110001111101110;
            14'h2480 	:	o_val <= 16'b0110001111110000;
            14'h2481 	:	o_val <= 16'b0110001111110010;
            14'h2482 	:	o_val <= 16'b0110001111110100;
            14'h2483 	:	o_val <= 16'b0110001111110110;
            14'h2484 	:	o_val <= 16'b0110001111111000;
            14'h2485 	:	o_val <= 16'b0110001111111001;
            14'h2486 	:	o_val <= 16'b0110001111111011;
            14'h2487 	:	o_val <= 16'b0110001111111101;
            14'h2488 	:	o_val <= 16'b0110001111111111;
            14'h2489 	:	o_val <= 16'b0110010000000001;
            14'h248a 	:	o_val <= 16'b0110010000000011;
            14'h248b 	:	o_val <= 16'b0110010000000101;
            14'h248c 	:	o_val <= 16'b0110010000000111;
            14'h248d 	:	o_val <= 16'b0110010000001001;
            14'h248e 	:	o_val <= 16'b0110010000001011;
            14'h248f 	:	o_val <= 16'b0110010000001101;
            14'h2490 	:	o_val <= 16'b0110010000001111;
            14'h2491 	:	o_val <= 16'b0110010000010001;
            14'h2492 	:	o_val <= 16'b0110010000010011;
            14'h2493 	:	o_val <= 16'b0110010000010101;
            14'h2494 	:	o_val <= 16'b0110010000010111;
            14'h2495 	:	o_val <= 16'b0110010000011001;
            14'h2496 	:	o_val <= 16'b0110010000011011;
            14'h2497 	:	o_val <= 16'b0110010000011101;
            14'h2498 	:	o_val <= 16'b0110010000011111;
            14'h2499 	:	o_val <= 16'b0110010000100001;
            14'h249a 	:	o_val <= 16'b0110010000100011;
            14'h249b 	:	o_val <= 16'b0110010000100101;
            14'h249c 	:	o_val <= 16'b0110010000100111;
            14'h249d 	:	o_val <= 16'b0110010000101001;
            14'h249e 	:	o_val <= 16'b0110010000101010;
            14'h249f 	:	o_val <= 16'b0110010000101100;
            14'h24a0 	:	o_val <= 16'b0110010000101110;
            14'h24a1 	:	o_val <= 16'b0110010000110000;
            14'h24a2 	:	o_val <= 16'b0110010000110010;
            14'h24a3 	:	o_val <= 16'b0110010000110100;
            14'h24a4 	:	o_val <= 16'b0110010000110110;
            14'h24a5 	:	o_val <= 16'b0110010000111000;
            14'h24a6 	:	o_val <= 16'b0110010000111010;
            14'h24a7 	:	o_val <= 16'b0110010000111100;
            14'h24a8 	:	o_val <= 16'b0110010000111110;
            14'h24a9 	:	o_val <= 16'b0110010001000000;
            14'h24aa 	:	o_val <= 16'b0110010001000010;
            14'h24ab 	:	o_val <= 16'b0110010001000100;
            14'h24ac 	:	o_val <= 16'b0110010001000110;
            14'h24ad 	:	o_val <= 16'b0110010001001000;
            14'h24ae 	:	o_val <= 16'b0110010001001010;
            14'h24af 	:	o_val <= 16'b0110010001001100;
            14'h24b0 	:	o_val <= 16'b0110010001001110;
            14'h24b1 	:	o_val <= 16'b0110010001010000;
            14'h24b2 	:	o_val <= 16'b0110010001010010;
            14'h24b3 	:	o_val <= 16'b0110010001010011;
            14'h24b4 	:	o_val <= 16'b0110010001010101;
            14'h24b5 	:	o_val <= 16'b0110010001010111;
            14'h24b6 	:	o_val <= 16'b0110010001011001;
            14'h24b7 	:	o_val <= 16'b0110010001011011;
            14'h24b8 	:	o_val <= 16'b0110010001011101;
            14'h24b9 	:	o_val <= 16'b0110010001011111;
            14'h24ba 	:	o_val <= 16'b0110010001100001;
            14'h24bb 	:	o_val <= 16'b0110010001100011;
            14'h24bc 	:	o_val <= 16'b0110010001100101;
            14'h24bd 	:	o_val <= 16'b0110010001100111;
            14'h24be 	:	o_val <= 16'b0110010001101001;
            14'h24bf 	:	o_val <= 16'b0110010001101011;
            14'h24c0 	:	o_val <= 16'b0110010001101101;
            14'h24c1 	:	o_val <= 16'b0110010001101111;
            14'h24c2 	:	o_val <= 16'b0110010001110001;
            14'h24c3 	:	o_val <= 16'b0110010001110011;
            14'h24c4 	:	o_val <= 16'b0110010001110101;
            14'h24c5 	:	o_val <= 16'b0110010001110111;
            14'h24c6 	:	o_val <= 16'b0110010001111001;
            14'h24c7 	:	o_val <= 16'b0110010001111010;
            14'h24c8 	:	o_val <= 16'b0110010001111100;
            14'h24c9 	:	o_val <= 16'b0110010001111110;
            14'h24ca 	:	o_val <= 16'b0110010010000000;
            14'h24cb 	:	o_val <= 16'b0110010010000010;
            14'h24cc 	:	o_val <= 16'b0110010010000100;
            14'h24cd 	:	o_val <= 16'b0110010010000110;
            14'h24ce 	:	o_val <= 16'b0110010010001000;
            14'h24cf 	:	o_val <= 16'b0110010010001010;
            14'h24d0 	:	o_val <= 16'b0110010010001100;
            14'h24d1 	:	o_val <= 16'b0110010010001110;
            14'h24d2 	:	o_val <= 16'b0110010010010000;
            14'h24d3 	:	o_val <= 16'b0110010010010010;
            14'h24d4 	:	o_val <= 16'b0110010010010100;
            14'h24d5 	:	o_val <= 16'b0110010010010110;
            14'h24d6 	:	o_val <= 16'b0110010010011000;
            14'h24d7 	:	o_val <= 16'b0110010010011010;
            14'h24d8 	:	o_val <= 16'b0110010010011100;
            14'h24d9 	:	o_val <= 16'b0110010010011101;
            14'h24da 	:	o_val <= 16'b0110010010011111;
            14'h24db 	:	o_val <= 16'b0110010010100001;
            14'h24dc 	:	o_val <= 16'b0110010010100011;
            14'h24dd 	:	o_val <= 16'b0110010010100101;
            14'h24de 	:	o_val <= 16'b0110010010100111;
            14'h24df 	:	o_val <= 16'b0110010010101001;
            14'h24e0 	:	o_val <= 16'b0110010010101011;
            14'h24e1 	:	o_val <= 16'b0110010010101101;
            14'h24e2 	:	o_val <= 16'b0110010010101111;
            14'h24e3 	:	o_val <= 16'b0110010010110001;
            14'h24e4 	:	o_val <= 16'b0110010010110011;
            14'h24e5 	:	o_val <= 16'b0110010010110101;
            14'h24e6 	:	o_val <= 16'b0110010010110111;
            14'h24e7 	:	o_val <= 16'b0110010010111001;
            14'h24e8 	:	o_val <= 16'b0110010010111011;
            14'h24e9 	:	o_val <= 16'b0110010010111100;
            14'h24ea 	:	o_val <= 16'b0110010010111110;
            14'h24eb 	:	o_val <= 16'b0110010011000000;
            14'h24ec 	:	o_val <= 16'b0110010011000010;
            14'h24ed 	:	o_val <= 16'b0110010011000100;
            14'h24ee 	:	o_val <= 16'b0110010011000110;
            14'h24ef 	:	o_val <= 16'b0110010011001000;
            14'h24f0 	:	o_val <= 16'b0110010011001010;
            14'h24f1 	:	o_val <= 16'b0110010011001100;
            14'h24f2 	:	o_val <= 16'b0110010011001110;
            14'h24f3 	:	o_val <= 16'b0110010011010000;
            14'h24f4 	:	o_val <= 16'b0110010011010010;
            14'h24f5 	:	o_val <= 16'b0110010011010100;
            14'h24f6 	:	o_val <= 16'b0110010011010110;
            14'h24f7 	:	o_val <= 16'b0110010011011000;
            14'h24f8 	:	o_val <= 16'b0110010011011010;
            14'h24f9 	:	o_val <= 16'b0110010011011011;
            14'h24fa 	:	o_val <= 16'b0110010011011101;
            14'h24fb 	:	o_val <= 16'b0110010011011111;
            14'h24fc 	:	o_val <= 16'b0110010011100001;
            14'h24fd 	:	o_val <= 16'b0110010011100011;
            14'h24fe 	:	o_val <= 16'b0110010011100101;
            14'h24ff 	:	o_val <= 16'b0110010011100111;
            14'h2500 	:	o_val <= 16'b0110010011101001;
            14'h2501 	:	o_val <= 16'b0110010011101011;
            14'h2502 	:	o_val <= 16'b0110010011101101;
            14'h2503 	:	o_val <= 16'b0110010011101111;
            14'h2504 	:	o_val <= 16'b0110010011110001;
            14'h2505 	:	o_val <= 16'b0110010011110011;
            14'h2506 	:	o_val <= 16'b0110010011110101;
            14'h2507 	:	o_val <= 16'b0110010011110111;
            14'h2508 	:	o_val <= 16'b0110010011111000;
            14'h2509 	:	o_val <= 16'b0110010011111010;
            14'h250a 	:	o_val <= 16'b0110010011111100;
            14'h250b 	:	o_val <= 16'b0110010011111110;
            14'h250c 	:	o_val <= 16'b0110010100000000;
            14'h250d 	:	o_val <= 16'b0110010100000010;
            14'h250e 	:	o_val <= 16'b0110010100000100;
            14'h250f 	:	o_val <= 16'b0110010100000110;
            14'h2510 	:	o_val <= 16'b0110010100001000;
            14'h2511 	:	o_val <= 16'b0110010100001010;
            14'h2512 	:	o_val <= 16'b0110010100001100;
            14'h2513 	:	o_val <= 16'b0110010100001110;
            14'h2514 	:	o_val <= 16'b0110010100010000;
            14'h2515 	:	o_val <= 16'b0110010100010010;
            14'h2516 	:	o_val <= 16'b0110010100010011;
            14'h2517 	:	o_val <= 16'b0110010100010101;
            14'h2518 	:	o_val <= 16'b0110010100010111;
            14'h2519 	:	o_val <= 16'b0110010100011001;
            14'h251a 	:	o_val <= 16'b0110010100011011;
            14'h251b 	:	o_val <= 16'b0110010100011101;
            14'h251c 	:	o_val <= 16'b0110010100011111;
            14'h251d 	:	o_val <= 16'b0110010100100001;
            14'h251e 	:	o_val <= 16'b0110010100100011;
            14'h251f 	:	o_val <= 16'b0110010100100101;
            14'h2520 	:	o_val <= 16'b0110010100100111;
            14'h2521 	:	o_val <= 16'b0110010100101001;
            14'h2522 	:	o_val <= 16'b0110010100101011;
            14'h2523 	:	o_val <= 16'b0110010100101101;
            14'h2524 	:	o_val <= 16'b0110010100101110;
            14'h2525 	:	o_val <= 16'b0110010100110000;
            14'h2526 	:	o_val <= 16'b0110010100110010;
            14'h2527 	:	o_val <= 16'b0110010100110100;
            14'h2528 	:	o_val <= 16'b0110010100110110;
            14'h2529 	:	o_val <= 16'b0110010100111000;
            14'h252a 	:	o_val <= 16'b0110010100111010;
            14'h252b 	:	o_val <= 16'b0110010100111100;
            14'h252c 	:	o_val <= 16'b0110010100111110;
            14'h252d 	:	o_val <= 16'b0110010101000000;
            14'h252e 	:	o_val <= 16'b0110010101000010;
            14'h252f 	:	o_val <= 16'b0110010101000100;
            14'h2530 	:	o_val <= 16'b0110010101000101;
            14'h2531 	:	o_val <= 16'b0110010101000111;
            14'h2532 	:	o_val <= 16'b0110010101001001;
            14'h2533 	:	o_val <= 16'b0110010101001011;
            14'h2534 	:	o_val <= 16'b0110010101001101;
            14'h2535 	:	o_val <= 16'b0110010101001111;
            14'h2536 	:	o_val <= 16'b0110010101010001;
            14'h2537 	:	o_val <= 16'b0110010101010011;
            14'h2538 	:	o_val <= 16'b0110010101010101;
            14'h2539 	:	o_val <= 16'b0110010101010111;
            14'h253a 	:	o_val <= 16'b0110010101011001;
            14'h253b 	:	o_val <= 16'b0110010101011011;
            14'h253c 	:	o_val <= 16'b0110010101011101;
            14'h253d 	:	o_val <= 16'b0110010101011110;
            14'h253e 	:	o_val <= 16'b0110010101100000;
            14'h253f 	:	o_val <= 16'b0110010101100010;
            14'h2540 	:	o_val <= 16'b0110010101100100;
            14'h2541 	:	o_val <= 16'b0110010101100110;
            14'h2542 	:	o_val <= 16'b0110010101101000;
            14'h2543 	:	o_val <= 16'b0110010101101010;
            14'h2544 	:	o_val <= 16'b0110010101101100;
            14'h2545 	:	o_val <= 16'b0110010101101110;
            14'h2546 	:	o_val <= 16'b0110010101110000;
            14'h2547 	:	o_val <= 16'b0110010101110010;
            14'h2548 	:	o_val <= 16'b0110010101110100;
            14'h2549 	:	o_val <= 16'b0110010101110101;
            14'h254a 	:	o_val <= 16'b0110010101110111;
            14'h254b 	:	o_val <= 16'b0110010101111001;
            14'h254c 	:	o_val <= 16'b0110010101111011;
            14'h254d 	:	o_val <= 16'b0110010101111101;
            14'h254e 	:	o_val <= 16'b0110010101111111;
            14'h254f 	:	o_val <= 16'b0110010110000001;
            14'h2550 	:	o_val <= 16'b0110010110000011;
            14'h2551 	:	o_val <= 16'b0110010110000101;
            14'h2552 	:	o_val <= 16'b0110010110000111;
            14'h2553 	:	o_val <= 16'b0110010110001001;
            14'h2554 	:	o_val <= 16'b0110010110001011;
            14'h2555 	:	o_val <= 16'b0110010110001100;
            14'h2556 	:	o_val <= 16'b0110010110001110;
            14'h2557 	:	o_val <= 16'b0110010110010000;
            14'h2558 	:	o_val <= 16'b0110010110010010;
            14'h2559 	:	o_val <= 16'b0110010110010100;
            14'h255a 	:	o_val <= 16'b0110010110010110;
            14'h255b 	:	o_val <= 16'b0110010110011000;
            14'h255c 	:	o_val <= 16'b0110010110011010;
            14'h255d 	:	o_val <= 16'b0110010110011100;
            14'h255e 	:	o_val <= 16'b0110010110011110;
            14'h255f 	:	o_val <= 16'b0110010110100000;
            14'h2560 	:	o_val <= 16'b0110010110100001;
            14'h2561 	:	o_val <= 16'b0110010110100011;
            14'h2562 	:	o_val <= 16'b0110010110100101;
            14'h2563 	:	o_val <= 16'b0110010110100111;
            14'h2564 	:	o_val <= 16'b0110010110101001;
            14'h2565 	:	o_val <= 16'b0110010110101011;
            14'h2566 	:	o_val <= 16'b0110010110101101;
            14'h2567 	:	o_val <= 16'b0110010110101111;
            14'h2568 	:	o_val <= 16'b0110010110110001;
            14'h2569 	:	o_val <= 16'b0110010110110011;
            14'h256a 	:	o_val <= 16'b0110010110110101;
            14'h256b 	:	o_val <= 16'b0110010110110110;
            14'h256c 	:	o_val <= 16'b0110010110111000;
            14'h256d 	:	o_val <= 16'b0110010110111010;
            14'h256e 	:	o_val <= 16'b0110010110111100;
            14'h256f 	:	o_val <= 16'b0110010110111110;
            14'h2570 	:	o_val <= 16'b0110010111000000;
            14'h2571 	:	o_val <= 16'b0110010111000010;
            14'h2572 	:	o_val <= 16'b0110010111000100;
            14'h2573 	:	o_val <= 16'b0110010111000110;
            14'h2574 	:	o_val <= 16'b0110010111001000;
            14'h2575 	:	o_val <= 16'b0110010111001001;
            14'h2576 	:	o_val <= 16'b0110010111001011;
            14'h2577 	:	o_val <= 16'b0110010111001101;
            14'h2578 	:	o_val <= 16'b0110010111001111;
            14'h2579 	:	o_val <= 16'b0110010111010001;
            14'h257a 	:	o_val <= 16'b0110010111010011;
            14'h257b 	:	o_val <= 16'b0110010111010101;
            14'h257c 	:	o_val <= 16'b0110010111010111;
            14'h257d 	:	o_val <= 16'b0110010111011001;
            14'h257e 	:	o_val <= 16'b0110010111011011;
            14'h257f 	:	o_val <= 16'b0110010111011101;
            14'h2580 	:	o_val <= 16'b0110010111011110;
            14'h2581 	:	o_val <= 16'b0110010111100000;
            14'h2582 	:	o_val <= 16'b0110010111100010;
            14'h2583 	:	o_val <= 16'b0110010111100100;
            14'h2584 	:	o_val <= 16'b0110010111100110;
            14'h2585 	:	o_val <= 16'b0110010111101000;
            14'h2586 	:	o_val <= 16'b0110010111101010;
            14'h2587 	:	o_val <= 16'b0110010111101100;
            14'h2588 	:	o_val <= 16'b0110010111101110;
            14'h2589 	:	o_val <= 16'b0110010111110000;
            14'h258a 	:	o_val <= 16'b0110010111110001;
            14'h258b 	:	o_val <= 16'b0110010111110011;
            14'h258c 	:	o_val <= 16'b0110010111110101;
            14'h258d 	:	o_val <= 16'b0110010111110111;
            14'h258e 	:	o_val <= 16'b0110010111111001;
            14'h258f 	:	o_val <= 16'b0110010111111011;
            14'h2590 	:	o_val <= 16'b0110010111111101;
            14'h2591 	:	o_val <= 16'b0110010111111111;
            14'h2592 	:	o_val <= 16'b0110011000000001;
            14'h2593 	:	o_val <= 16'b0110011000000011;
            14'h2594 	:	o_val <= 16'b0110011000000100;
            14'h2595 	:	o_val <= 16'b0110011000000110;
            14'h2596 	:	o_val <= 16'b0110011000001000;
            14'h2597 	:	o_val <= 16'b0110011000001010;
            14'h2598 	:	o_val <= 16'b0110011000001100;
            14'h2599 	:	o_val <= 16'b0110011000001110;
            14'h259a 	:	o_val <= 16'b0110011000010000;
            14'h259b 	:	o_val <= 16'b0110011000010010;
            14'h259c 	:	o_val <= 16'b0110011000010100;
            14'h259d 	:	o_val <= 16'b0110011000010101;
            14'h259e 	:	o_val <= 16'b0110011000010111;
            14'h259f 	:	o_val <= 16'b0110011000011001;
            14'h25a0 	:	o_val <= 16'b0110011000011011;
            14'h25a1 	:	o_val <= 16'b0110011000011101;
            14'h25a2 	:	o_val <= 16'b0110011000011111;
            14'h25a3 	:	o_val <= 16'b0110011000100001;
            14'h25a4 	:	o_val <= 16'b0110011000100011;
            14'h25a5 	:	o_val <= 16'b0110011000100101;
            14'h25a6 	:	o_val <= 16'b0110011000100111;
            14'h25a7 	:	o_val <= 16'b0110011000101000;
            14'h25a8 	:	o_val <= 16'b0110011000101010;
            14'h25a9 	:	o_val <= 16'b0110011000101100;
            14'h25aa 	:	o_val <= 16'b0110011000101110;
            14'h25ab 	:	o_val <= 16'b0110011000110000;
            14'h25ac 	:	o_val <= 16'b0110011000110010;
            14'h25ad 	:	o_val <= 16'b0110011000110100;
            14'h25ae 	:	o_val <= 16'b0110011000110110;
            14'h25af 	:	o_val <= 16'b0110011000111000;
            14'h25b0 	:	o_val <= 16'b0110011000111001;
            14'h25b1 	:	o_val <= 16'b0110011000111011;
            14'h25b2 	:	o_val <= 16'b0110011000111101;
            14'h25b3 	:	o_val <= 16'b0110011000111111;
            14'h25b4 	:	o_val <= 16'b0110011001000001;
            14'h25b5 	:	o_val <= 16'b0110011001000011;
            14'h25b6 	:	o_val <= 16'b0110011001000101;
            14'h25b7 	:	o_val <= 16'b0110011001000111;
            14'h25b8 	:	o_val <= 16'b0110011001001001;
            14'h25b9 	:	o_val <= 16'b0110011001001010;
            14'h25ba 	:	o_val <= 16'b0110011001001100;
            14'h25bb 	:	o_val <= 16'b0110011001001110;
            14'h25bc 	:	o_val <= 16'b0110011001010000;
            14'h25bd 	:	o_val <= 16'b0110011001010010;
            14'h25be 	:	o_val <= 16'b0110011001010100;
            14'h25bf 	:	o_val <= 16'b0110011001010110;
            14'h25c0 	:	o_val <= 16'b0110011001011000;
            14'h25c1 	:	o_val <= 16'b0110011001011010;
            14'h25c2 	:	o_val <= 16'b0110011001011011;
            14'h25c3 	:	o_val <= 16'b0110011001011101;
            14'h25c4 	:	o_val <= 16'b0110011001011111;
            14'h25c5 	:	o_val <= 16'b0110011001100001;
            14'h25c6 	:	o_val <= 16'b0110011001100011;
            14'h25c7 	:	o_val <= 16'b0110011001100101;
            14'h25c8 	:	o_val <= 16'b0110011001100111;
            14'h25c9 	:	o_val <= 16'b0110011001101001;
            14'h25ca 	:	o_val <= 16'b0110011001101011;
            14'h25cb 	:	o_val <= 16'b0110011001101100;
            14'h25cc 	:	o_val <= 16'b0110011001101110;
            14'h25cd 	:	o_val <= 16'b0110011001110000;
            14'h25ce 	:	o_val <= 16'b0110011001110010;
            14'h25cf 	:	o_val <= 16'b0110011001110100;
            14'h25d0 	:	o_val <= 16'b0110011001110110;
            14'h25d1 	:	o_val <= 16'b0110011001111000;
            14'h25d2 	:	o_val <= 16'b0110011001111010;
            14'h25d3 	:	o_val <= 16'b0110011001111011;
            14'h25d4 	:	o_val <= 16'b0110011001111101;
            14'h25d5 	:	o_val <= 16'b0110011001111111;
            14'h25d6 	:	o_val <= 16'b0110011010000001;
            14'h25d7 	:	o_val <= 16'b0110011010000011;
            14'h25d8 	:	o_val <= 16'b0110011010000101;
            14'h25d9 	:	o_val <= 16'b0110011010000111;
            14'h25da 	:	o_val <= 16'b0110011010001001;
            14'h25db 	:	o_val <= 16'b0110011010001011;
            14'h25dc 	:	o_val <= 16'b0110011010001100;
            14'h25dd 	:	o_val <= 16'b0110011010001110;
            14'h25de 	:	o_val <= 16'b0110011010010000;
            14'h25df 	:	o_val <= 16'b0110011010010010;
            14'h25e0 	:	o_val <= 16'b0110011010010100;
            14'h25e1 	:	o_val <= 16'b0110011010010110;
            14'h25e2 	:	o_val <= 16'b0110011010011000;
            14'h25e3 	:	o_val <= 16'b0110011010011010;
            14'h25e4 	:	o_val <= 16'b0110011010011011;
            14'h25e5 	:	o_val <= 16'b0110011010011101;
            14'h25e6 	:	o_val <= 16'b0110011010011111;
            14'h25e7 	:	o_val <= 16'b0110011010100001;
            14'h25e8 	:	o_val <= 16'b0110011010100011;
            14'h25e9 	:	o_val <= 16'b0110011010100101;
            14'h25ea 	:	o_val <= 16'b0110011010100111;
            14'h25eb 	:	o_val <= 16'b0110011010101001;
            14'h25ec 	:	o_val <= 16'b0110011010101010;
            14'h25ed 	:	o_val <= 16'b0110011010101100;
            14'h25ee 	:	o_val <= 16'b0110011010101110;
            14'h25ef 	:	o_val <= 16'b0110011010110000;
            14'h25f0 	:	o_val <= 16'b0110011010110010;
            14'h25f1 	:	o_val <= 16'b0110011010110100;
            14'h25f2 	:	o_val <= 16'b0110011010110110;
            14'h25f3 	:	o_val <= 16'b0110011010111000;
            14'h25f4 	:	o_val <= 16'b0110011010111001;
            14'h25f5 	:	o_val <= 16'b0110011010111011;
            14'h25f6 	:	o_val <= 16'b0110011010111101;
            14'h25f7 	:	o_val <= 16'b0110011010111111;
            14'h25f8 	:	o_val <= 16'b0110011011000001;
            14'h25f9 	:	o_val <= 16'b0110011011000011;
            14'h25fa 	:	o_val <= 16'b0110011011000101;
            14'h25fb 	:	o_val <= 16'b0110011011000111;
            14'h25fc 	:	o_val <= 16'b0110011011001000;
            14'h25fd 	:	o_val <= 16'b0110011011001010;
            14'h25fe 	:	o_val <= 16'b0110011011001100;
            14'h25ff 	:	o_val <= 16'b0110011011001110;
            14'h2600 	:	o_val <= 16'b0110011011010000;
            14'h2601 	:	o_val <= 16'b0110011011010010;
            14'h2602 	:	o_val <= 16'b0110011011010100;
            14'h2603 	:	o_val <= 16'b0110011011010110;
            14'h2604 	:	o_val <= 16'b0110011011010111;
            14'h2605 	:	o_val <= 16'b0110011011011001;
            14'h2606 	:	o_val <= 16'b0110011011011011;
            14'h2607 	:	o_val <= 16'b0110011011011101;
            14'h2608 	:	o_val <= 16'b0110011011011111;
            14'h2609 	:	o_val <= 16'b0110011011100001;
            14'h260a 	:	o_val <= 16'b0110011011100011;
            14'h260b 	:	o_val <= 16'b0110011011100101;
            14'h260c 	:	o_val <= 16'b0110011011100110;
            14'h260d 	:	o_val <= 16'b0110011011101000;
            14'h260e 	:	o_val <= 16'b0110011011101010;
            14'h260f 	:	o_val <= 16'b0110011011101100;
            14'h2610 	:	o_val <= 16'b0110011011101110;
            14'h2611 	:	o_val <= 16'b0110011011110000;
            14'h2612 	:	o_val <= 16'b0110011011110010;
            14'h2613 	:	o_val <= 16'b0110011011110011;
            14'h2614 	:	o_val <= 16'b0110011011110101;
            14'h2615 	:	o_val <= 16'b0110011011110111;
            14'h2616 	:	o_val <= 16'b0110011011111001;
            14'h2617 	:	o_val <= 16'b0110011011111011;
            14'h2618 	:	o_val <= 16'b0110011011111101;
            14'h2619 	:	o_val <= 16'b0110011011111111;
            14'h261a 	:	o_val <= 16'b0110011100000001;
            14'h261b 	:	o_val <= 16'b0110011100000010;
            14'h261c 	:	o_val <= 16'b0110011100000100;
            14'h261d 	:	o_val <= 16'b0110011100000110;
            14'h261e 	:	o_val <= 16'b0110011100001000;
            14'h261f 	:	o_val <= 16'b0110011100001010;
            14'h2620 	:	o_val <= 16'b0110011100001100;
            14'h2621 	:	o_val <= 16'b0110011100001110;
            14'h2622 	:	o_val <= 16'b0110011100001111;
            14'h2623 	:	o_val <= 16'b0110011100010001;
            14'h2624 	:	o_val <= 16'b0110011100010011;
            14'h2625 	:	o_val <= 16'b0110011100010101;
            14'h2626 	:	o_val <= 16'b0110011100010111;
            14'h2627 	:	o_val <= 16'b0110011100011001;
            14'h2628 	:	o_val <= 16'b0110011100011011;
            14'h2629 	:	o_val <= 16'b0110011100011100;
            14'h262a 	:	o_val <= 16'b0110011100011110;
            14'h262b 	:	o_val <= 16'b0110011100100000;
            14'h262c 	:	o_val <= 16'b0110011100100010;
            14'h262d 	:	o_val <= 16'b0110011100100100;
            14'h262e 	:	o_val <= 16'b0110011100100110;
            14'h262f 	:	o_val <= 16'b0110011100101000;
            14'h2630 	:	o_val <= 16'b0110011100101001;
            14'h2631 	:	o_val <= 16'b0110011100101011;
            14'h2632 	:	o_val <= 16'b0110011100101101;
            14'h2633 	:	o_val <= 16'b0110011100101111;
            14'h2634 	:	o_val <= 16'b0110011100110001;
            14'h2635 	:	o_val <= 16'b0110011100110011;
            14'h2636 	:	o_val <= 16'b0110011100110101;
            14'h2637 	:	o_val <= 16'b0110011100110110;
            14'h2638 	:	o_val <= 16'b0110011100111000;
            14'h2639 	:	o_val <= 16'b0110011100111010;
            14'h263a 	:	o_val <= 16'b0110011100111100;
            14'h263b 	:	o_val <= 16'b0110011100111110;
            14'h263c 	:	o_val <= 16'b0110011101000000;
            14'h263d 	:	o_val <= 16'b0110011101000010;
            14'h263e 	:	o_val <= 16'b0110011101000011;
            14'h263f 	:	o_val <= 16'b0110011101000101;
            14'h2640 	:	o_val <= 16'b0110011101000111;
            14'h2641 	:	o_val <= 16'b0110011101001001;
            14'h2642 	:	o_val <= 16'b0110011101001011;
            14'h2643 	:	o_val <= 16'b0110011101001101;
            14'h2644 	:	o_val <= 16'b0110011101001111;
            14'h2645 	:	o_val <= 16'b0110011101010000;
            14'h2646 	:	o_val <= 16'b0110011101010010;
            14'h2647 	:	o_val <= 16'b0110011101010100;
            14'h2648 	:	o_val <= 16'b0110011101010110;
            14'h2649 	:	o_val <= 16'b0110011101011000;
            14'h264a 	:	o_val <= 16'b0110011101011010;
            14'h264b 	:	o_val <= 16'b0110011101011100;
            14'h264c 	:	o_val <= 16'b0110011101011101;
            14'h264d 	:	o_val <= 16'b0110011101011111;
            14'h264e 	:	o_val <= 16'b0110011101100001;
            14'h264f 	:	o_val <= 16'b0110011101100011;
            14'h2650 	:	o_val <= 16'b0110011101100101;
            14'h2651 	:	o_val <= 16'b0110011101100111;
            14'h2652 	:	o_val <= 16'b0110011101101001;
            14'h2653 	:	o_val <= 16'b0110011101101010;
            14'h2654 	:	o_val <= 16'b0110011101101100;
            14'h2655 	:	o_val <= 16'b0110011101101110;
            14'h2656 	:	o_val <= 16'b0110011101110000;
            14'h2657 	:	o_val <= 16'b0110011101110010;
            14'h2658 	:	o_val <= 16'b0110011101110100;
            14'h2659 	:	o_val <= 16'b0110011101110110;
            14'h265a 	:	o_val <= 16'b0110011101110111;
            14'h265b 	:	o_val <= 16'b0110011101111001;
            14'h265c 	:	o_val <= 16'b0110011101111011;
            14'h265d 	:	o_val <= 16'b0110011101111101;
            14'h265e 	:	o_val <= 16'b0110011101111111;
            14'h265f 	:	o_val <= 16'b0110011110000001;
            14'h2660 	:	o_val <= 16'b0110011110000010;
            14'h2661 	:	o_val <= 16'b0110011110000100;
            14'h2662 	:	o_val <= 16'b0110011110000110;
            14'h2663 	:	o_val <= 16'b0110011110001000;
            14'h2664 	:	o_val <= 16'b0110011110001010;
            14'h2665 	:	o_val <= 16'b0110011110001100;
            14'h2666 	:	o_val <= 16'b0110011110001110;
            14'h2667 	:	o_val <= 16'b0110011110001111;
            14'h2668 	:	o_val <= 16'b0110011110010001;
            14'h2669 	:	o_val <= 16'b0110011110010011;
            14'h266a 	:	o_val <= 16'b0110011110010101;
            14'h266b 	:	o_val <= 16'b0110011110010111;
            14'h266c 	:	o_val <= 16'b0110011110011001;
            14'h266d 	:	o_val <= 16'b0110011110011010;
            14'h266e 	:	o_val <= 16'b0110011110011100;
            14'h266f 	:	o_val <= 16'b0110011110011110;
            14'h2670 	:	o_val <= 16'b0110011110100000;
            14'h2671 	:	o_val <= 16'b0110011110100010;
            14'h2672 	:	o_val <= 16'b0110011110100100;
            14'h2673 	:	o_val <= 16'b0110011110100110;
            14'h2674 	:	o_val <= 16'b0110011110100111;
            14'h2675 	:	o_val <= 16'b0110011110101001;
            14'h2676 	:	o_val <= 16'b0110011110101011;
            14'h2677 	:	o_val <= 16'b0110011110101101;
            14'h2678 	:	o_val <= 16'b0110011110101111;
            14'h2679 	:	o_val <= 16'b0110011110110001;
            14'h267a 	:	o_val <= 16'b0110011110110010;
            14'h267b 	:	o_val <= 16'b0110011110110100;
            14'h267c 	:	o_val <= 16'b0110011110110110;
            14'h267d 	:	o_val <= 16'b0110011110111000;
            14'h267e 	:	o_val <= 16'b0110011110111010;
            14'h267f 	:	o_val <= 16'b0110011110111100;
            14'h2680 	:	o_val <= 16'b0110011110111101;
            14'h2681 	:	o_val <= 16'b0110011110111111;
            14'h2682 	:	o_val <= 16'b0110011111000001;
            14'h2683 	:	o_val <= 16'b0110011111000011;
            14'h2684 	:	o_val <= 16'b0110011111000101;
            14'h2685 	:	o_val <= 16'b0110011111000111;
            14'h2686 	:	o_val <= 16'b0110011111001001;
            14'h2687 	:	o_val <= 16'b0110011111001010;
            14'h2688 	:	o_val <= 16'b0110011111001100;
            14'h2689 	:	o_val <= 16'b0110011111001110;
            14'h268a 	:	o_val <= 16'b0110011111010000;
            14'h268b 	:	o_val <= 16'b0110011111010010;
            14'h268c 	:	o_val <= 16'b0110011111010100;
            14'h268d 	:	o_val <= 16'b0110011111010101;
            14'h268e 	:	o_val <= 16'b0110011111010111;
            14'h268f 	:	o_val <= 16'b0110011111011001;
            14'h2690 	:	o_val <= 16'b0110011111011011;
            14'h2691 	:	o_val <= 16'b0110011111011101;
            14'h2692 	:	o_val <= 16'b0110011111011111;
            14'h2693 	:	o_val <= 16'b0110011111100000;
            14'h2694 	:	o_val <= 16'b0110011111100010;
            14'h2695 	:	o_val <= 16'b0110011111100100;
            14'h2696 	:	o_val <= 16'b0110011111100110;
            14'h2697 	:	o_val <= 16'b0110011111101000;
            14'h2698 	:	o_val <= 16'b0110011111101010;
            14'h2699 	:	o_val <= 16'b0110011111101011;
            14'h269a 	:	o_val <= 16'b0110011111101101;
            14'h269b 	:	o_val <= 16'b0110011111101111;
            14'h269c 	:	o_val <= 16'b0110011111110001;
            14'h269d 	:	o_val <= 16'b0110011111110011;
            14'h269e 	:	o_val <= 16'b0110011111110101;
            14'h269f 	:	o_val <= 16'b0110011111110110;
            14'h26a0 	:	o_val <= 16'b0110011111111000;
            14'h26a1 	:	o_val <= 16'b0110011111111010;
            14'h26a2 	:	o_val <= 16'b0110011111111100;
            14'h26a3 	:	o_val <= 16'b0110011111111110;
            14'h26a4 	:	o_val <= 16'b0110100000000000;
            14'h26a5 	:	o_val <= 16'b0110100000000001;
            14'h26a6 	:	o_val <= 16'b0110100000000011;
            14'h26a7 	:	o_val <= 16'b0110100000000101;
            14'h26a8 	:	o_val <= 16'b0110100000000111;
            14'h26a9 	:	o_val <= 16'b0110100000001001;
            14'h26aa 	:	o_val <= 16'b0110100000001011;
            14'h26ab 	:	o_val <= 16'b0110100000001100;
            14'h26ac 	:	o_val <= 16'b0110100000001110;
            14'h26ad 	:	o_val <= 16'b0110100000010000;
            14'h26ae 	:	o_val <= 16'b0110100000010010;
            14'h26af 	:	o_val <= 16'b0110100000010100;
            14'h26b0 	:	o_val <= 16'b0110100000010110;
            14'h26b1 	:	o_val <= 16'b0110100000010111;
            14'h26b2 	:	o_val <= 16'b0110100000011001;
            14'h26b3 	:	o_val <= 16'b0110100000011011;
            14'h26b4 	:	o_val <= 16'b0110100000011101;
            14'h26b5 	:	o_val <= 16'b0110100000011111;
            14'h26b6 	:	o_val <= 16'b0110100000100000;
            14'h26b7 	:	o_val <= 16'b0110100000100010;
            14'h26b8 	:	o_val <= 16'b0110100000100100;
            14'h26b9 	:	o_val <= 16'b0110100000100110;
            14'h26ba 	:	o_val <= 16'b0110100000101000;
            14'h26bb 	:	o_val <= 16'b0110100000101010;
            14'h26bc 	:	o_val <= 16'b0110100000101011;
            14'h26bd 	:	o_val <= 16'b0110100000101101;
            14'h26be 	:	o_val <= 16'b0110100000101111;
            14'h26bf 	:	o_val <= 16'b0110100000110001;
            14'h26c0 	:	o_val <= 16'b0110100000110011;
            14'h26c1 	:	o_val <= 16'b0110100000110101;
            14'h26c2 	:	o_val <= 16'b0110100000110110;
            14'h26c3 	:	o_val <= 16'b0110100000111000;
            14'h26c4 	:	o_val <= 16'b0110100000111010;
            14'h26c5 	:	o_val <= 16'b0110100000111100;
            14'h26c6 	:	o_val <= 16'b0110100000111110;
            14'h26c7 	:	o_val <= 16'b0110100001000000;
            14'h26c8 	:	o_val <= 16'b0110100001000001;
            14'h26c9 	:	o_val <= 16'b0110100001000011;
            14'h26ca 	:	o_val <= 16'b0110100001000101;
            14'h26cb 	:	o_val <= 16'b0110100001000111;
            14'h26cc 	:	o_val <= 16'b0110100001001001;
            14'h26cd 	:	o_val <= 16'b0110100001001010;
            14'h26ce 	:	o_val <= 16'b0110100001001100;
            14'h26cf 	:	o_val <= 16'b0110100001001110;
            14'h26d0 	:	o_val <= 16'b0110100001010000;
            14'h26d1 	:	o_val <= 16'b0110100001010010;
            14'h26d2 	:	o_val <= 16'b0110100001010100;
            14'h26d3 	:	o_val <= 16'b0110100001010101;
            14'h26d4 	:	o_val <= 16'b0110100001010111;
            14'h26d5 	:	o_val <= 16'b0110100001011001;
            14'h26d6 	:	o_val <= 16'b0110100001011011;
            14'h26d7 	:	o_val <= 16'b0110100001011101;
            14'h26d8 	:	o_val <= 16'b0110100001011110;
            14'h26d9 	:	o_val <= 16'b0110100001100000;
            14'h26da 	:	o_val <= 16'b0110100001100010;
            14'h26db 	:	o_val <= 16'b0110100001100100;
            14'h26dc 	:	o_val <= 16'b0110100001100110;
            14'h26dd 	:	o_val <= 16'b0110100001101000;
            14'h26de 	:	o_val <= 16'b0110100001101001;
            14'h26df 	:	o_val <= 16'b0110100001101011;
            14'h26e0 	:	o_val <= 16'b0110100001101101;
            14'h26e1 	:	o_val <= 16'b0110100001101111;
            14'h26e2 	:	o_val <= 16'b0110100001110001;
            14'h26e3 	:	o_val <= 16'b0110100001110010;
            14'h26e4 	:	o_val <= 16'b0110100001110100;
            14'h26e5 	:	o_val <= 16'b0110100001110110;
            14'h26e6 	:	o_val <= 16'b0110100001111000;
            14'h26e7 	:	o_val <= 16'b0110100001111010;
            14'h26e8 	:	o_val <= 16'b0110100001111100;
            14'h26e9 	:	o_val <= 16'b0110100001111101;
            14'h26ea 	:	o_val <= 16'b0110100001111111;
            14'h26eb 	:	o_val <= 16'b0110100010000001;
            14'h26ec 	:	o_val <= 16'b0110100010000011;
            14'h26ed 	:	o_val <= 16'b0110100010000101;
            14'h26ee 	:	o_val <= 16'b0110100010000110;
            14'h26ef 	:	o_val <= 16'b0110100010001000;
            14'h26f0 	:	o_val <= 16'b0110100010001010;
            14'h26f1 	:	o_val <= 16'b0110100010001100;
            14'h26f2 	:	o_val <= 16'b0110100010001110;
            14'h26f3 	:	o_val <= 16'b0110100010001111;
            14'h26f4 	:	o_val <= 16'b0110100010010001;
            14'h26f5 	:	o_val <= 16'b0110100010010011;
            14'h26f6 	:	o_val <= 16'b0110100010010101;
            14'h26f7 	:	o_val <= 16'b0110100010010111;
            14'h26f8 	:	o_val <= 16'b0110100010011001;
            14'h26f9 	:	o_val <= 16'b0110100010011010;
            14'h26fa 	:	o_val <= 16'b0110100010011100;
            14'h26fb 	:	o_val <= 16'b0110100010011110;
            14'h26fc 	:	o_val <= 16'b0110100010100000;
            14'h26fd 	:	o_val <= 16'b0110100010100010;
            14'h26fe 	:	o_val <= 16'b0110100010100011;
            14'h26ff 	:	o_val <= 16'b0110100010100101;
            14'h2700 	:	o_val <= 16'b0110100010100111;
            14'h2701 	:	o_val <= 16'b0110100010101001;
            14'h2702 	:	o_val <= 16'b0110100010101011;
            14'h2703 	:	o_val <= 16'b0110100010101100;
            14'h2704 	:	o_val <= 16'b0110100010101110;
            14'h2705 	:	o_val <= 16'b0110100010110000;
            14'h2706 	:	o_val <= 16'b0110100010110010;
            14'h2707 	:	o_val <= 16'b0110100010110100;
            14'h2708 	:	o_val <= 16'b0110100010110101;
            14'h2709 	:	o_val <= 16'b0110100010110111;
            14'h270a 	:	o_val <= 16'b0110100010111001;
            14'h270b 	:	o_val <= 16'b0110100010111011;
            14'h270c 	:	o_val <= 16'b0110100010111101;
            14'h270d 	:	o_val <= 16'b0110100010111111;
            14'h270e 	:	o_val <= 16'b0110100011000000;
            14'h270f 	:	o_val <= 16'b0110100011000010;
            14'h2710 	:	o_val <= 16'b0110100011000100;
            14'h2711 	:	o_val <= 16'b0110100011000110;
            14'h2712 	:	o_val <= 16'b0110100011001000;
            14'h2713 	:	o_val <= 16'b0110100011001001;
            14'h2714 	:	o_val <= 16'b0110100011001011;
            14'h2715 	:	o_val <= 16'b0110100011001101;
            14'h2716 	:	o_val <= 16'b0110100011001111;
            14'h2717 	:	o_val <= 16'b0110100011010001;
            14'h2718 	:	o_val <= 16'b0110100011010010;
            14'h2719 	:	o_val <= 16'b0110100011010100;
            14'h271a 	:	o_val <= 16'b0110100011010110;
            14'h271b 	:	o_val <= 16'b0110100011011000;
            14'h271c 	:	o_val <= 16'b0110100011011010;
            14'h271d 	:	o_val <= 16'b0110100011011011;
            14'h271e 	:	o_val <= 16'b0110100011011101;
            14'h271f 	:	o_val <= 16'b0110100011011111;
            14'h2720 	:	o_val <= 16'b0110100011100001;
            14'h2721 	:	o_val <= 16'b0110100011100011;
            14'h2722 	:	o_val <= 16'b0110100011100100;
            14'h2723 	:	o_val <= 16'b0110100011100110;
            14'h2724 	:	o_val <= 16'b0110100011101000;
            14'h2725 	:	o_val <= 16'b0110100011101010;
            14'h2726 	:	o_val <= 16'b0110100011101100;
            14'h2727 	:	o_val <= 16'b0110100011101101;
            14'h2728 	:	o_val <= 16'b0110100011101111;
            14'h2729 	:	o_val <= 16'b0110100011110001;
            14'h272a 	:	o_val <= 16'b0110100011110011;
            14'h272b 	:	o_val <= 16'b0110100011110101;
            14'h272c 	:	o_val <= 16'b0110100011110110;
            14'h272d 	:	o_val <= 16'b0110100011111000;
            14'h272e 	:	o_val <= 16'b0110100011111010;
            14'h272f 	:	o_val <= 16'b0110100011111100;
            14'h2730 	:	o_val <= 16'b0110100011111110;
            14'h2731 	:	o_val <= 16'b0110100011111111;
            14'h2732 	:	o_val <= 16'b0110100100000001;
            14'h2733 	:	o_val <= 16'b0110100100000011;
            14'h2734 	:	o_val <= 16'b0110100100000101;
            14'h2735 	:	o_val <= 16'b0110100100000111;
            14'h2736 	:	o_val <= 16'b0110100100001000;
            14'h2737 	:	o_val <= 16'b0110100100001010;
            14'h2738 	:	o_val <= 16'b0110100100001100;
            14'h2739 	:	o_val <= 16'b0110100100001110;
            14'h273a 	:	o_val <= 16'b0110100100010000;
            14'h273b 	:	o_val <= 16'b0110100100010001;
            14'h273c 	:	o_val <= 16'b0110100100010011;
            14'h273d 	:	o_val <= 16'b0110100100010101;
            14'h273e 	:	o_val <= 16'b0110100100010111;
            14'h273f 	:	o_val <= 16'b0110100100011000;
            14'h2740 	:	o_val <= 16'b0110100100011010;
            14'h2741 	:	o_val <= 16'b0110100100011100;
            14'h2742 	:	o_val <= 16'b0110100100011110;
            14'h2743 	:	o_val <= 16'b0110100100100000;
            14'h2744 	:	o_val <= 16'b0110100100100001;
            14'h2745 	:	o_val <= 16'b0110100100100011;
            14'h2746 	:	o_val <= 16'b0110100100100101;
            14'h2747 	:	o_val <= 16'b0110100100100111;
            14'h2748 	:	o_val <= 16'b0110100100101001;
            14'h2749 	:	o_val <= 16'b0110100100101010;
            14'h274a 	:	o_val <= 16'b0110100100101100;
            14'h274b 	:	o_val <= 16'b0110100100101110;
            14'h274c 	:	o_val <= 16'b0110100100110000;
            14'h274d 	:	o_val <= 16'b0110100100110010;
            14'h274e 	:	o_val <= 16'b0110100100110011;
            14'h274f 	:	o_val <= 16'b0110100100110101;
            14'h2750 	:	o_val <= 16'b0110100100110111;
            14'h2751 	:	o_val <= 16'b0110100100111001;
            14'h2752 	:	o_val <= 16'b0110100100111011;
            14'h2753 	:	o_val <= 16'b0110100100111100;
            14'h2754 	:	o_val <= 16'b0110100100111110;
            14'h2755 	:	o_val <= 16'b0110100101000000;
            14'h2756 	:	o_val <= 16'b0110100101000010;
            14'h2757 	:	o_val <= 16'b0110100101000011;
            14'h2758 	:	o_val <= 16'b0110100101000101;
            14'h2759 	:	o_val <= 16'b0110100101000111;
            14'h275a 	:	o_val <= 16'b0110100101001001;
            14'h275b 	:	o_val <= 16'b0110100101001011;
            14'h275c 	:	o_val <= 16'b0110100101001100;
            14'h275d 	:	o_val <= 16'b0110100101001110;
            14'h275e 	:	o_val <= 16'b0110100101010000;
            14'h275f 	:	o_val <= 16'b0110100101010010;
            14'h2760 	:	o_val <= 16'b0110100101010100;
            14'h2761 	:	o_val <= 16'b0110100101010101;
            14'h2762 	:	o_val <= 16'b0110100101010111;
            14'h2763 	:	o_val <= 16'b0110100101011001;
            14'h2764 	:	o_val <= 16'b0110100101011011;
            14'h2765 	:	o_val <= 16'b0110100101011100;
            14'h2766 	:	o_val <= 16'b0110100101011110;
            14'h2767 	:	o_val <= 16'b0110100101100000;
            14'h2768 	:	o_val <= 16'b0110100101100010;
            14'h2769 	:	o_val <= 16'b0110100101100100;
            14'h276a 	:	o_val <= 16'b0110100101100101;
            14'h276b 	:	o_val <= 16'b0110100101100111;
            14'h276c 	:	o_val <= 16'b0110100101101001;
            14'h276d 	:	o_val <= 16'b0110100101101011;
            14'h276e 	:	o_val <= 16'b0110100101101101;
            14'h276f 	:	o_val <= 16'b0110100101101110;
            14'h2770 	:	o_val <= 16'b0110100101110000;
            14'h2771 	:	o_val <= 16'b0110100101110010;
            14'h2772 	:	o_val <= 16'b0110100101110100;
            14'h2773 	:	o_val <= 16'b0110100101110101;
            14'h2774 	:	o_val <= 16'b0110100101110111;
            14'h2775 	:	o_val <= 16'b0110100101111001;
            14'h2776 	:	o_val <= 16'b0110100101111011;
            14'h2777 	:	o_val <= 16'b0110100101111101;
            14'h2778 	:	o_val <= 16'b0110100101111110;
            14'h2779 	:	o_val <= 16'b0110100110000000;
            14'h277a 	:	o_val <= 16'b0110100110000010;
            14'h277b 	:	o_val <= 16'b0110100110000100;
            14'h277c 	:	o_val <= 16'b0110100110000101;
            14'h277d 	:	o_val <= 16'b0110100110000111;
            14'h277e 	:	o_val <= 16'b0110100110001001;
            14'h277f 	:	o_val <= 16'b0110100110001011;
            14'h2780 	:	o_val <= 16'b0110100110001101;
            14'h2781 	:	o_val <= 16'b0110100110001110;
            14'h2782 	:	o_val <= 16'b0110100110010000;
            14'h2783 	:	o_val <= 16'b0110100110010010;
            14'h2784 	:	o_val <= 16'b0110100110010100;
            14'h2785 	:	o_val <= 16'b0110100110010101;
            14'h2786 	:	o_val <= 16'b0110100110010111;
            14'h2787 	:	o_val <= 16'b0110100110011001;
            14'h2788 	:	o_val <= 16'b0110100110011011;
            14'h2789 	:	o_val <= 16'b0110100110011101;
            14'h278a 	:	o_val <= 16'b0110100110011110;
            14'h278b 	:	o_val <= 16'b0110100110100000;
            14'h278c 	:	o_val <= 16'b0110100110100010;
            14'h278d 	:	o_val <= 16'b0110100110100100;
            14'h278e 	:	o_val <= 16'b0110100110100101;
            14'h278f 	:	o_val <= 16'b0110100110100111;
            14'h2790 	:	o_val <= 16'b0110100110101001;
            14'h2791 	:	o_val <= 16'b0110100110101011;
            14'h2792 	:	o_val <= 16'b0110100110101100;
            14'h2793 	:	o_val <= 16'b0110100110101110;
            14'h2794 	:	o_val <= 16'b0110100110110000;
            14'h2795 	:	o_val <= 16'b0110100110110010;
            14'h2796 	:	o_val <= 16'b0110100110110100;
            14'h2797 	:	o_val <= 16'b0110100110110101;
            14'h2798 	:	o_val <= 16'b0110100110110111;
            14'h2799 	:	o_val <= 16'b0110100110111001;
            14'h279a 	:	o_val <= 16'b0110100110111011;
            14'h279b 	:	o_val <= 16'b0110100110111100;
            14'h279c 	:	o_val <= 16'b0110100110111110;
            14'h279d 	:	o_val <= 16'b0110100111000000;
            14'h279e 	:	o_val <= 16'b0110100111000010;
            14'h279f 	:	o_val <= 16'b0110100111000100;
            14'h27a0 	:	o_val <= 16'b0110100111000101;
            14'h27a1 	:	o_val <= 16'b0110100111000111;
            14'h27a2 	:	o_val <= 16'b0110100111001001;
            14'h27a3 	:	o_val <= 16'b0110100111001011;
            14'h27a4 	:	o_val <= 16'b0110100111001100;
            14'h27a5 	:	o_val <= 16'b0110100111001110;
            14'h27a6 	:	o_val <= 16'b0110100111010000;
            14'h27a7 	:	o_val <= 16'b0110100111010010;
            14'h27a8 	:	o_val <= 16'b0110100111010011;
            14'h27a9 	:	o_val <= 16'b0110100111010101;
            14'h27aa 	:	o_val <= 16'b0110100111010111;
            14'h27ab 	:	o_val <= 16'b0110100111011001;
            14'h27ac 	:	o_val <= 16'b0110100111011010;
            14'h27ad 	:	o_val <= 16'b0110100111011100;
            14'h27ae 	:	o_val <= 16'b0110100111011110;
            14'h27af 	:	o_val <= 16'b0110100111100000;
            14'h27b0 	:	o_val <= 16'b0110100111100010;
            14'h27b1 	:	o_val <= 16'b0110100111100011;
            14'h27b2 	:	o_val <= 16'b0110100111100101;
            14'h27b3 	:	o_val <= 16'b0110100111100111;
            14'h27b4 	:	o_val <= 16'b0110100111101001;
            14'h27b5 	:	o_val <= 16'b0110100111101010;
            14'h27b6 	:	o_val <= 16'b0110100111101100;
            14'h27b7 	:	o_val <= 16'b0110100111101110;
            14'h27b8 	:	o_val <= 16'b0110100111110000;
            14'h27b9 	:	o_val <= 16'b0110100111110001;
            14'h27ba 	:	o_val <= 16'b0110100111110011;
            14'h27bb 	:	o_val <= 16'b0110100111110101;
            14'h27bc 	:	o_val <= 16'b0110100111110111;
            14'h27bd 	:	o_val <= 16'b0110100111111000;
            14'h27be 	:	o_val <= 16'b0110100111111010;
            14'h27bf 	:	o_val <= 16'b0110100111111100;
            14'h27c0 	:	o_val <= 16'b0110100111111110;
            14'h27c1 	:	o_val <= 16'b0110101000000000;
            14'h27c2 	:	o_val <= 16'b0110101000000001;
            14'h27c3 	:	o_val <= 16'b0110101000000011;
            14'h27c4 	:	o_val <= 16'b0110101000000101;
            14'h27c5 	:	o_val <= 16'b0110101000000111;
            14'h27c6 	:	o_val <= 16'b0110101000001000;
            14'h27c7 	:	o_val <= 16'b0110101000001010;
            14'h27c8 	:	o_val <= 16'b0110101000001100;
            14'h27c9 	:	o_val <= 16'b0110101000001110;
            14'h27ca 	:	o_val <= 16'b0110101000001111;
            14'h27cb 	:	o_val <= 16'b0110101000010001;
            14'h27cc 	:	o_val <= 16'b0110101000010011;
            14'h27cd 	:	o_val <= 16'b0110101000010101;
            14'h27ce 	:	o_val <= 16'b0110101000010110;
            14'h27cf 	:	o_val <= 16'b0110101000011000;
            14'h27d0 	:	o_val <= 16'b0110101000011010;
            14'h27d1 	:	o_val <= 16'b0110101000011100;
            14'h27d2 	:	o_val <= 16'b0110101000011101;
            14'h27d3 	:	o_val <= 16'b0110101000011111;
            14'h27d4 	:	o_val <= 16'b0110101000100001;
            14'h27d5 	:	o_val <= 16'b0110101000100011;
            14'h27d6 	:	o_val <= 16'b0110101000100100;
            14'h27d7 	:	o_val <= 16'b0110101000100110;
            14'h27d8 	:	o_val <= 16'b0110101000101000;
            14'h27d9 	:	o_val <= 16'b0110101000101010;
            14'h27da 	:	o_val <= 16'b0110101000101011;
            14'h27db 	:	o_val <= 16'b0110101000101101;
            14'h27dc 	:	o_val <= 16'b0110101000101111;
            14'h27dd 	:	o_val <= 16'b0110101000110001;
            14'h27de 	:	o_val <= 16'b0110101000110010;
            14'h27df 	:	o_val <= 16'b0110101000110100;
            14'h27e0 	:	o_val <= 16'b0110101000110110;
            14'h27e1 	:	o_val <= 16'b0110101000111000;
            14'h27e2 	:	o_val <= 16'b0110101000111001;
            14'h27e3 	:	o_val <= 16'b0110101000111011;
            14'h27e4 	:	o_val <= 16'b0110101000111101;
            14'h27e5 	:	o_val <= 16'b0110101000111111;
            14'h27e6 	:	o_val <= 16'b0110101001000001;
            14'h27e7 	:	o_val <= 16'b0110101001000010;
            14'h27e8 	:	o_val <= 16'b0110101001000100;
            14'h27e9 	:	o_val <= 16'b0110101001000110;
            14'h27ea 	:	o_val <= 16'b0110101001001000;
            14'h27eb 	:	o_val <= 16'b0110101001001001;
            14'h27ec 	:	o_val <= 16'b0110101001001011;
            14'h27ed 	:	o_val <= 16'b0110101001001101;
            14'h27ee 	:	o_val <= 16'b0110101001001111;
            14'h27ef 	:	o_val <= 16'b0110101001010000;
            14'h27f0 	:	o_val <= 16'b0110101001010010;
            14'h27f1 	:	o_val <= 16'b0110101001010100;
            14'h27f2 	:	o_val <= 16'b0110101001010110;
            14'h27f3 	:	o_val <= 16'b0110101001010111;
            14'h27f4 	:	o_val <= 16'b0110101001011001;
            14'h27f5 	:	o_val <= 16'b0110101001011011;
            14'h27f6 	:	o_val <= 16'b0110101001011101;
            14'h27f7 	:	o_val <= 16'b0110101001011110;
            14'h27f8 	:	o_val <= 16'b0110101001100000;
            14'h27f9 	:	o_val <= 16'b0110101001100010;
            14'h27fa 	:	o_val <= 16'b0110101001100011;
            14'h27fb 	:	o_val <= 16'b0110101001100101;
            14'h27fc 	:	o_val <= 16'b0110101001100111;
            14'h27fd 	:	o_val <= 16'b0110101001101001;
            14'h27fe 	:	o_val <= 16'b0110101001101010;
            14'h27ff 	:	o_val <= 16'b0110101001101100;
            14'h2800 	:	o_val <= 16'b0110101001101110;
            14'h2801 	:	o_val <= 16'b0110101001110000;
            14'h2802 	:	o_val <= 16'b0110101001110001;
            14'h2803 	:	o_val <= 16'b0110101001110011;
            14'h2804 	:	o_val <= 16'b0110101001110101;
            14'h2805 	:	o_val <= 16'b0110101001110111;
            14'h2806 	:	o_val <= 16'b0110101001111000;
            14'h2807 	:	o_val <= 16'b0110101001111010;
            14'h2808 	:	o_val <= 16'b0110101001111100;
            14'h2809 	:	o_val <= 16'b0110101001111110;
            14'h280a 	:	o_val <= 16'b0110101001111111;
            14'h280b 	:	o_val <= 16'b0110101010000001;
            14'h280c 	:	o_val <= 16'b0110101010000011;
            14'h280d 	:	o_val <= 16'b0110101010000101;
            14'h280e 	:	o_val <= 16'b0110101010000110;
            14'h280f 	:	o_val <= 16'b0110101010001000;
            14'h2810 	:	o_val <= 16'b0110101010001010;
            14'h2811 	:	o_val <= 16'b0110101010001100;
            14'h2812 	:	o_val <= 16'b0110101010001101;
            14'h2813 	:	o_val <= 16'b0110101010001111;
            14'h2814 	:	o_val <= 16'b0110101010010001;
            14'h2815 	:	o_val <= 16'b0110101010010011;
            14'h2816 	:	o_val <= 16'b0110101010010100;
            14'h2817 	:	o_val <= 16'b0110101010010110;
            14'h2818 	:	o_val <= 16'b0110101010011000;
            14'h2819 	:	o_val <= 16'b0110101010011010;
            14'h281a 	:	o_val <= 16'b0110101010011011;
            14'h281b 	:	o_val <= 16'b0110101010011101;
            14'h281c 	:	o_val <= 16'b0110101010011111;
            14'h281d 	:	o_val <= 16'b0110101010100000;
            14'h281e 	:	o_val <= 16'b0110101010100010;
            14'h281f 	:	o_val <= 16'b0110101010100100;
            14'h2820 	:	o_val <= 16'b0110101010100110;
            14'h2821 	:	o_val <= 16'b0110101010100111;
            14'h2822 	:	o_val <= 16'b0110101010101001;
            14'h2823 	:	o_val <= 16'b0110101010101011;
            14'h2824 	:	o_val <= 16'b0110101010101101;
            14'h2825 	:	o_val <= 16'b0110101010101110;
            14'h2826 	:	o_val <= 16'b0110101010110000;
            14'h2827 	:	o_val <= 16'b0110101010110010;
            14'h2828 	:	o_val <= 16'b0110101010110100;
            14'h2829 	:	o_val <= 16'b0110101010110101;
            14'h282a 	:	o_val <= 16'b0110101010110111;
            14'h282b 	:	o_val <= 16'b0110101010111001;
            14'h282c 	:	o_val <= 16'b0110101010111011;
            14'h282d 	:	o_val <= 16'b0110101010111100;
            14'h282e 	:	o_val <= 16'b0110101010111110;
            14'h282f 	:	o_val <= 16'b0110101011000000;
            14'h2830 	:	o_val <= 16'b0110101011000001;
            14'h2831 	:	o_val <= 16'b0110101011000011;
            14'h2832 	:	o_val <= 16'b0110101011000101;
            14'h2833 	:	o_val <= 16'b0110101011000111;
            14'h2834 	:	o_val <= 16'b0110101011001000;
            14'h2835 	:	o_val <= 16'b0110101011001010;
            14'h2836 	:	o_val <= 16'b0110101011001100;
            14'h2837 	:	o_val <= 16'b0110101011001110;
            14'h2838 	:	o_val <= 16'b0110101011001111;
            14'h2839 	:	o_val <= 16'b0110101011010001;
            14'h283a 	:	o_val <= 16'b0110101011010011;
            14'h283b 	:	o_val <= 16'b0110101011010101;
            14'h283c 	:	o_val <= 16'b0110101011010110;
            14'h283d 	:	o_val <= 16'b0110101011011000;
            14'h283e 	:	o_val <= 16'b0110101011011010;
            14'h283f 	:	o_val <= 16'b0110101011011011;
            14'h2840 	:	o_val <= 16'b0110101011011101;
            14'h2841 	:	o_val <= 16'b0110101011011111;
            14'h2842 	:	o_val <= 16'b0110101011100001;
            14'h2843 	:	o_val <= 16'b0110101011100010;
            14'h2844 	:	o_val <= 16'b0110101011100100;
            14'h2845 	:	o_val <= 16'b0110101011100110;
            14'h2846 	:	o_val <= 16'b0110101011101000;
            14'h2847 	:	o_val <= 16'b0110101011101001;
            14'h2848 	:	o_val <= 16'b0110101011101011;
            14'h2849 	:	o_val <= 16'b0110101011101101;
            14'h284a 	:	o_val <= 16'b0110101011101110;
            14'h284b 	:	o_val <= 16'b0110101011110000;
            14'h284c 	:	o_val <= 16'b0110101011110010;
            14'h284d 	:	o_val <= 16'b0110101011110100;
            14'h284e 	:	o_val <= 16'b0110101011110101;
            14'h284f 	:	o_val <= 16'b0110101011110111;
            14'h2850 	:	o_val <= 16'b0110101011111001;
            14'h2851 	:	o_val <= 16'b0110101011111011;
            14'h2852 	:	o_val <= 16'b0110101011111100;
            14'h2853 	:	o_val <= 16'b0110101011111110;
            14'h2854 	:	o_val <= 16'b0110101100000000;
            14'h2855 	:	o_val <= 16'b0110101100000001;
            14'h2856 	:	o_val <= 16'b0110101100000011;
            14'h2857 	:	o_val <= 16'b0110101100000101;
            14'h2858 	:	o_val <= 16'b0110101100000111;
            14'h2859 	:	o_val <= 16'b0110101100001000;
            14'h285a 	:	o_val <= 16'b0110101100001010;
            14'h285b 	:	o_val <= 16'b0110101100001100;
            14'h285c 	:	o_val <= 16'b0110101100001101;
            14'h285d 	:	o_val <= 16'b0110101100001111;
            14'h285e 	:	o_val <= 16'b0110101100010001;
            14'h285f 	:	o_val <= 16'b0110101100010011;
            14'h2860 	:	o_val <= 16'b0110101100010100;
            14'h2861 	:	o_val <= 16'b0110101100010110;
            14'h2862 	:	o_val <= 16'b0110101100011000;
            14'h2863 	:	o_val <= 16'b0110101100011010;
            14'h2864 	:	o_val <= 16'b0110101100011011;
            14'h2865 	:	o_val <= 16'b0110101100011101;
            14'h2866 	:	o_val <= 16'b0110101100011111;
            14'h2867 	:	o_val <= 16'b0110101100100000;
            14'h2868 	:	o_val <= 16'b0110101100100010;
            14'h2869 	:	o_val <= 16'b0110101100100100;
            14'h286a 	:	o_val <= 16'b0110101100100110;
            14'h286b 	:	o_val <= 16'b0110101100100111;
            14'h286c 	:	o_val <= 16'b0110101100101001;
            14'h286d 	:	o_val <= 16'b0110101100101011;
            14'h286e 	:	o_val <= 16'b0110101100101100;
            14'h286f 	:	o_val <= 16'b0110101100101110;
            14'h2870 	:	o_val <= 16'b0110101100110000;
            14'h2871 	:	o_val <= 16'b0110101100110010;
            14'h2872 	:	o_val <= 16'b0110101100110011;
            14'h2873 	:	o_val <= 16'b0110101100110101;
            14'h2874 	:	o_val <= 16'b0110101100110111;
            14'h2875 	:	o_val <= 16'b0110101100111000;
            14'h2876 	:	o_val <= 16'b0110101100111010;
            14'h2877 	:	o_val <= 16'b0110101100111100;
            14'h2878 	:	o_val <= 16'b0110101100111110;
            14'h2879 	:	o_val <= 16'b0110101100111111;
            14'h287a 	:	o_val <= 16'b0110101101000001;
            14'h287b 	:	o_val <= 16'b0110101101000011;
            14'h287c 	:	o_val <= 16'b0110101101000100;
            14'h287d 	:	o_val <= 16'b0110101101000110;
            14'h287e 	:	o_val <= 16'b0110101101001000;
            14'h287f 	:	o_val <= 16'b0110101101001010;
            14'h2880 	:	o_val <= 16'b0110101101001011;
            14'h2881 	:	o_val <= 16'b0110101101001101;
            14'h2882 	:	o_val <= 16'b0110101101001111;
            14'h2883 	:	o_val <= 16'b0110101101010000;
            14'h2884 	:	o_val <= 16'b0110101101010010;
            14'h2885 	:	o_val <= 16'b0110101101010100;
            14'h2886 	:	o_val <= 16'b0110101101010110;
            14'h2887 	:	o_val <= 16'b0110101101010111;
            14'h2888 	:	o_val <= 16'b0110101101011001;
            14'h2889 	:	o_val <= 16'b0110101101011011;
            14'h288a 	:	o_val <= 16'b0110101101011100;
            14'h288b 	:	o_val <= 16'b0110101101011110;
            14'h288c 	:	o_val <= 16'b0110101101100000;
            14'h288d 	:	o_val <= 16'b0110101101100010;
            14'h288e 	:	o_val <= 16'b0110101101100011;
            14'h288f 	:	o_val <= 16'b0110101101100101;
            14'h2890 	:	o_val <= 16'b0110101101100111;
            14'h2891 	:	o_val <= 16'b0110101101101000;
            14'h2892 	:	o_val <= 16'b0110101101101010;
            14'h2893 	:	o_val <= 16'b0110101101101100;
            14'h2894 	:	o_val <= 16'b0110101101101110;
            14'h2895 	:	o_val <= 16'b0110101101101111;
            14'h2896 	:	o_val <= 16'b0110101101110001;
            14'h2897 	:	o_val <= 16'b0110101101110011;
            14'h2898 	:	o_val <= 16'b0110101101110100;
            14'h2899 	:	o_val <= 16'b0110101101110110;
            14'h289a 	:	o_val <= 16'b0110101101111000;
            14'h289b 	:	o_val <= 16'b0110101101111001;
            14'h289c 	:	o_val <= 16'b0110101101111011;
            14'h289d 	:	o_val <= 16'b0110101101111101;
            14'h289e 	:	o_val <= 16'b0110101101111111;
            14'h289f 	:	o_val <= 16'b0110101110000000;
            14'h28a0 	:	o_val <= 16'b0110101110000010;
            14'h28a1 	:	o_val <= 16'b0110101110000100;
            14'h28a2 	:	o_val <= 16'b0110101110000101;
            14'h28a3 	:	o_val <= 16'b0110101110000111;
            14'h28a4 	:	o_val <= 16'b0110101110001001;
            14'h28a5 	:	o_val <= 16'b0110101110001011;
            14'h28a6 	:	o_val <= 16'b0110101110001100;
            14'h28a7 	:	o_val <= 16'b0110101110001110;
            14'h28a8 	:	o_val <= 16'b0110101110010000;
            14'h28a9 	:	o_val <= 16'b0110101110010001;
            14'h28aa 	:	o_val <= 16'b0110101110010011;
            14'h28ab 	:	o_val <= 16'b0110101110010101;
            14'h28ac 	:	o_val <= 16'b0110101110010110;
            14'h28ad 	:	o_val <= 16'b0110101110011000;
            14'h28ae 	:	o_val <= 16'b0110101110011010;
            14'h28af 	:	o_val <= 16'b0110101110011100;
            14'h28b0 	:	o_val <= 16'b0110101110011101;
            14'h28b1 	:	o_val <= 16'b0110101110011111;
            14'h28b2 	:	o_val <= 16'b0110101110100001;
            14'h28b3 	:	o_val <= 16'b0110101110100010;
            14'h28b4 	:	o_val <= 16'b0110101110100100;
            14'h28b5 	:	o_val <= 16'b0110101110100110;
            14'h28b6 	:	o_val <= 16'b0110101110100111;
            14'h28b7 	:	o_val <= 16'b0110101110101001;
            14'h28b8 	:	o_val <= 16'b0110101110101011;
            14'h28b9 	:	o_val <= 16'b0110101110101101;
            14'h28ba 	:	o_val <= 16'b0110101110101110;
            14'h28bb 	:	o_val <= 16'b0110101110110000;
            14'h28bc 	:	o_val <= 16'b0110101110110010;
            14'h28bd 	:	o_val <= 16'b0110101110110011;
            14'h28be 	:	o_val <= 16'b0110101110110101;
            14'h28bf 	:	o_val <= 16'b0110101110110111;
            14'h28c0 	:	o_val <= 16'b0110101110111000;
            14'h28c1 	:	o_val <= 16'b0110101110111010;
            14'h28c2 	:	o_val <= 16'b0110101110111100;
            14'h28c3 	:	o_val <= 16'b0110101110111110;
            14'h28c4 	:	o_val <= 16'b0110101110111111;
            14'h28c5 	:	o_val <= 16'b0110101111000001;
            14'h28c6 	:	o_val <= 16'b0110101111000011;
            14'h28c7 	:	o_val <= 16'b0110101111000100;
            14'h28c8 	:	o_val <= 16'b0110101111000110;
            14'h28c9 	:	o_val <= 16'b0110101111001000;
            14'h28ca 	:	o_val <= 16'b0110101111001001;
            14'h28cb 	:	o_val <= 16'b0110101111001011;
            14'h28cc 	:	o_val <= 16'b0110101111001101;
            14'h28cd 	:	o_val <= 16'b0110101111001110;
            14'h28ce 	:	o_val <= 16'b0110101111010000;
            14'h28cf 	:	o_val <= 16'b0110101111010010;
            14'h28d0 	:	o_val <= 16'b0110101111010100;
            14'h28d1 	:	o_val <= 16'b0110101111010101;
            14'h28d2 	:	o_val <= 16'b0110101111010111;
            14'h28d3 	:	o_val <= 16'b0110101111011001;
            14'h28d4 	:	o_val <= 16'b0110101111011010;
            14'h28d5 	:	o_val <= 16'b0110101111011100;
            14'h28d6 	:	o_val <= 16'b0110101111011110;
            14'h28d7 	:	o_val <= 16'b0110101111011111;
            14'h28d8 	:	o_val <= 16'b0110101111100001;
            14'h28d9 	:	o_val <= 16'b0110101111100011;
            14'h28da 	:	o_val <= 16'b0110101111100100;
            14'h28db 	:	o_val <= 16'b0110101111100110;
            14'h28dc 	:	o_val <= 16'b0110101111101000;
            14'h28dd 	:	o_val <= 16'b0110101111101010;
            14'h28de 	:	o_val <= 16'b0110101111101011;
            14'h28df 	:	o_val <= 16'b0110101111101101;
            14'h28e0 	:	o_val <= 16'b0110101111101111;
            14'h28e1 	:	o_val <= 16'b0110101111110000;
            14'h28e2 	:	o_val <= 16'b0110101111110010;
            14'h28e3 	:	o_val <= 16'b0110101111110100;
            14'h28e4 	:	o_val <= 16'b0110101111110101;
            14'h28e5 	:	o_val <= 16'b0110101111110111;
            14'h28e6 	:	o_val <= 16'b0110101111111001;
            14'h28e7 	:	o_val <= 16'b0110101111111010;
            14'h28e8 	:	o_val <= 16'b0110101111111100;
            14'h28e9 	:	o_val <= 16'b0110101111111110;
            14'h28ea 	:	o_val <= 16'b0110101111111111;
            14'h28eb 	:	o_val <= 16'b0110110000000001;
            14'h28ec 	:	o_val <= 16'b0110110000000011;
            14'h28ed 	:	o_val <= 16'b0110110000000101;
            14'h28ee 	:	o_val <= 16'b0110110000000110;
            14'h28ef 	:	o_val <= 16'b0110110000001000;
            14'h28f0 	:	o_val <= 16'b0110110000001010;
            14'h28f1 	:	o_val <= 16'b0110110000001011;
            14'h28f2 	:	o_val <= 16'b0110110000001101;
            14'h28f3 	:	o_val <= 16'b0110110000001111;
            14'h28f4 	:	o_val <= 16'b0110110000010000;
            14'h28f5 	:	o_val <= 16'b0110110000010010;
            14'h28f6 	:	o_val <= 16'b0110110000010100;
            14'h28f7 	:	o_val <= 16'b0110110000010101;
            14'h28f8 	:	o_val <= 16'b0110110000010111;
            14'h28f9 	:	o_val <= 16'b0110110000011001;
            14'h28fa 	:	o_val <= 16'b0110110000011010;
            14'h28fb 	:	o_val <= 16'b0110110000011100;
            14'h28fc 	:	o_val <= 16'b0110110000011110;
            14'h28fd 	:	o_val <= 16'b0110110000011111;
            14'h28fe 	:	o_val <= 16'b0110110000100001;
            14'h28ff 	:	o_val <= 16'b0110110000100011;
            14'h2900 	:	o_val <= 16'b0110110000100101;
            14'h2901 	:	o_val <= 16'b0110110000100110;
            14'h2902 	:	o_val <= 16'b0110110000101000;
            14'h2903 	:	o_val <= 16'b0110110000101010;
            14'h2904 	:	o_val <= 16'b0110110000101011;
            14'h2905 	:	o_val <= 16'b0110110000101101;
            14'h2906 	:	o_val <= 16'b0110110000101111;
            14'h2907 	:	o_val <= 16'b0110110000110000;
            14'h2908 	:	o_val <= 16'b0110110000110010;
            14'h2909 	:	o_val <= 16'b0110110000110100;
            14'h290a 	:	o_val <= 16'b0110110000110101;
            14'h290b 	:	o_val <= 16'b0110110000110111;
            14'h290c 	:	o_val <= 16'b0110110000111001;
            14'h290d 	:	o_val <= 16'b0110110000111010;
            14'h290e 	:	o_val <= 16'b0110110000111100;
            14'h290f 	:	o_val <= 16'b0110110000111110;
            14'h2910 	:	o_val <= 16'b0110110000111111;
            14'h2911 	:	o_val <= 16'b0110110001000001;
            14'h2912 	:	o_val <= 16'b0110110001000011;
            14'h2913 	:	o_val <= 16'b0110110001000100;
            14'h2914 	:	o_val <= 16'b0110110001000110;
            14'h2915 	:	o_val <= 16'b0110110001001000;
            14'h2916 	:	o_val <= 16'b0110110001001001;
            14'h2917 	:	o_val <= 16'b0110110001001011;
            14'h2918 	:	o_val <= 16'b0110110001001101;
            14'h2919 	:	o_val <= 16'b0110110001001110;
            14'h291a 	:	o_val <= 16'b0110110001010000;
            14'h291b 	:	o_val <= 16'b0110110001010010;
            14'h291c 	:	o_val <= 16'b0110110001010011;
            14'h291d 	:	o_val <= 16'b0110110001010101;
            14'h291e 	:	o_val <= 16'b0110110001010111;
            14'h291f 	:	o_val <= 16'b0110110001011000;
            14'h2920 	:	o_val <= 16'b0110110001011010;
            14'h2921 	:	o_val <= 16'b0110110001011100;
            14'h2922 	:	o_val <= 16'b0110110001011101;
            14'h2923 	:	o_val <= 16'b0110110001011111;
            14'h2924 	:	o_val <= 16'b0110110001100001;
            14'h2925 	:	o_val <= 16'b0110110001100011;
            14'h2926 	:	o_val <= 16'b0110110001100100;
            14'h2927 	:	o_val <= 16'b0110110001100110;
            14'h2928 	:	o_val <= 16'b0110110001101000;
            14'h2929 	:	o_val <= 16'b0110110001101001;
            14'h292a 	:	o_val <= 16'b0110110001101011;
            14'h292b 	:	o_val <= 16'b0110110001101101;
            14'h292c 	:	o_val <= 16'b0110110001101110;
            14'h292d 	:	o_val <= 16'b0110110001110000;
            14'h292e 	:	o_val <= 16'b0110110001110010;
            14'h292f 	:	o_val <= 16'b0110110001110011;
            14'h2930 	:	o_val <= 16'b0110110001110101;
            14'h2931 	:	o_val <= 16'b0110110001110111;
            14'h2932 	:	o_val <= 16'b0110110001111000;
            14'h2933 	:	o_val <= 16'b0110110001111010;
            14'h2934 	:	o_val <= 16'b0110110001111100;
            14'h2935 	:	o_val <= 16'b0110110001111101;
            14'h2936 	:	o_val <= 16'b0110110001111111;
            14'h2937 	:	o_val <= 16'b0110110010000001;
            14'h2938 	:	o_val <= 16'b0110110010000010;
            14'h2939 	:	o_val <= 16'b0110110010000100;
            14'h293a 	:	o_val <= 16'b0110110010000110;
            14'h293b 	:	o_val <= 16'b0110110010000111;
            14'h293c 	:	o_val <= 16'b0110110010001001;
            14'h293d 	:	o_val <= 16'b0110110010001011;
            14'h293e 	:	o_val <= 16'b0110110010001100;
            14'h293f 	:	o_val <= 16'b0110110010001110;
            14'h2940 	:	o_val <= 16'b0110110010010000;
            14'h2941 	:	o_val <= 16'b0110110010010001;
            14'h2942 	:	o_val <= 16'b0110110010010011;
            14'h2943 	:	o_val <= 16'b0110110010010101;
            14'h2944 	:	o_val <= 16'b0110110010010110;
            14'h2945 	:	o_val <= 16'b0110110010011000;
            14'h2946 	:	o_val <= 16'b0110110010011010;
            14'h2947 	:	o_val <= 16'b0110110010011011;
            14'h2948 	:	o_val <= 16'b0110110010011101;
            14'h2949 	:	o_val <= 16'b0110110010011111;
            14'h294a 	:	o_val <= 16'b0110110010100000;
            14'h294b 	:	o_val <= 16'b0110110010100010;
            14'h294c 	:	o_val <= 16'b0110110010100011;
            14'h294d 	:	o_val <= 16'b0110110010100101;
            14'h294e 	:	o_val <= 16'b0110110010100111;
            14'h294f 	:	o_val <= 16'b0110110010101000;
            14'h2950 	:	o_val <= 16'b0110110010101010;
            14'h2951 	:	o_val <= 16'b0110110010101100;
            14'h2952 	:	o_val <= 16'b0110110010101101;
            14'h2953 	:	o_val <= 16'b0110110010101111;
            14'h2954 	:	o_val <= 16'b0110110010110001;
            14'h2955 	:	o_val <= 16'b0110110010110010;
            14'h2956 	:	o_val <= 16'b0110110010110100;
            14'h2957 	:	o_val <= 16'b0110110010110110;
            14'h2958 	:	o_val <= 16'b0110110010110111;
            14'h2959 	:	o_val <= 16'b0110110010111001;
            14'h295a 	:	o_val <= 16'b0110110010111011;
            14'h295b 	:	o_val <= 16'b0110110010111100;
            14'h295c 	:	o_val <= 16'b0110110010111110;
            14'h295d 	:	o_val <= 16'b0110110011000000;
            14'h295e 	:	o_val <= 16'b0110110011000001;
            14'h295f 	:	o_val <= 16'b0110110011000011;
            14'h2960 	:	o_val <= 16'b0110110011000101;
            14'h2961 	:	o_val <= 16'b0110110011000110;
            14'h2962 	:	o_val <= 16'b0110110011001000;
            14'h2963 	:	o_val <= 16'b0110110011001010;
            14'h2964 	:	o_val <= 16'b0110110011001011;
            14'h2965 	:	o_val <= 16'b0110110011001101;
            14'h2966 	:	o_val <= 16'b0110110011001111;
            14'h2967 	:	o_val <= 16'b0110110011010000;
            14'h2968 	:	o_val <= 16'b0110110011010010;
            14'h2969 	:	o_val <= 16'b0110110011010100;
            14'h296a 	:	o_val <= 16'b0110110011010101;
            14'h296b 	:	o_val <= 16'b0110110011010111;
            14'h296c 	:	o_val <= 16'b0110110011011001;
            14'h296d 	:	o_val <= 16'b0110110011011010;
            14'h296e 	:	o_val <= 16'b0110110011011100;
            14'h296f 	:	o_val <= 16'b0110110011011101;
            14'h2970 	:	o_val <= 16'b0110110011011111;
            14'h2971 	:	o_val <= 16'b0110110011100001;
            14'h2972 	:	o_val <= 16'b0110110011100010;
            14'h2973 	:	o_val <= 16'b0110110011100100;
            14'h2974 	:	o_val <= 16'b0110110011100110;
            14'h2975 	:	o_val <= 16'b0110110011100111;
            14'h2976 	:	o_val <= 16'b0110110011101001;
            14'h2977 	:	o_val <= 16'b0110110011101011;
            14'h2978 	:	o_val <= 16'b0110110011101100;
            14'h2979 	:	o_val <= 16'b0110110011101110;
            14'h297a 	:	o_val <= 16'b0110110011110000;
            14'h297b 	:	o_val <= 16'b0110110011110001;
            14'h297c 	:	o_val <= 16'b0110110011110011;
            14'h297d 	:	o_val <= 16'b0110110011110101;
            14'h297e 	:	o_val <= 16'b0110110011110110;
            14'h297f 	:	o_val <= 16'b0110110011111000;
            14'h2980 	:	o_val <= 16'b0110110011111010;
            14'h2981 	:	o_val <= 16'b0110110011111011;
            14'h2982 	:	o_val <= 16'b0110110011111101;
            14'h2983 	:	o_val <= 16'b0110110011111110;
            14'h2984 	:	o_val <= 16'b0110110100000000;
            14'h2985 	:	o_val <= 16'b0110110100000010;
            14'h2986 	:	o_val <= 16'b0110110100000011;
            14'h2987 	:	o_val <= 16'b0110110100000101;
            14'h2988 	:	o_val <= 16'b0110110100000111;
            14'h2989 	:	o_val <= 16'b0110110100001000;
            14'h298a 	:	o_val <= 16'b0110110100001010;
            14'h298b 	:	o_val <= 16'b0110110100001100;
            14'h298c 	:	o_val <= 16'b0110110100001101;
            14'h298d 	:	o_val <= 16'b0110110100001111;
            14'h298e 	:	o_val <= 16'b0110110100010001;
            14'h298f 	:	o_val <= 16'b0110110100010010;
            14'h2990 	:	o_val <= 16'b0110110100010100;
            14'h2991 	:	o_val <= 16'b0110110100010110;
            14'h2992 	:	o_val <= 16'b0110110100010111;
            14'h2993 	:	o_val <= 16'b0110110100011001;
            14'h2994 	:	o_val <= 16'b0110110100011010;
            14'h2995 	:	o_val <= 16'b0110110100011100;
            14'h2996 	:	o_val <= 16'b0110110100011110;
            14'h2997 	:	o_val <= 16'b0110110100011111;
            14'h2998 	:	o_val <= 16'b0110110100100001;
            14'h2999 	:	o_val <= 16'b0110110100100011;
            14'h299a 	:	o_val <= 16'b0110110100100100;
            14'h299b 	:	o_val <= 16'b0110110100100110;
            14'h299c 	:	o_val <= 16'b0110110100101000;
            14'h299d 	:	o_val <= 16'b0110110100101001;
            14'h299e 	:	o_val <= 16'b0110110100101011;
            14'h299f 	:	o_val <= 16'b0110110100101100;
            14'h29a0 	:	o_val <= 16'b0110110100101110;
            14'h29a1 	:	o_val <= 16'b0110110100110000;
            14'h29a2 	:	o_val <= 16'b0110110100110001;
            14'h29a3 	:	o_val <= 16'b0110110100110011;
            14'h29a4 	:	o_val <= 16'b0110110100110101;
            14'h29a5 	:	o_val <= 16'b0110110100110110;
            14'h29a6 	:	o_val <= 16'b0110110100111000;
            14'h29a7 	:	o_val <= 16'b0110110100111010;
            14'h29a8 	:	o_val <= 16'b0110110100111011;
            14'h29a9 	:	o_val <= 16'b0110110100111101;
            14'h29aa 	:	o_val <= 16'b0110110100111111;
            14'h29ab 	:	o_val <= 16'b0110110101000000;
            14'h29ac 	:	o_val <= 16'b0110110101000010;
            14'h29ad 	:	o_val <= 16'b0110110101000011;
            14'h29ae 	:	o_val <= 16'b0110110101000101;
            14'h29af 	:	o_val <= 16'b0110110101000111;
            14'h29b0 	:	o_val <= 16'b0110110101001000;
            14'h29b1 	:	o_val <= 16'b0110110101001010;
            14'h29b2 	:	o_val <= 16'b0110110101001100;
            14'h29b3 	:	o_val <= 16'b0110110101001101;
            14'h29b4 	:	o_val <= 16'b0110110101001111;
            14'h29b5 	:	o_val <= 16'b0110110101010001;
            14'h29b6 	:	o_val <= 16'b0110110101010010;
            14'h29b7 	:	o_val <= 16'b0110110101010100;
            14'h29b8 	:	o_val <= 16'b0110110101010101;
            14'h29b9 	:	o_val <= 16'b0110110101010111;
            14'h29ba 	:	o_val <= 16'b0110110101011001;
            14'h29bb 	:	o_val <= 16'b0110110101011010;
            14'h29bc 	:	o_val <= 16'b0110110101011100;
            14'h29bd 	:	o_val <= 16'b0110110101011110;
            14'h29be 	:	o_val <= 16'b0110110101011111;
            14'h29bf 	:	o_val <= 16'b0110110101100001;
            14'h29c0 	:	o_val <= 16'b0110110101100010;
            14'h29c1 	:	o_val <= 16'b0110110101100100;
            14'h29c2 	:	o_val <= 16'b0110110101100110;
            14'h29c3 	:	o_val <= 16'b0110110101100111;
            14'h29c4 	:	o_val <= 16'b0110110101101001;
            14'h29c5 	:	o_val <= 16'b0110110101101011;
            14'h29c6 	:	o_val <= 16'b0110110101101100;
            14'h29c7 	:	o_val <= 16'b0110110101101110;
            14'h29c8 	:	o_val <= 16'b0110110101110000;
            14'h29c9 	:	o_val <= 16'b0110110101110001;
            14'h29ca 	:	o_val <= 16'b0110110101110011;
            14'h29cb 	:	o_val <= 16'b0110110101110100;
            14'h29cc 	:	o_val <= 16'b0110110101110110;
            14'h29cd 	:	o_val <= 16'b0110110101111000;
            14'h29ce 	:	o_val <= 16'b0110110101111001;
            14'h29cf 	:	o_val <= 16'b0110110101111011;
            14'h29d0 	:	o_val <= 16'b0110110101111101;
            14'h29d1 	:	o_val <= 16'b0110110101111110;
            14'h29d2 	:	o_val <= 16'b0110110110000000;
            14'h29d3 	:	o_val <= 16'b0110110110000001;
            14'h29d4 	:	o_val <= 16'b0110110110000011;
            14'h29d5 	:	o_val <= 16'b0110110110000101;
            14'h29d6 	:	o_val <= 16'b0110110110000110;
            14'h29d7 	:	o_val <= 16'b0110110110001000;
            14'h29d8 	:	o_val <= 16'b0110110110001010;
            14'h29d9 	:	o_val <= 16'b0110110110001011;
            14'h29da 	:	o_val <= 16'b0110110110001101;
            14'h29db 	:	o_val <= 16'b0110110110001110;
            14'h29dc 	:	o_val <= 16'b0110110110010000;
            14'h29dd 	:	o_val <= 16'b0110110110010010;
            14'h29de 	:	o_val <= 16'b0110110110010011;
            14'h29df 	:	o_val <= 16'b0110110110010101;
            14'h29e0 	:	o_val <= 16'b0110110110010111;
            14'h29e1 	:	o_val <= 16'b0110110110011000;
            14'h29e2 	:	o_val <= 16'b0110110110011010;
            14'h29e3 	:	o_val <= 16'b0110110110011011;
            14'h29e4 	:	o_val <= 16'b0110110110011101;
            14'h29e5 	:	o_val <= 16'b0110110110011111;
            14'h29e6 	:	o_val <= 16'b0110110110100000;
            14'h29e7 	:	o_val <= 16'b0110110110100010;
            14'h29e8 	:	o_val <= 16'b0110110110100100;
            14'h29e9 	:	o_val <= 16'b0110110110100101;
            14'h29ea 	:	o_val <= 16'b0110110110100111;
            14'h29eb 	:	o_val <= 16'b0110110110101000;
            14'h29ec 	:	o_val <= 16'b0110110110101010;
            14'h29ed 	:	o_val <= 16'b0110110110101100;
            14'h29ee 	:	o_val <= 16'b0110110110101101;
            14'h29ef 	:	o_val <= 16'b0110110110101111;
            14'h29f0 	:	o_val <= 16'b0110110110110000;
            14'h29f1 	:	o_val <= 16'b0110110110110010;
            14'h29f2 	:	o_val <= 16'b0110110110110100;
            14'h29f3 	:	o_val <= 16'b0110110110110101;
            14'h29f4 	:	o_val <= 16'b0110110110110111;
            14'h29f5 	:	o_val <= 16'b0110110110111001;
            14'h29f6 	:	o_val <= 16'b0110110110111010;
            14'h29f7 	:	o_val <= 16'b0110110110111100;
            14'h29f8 	:	o_val <= 16'b0110110110111101;
            14'h29f9 	:	o_val <= 16'b0110110110111111;
            14'h29fa 	:	o_val <= 16'b0110110111000001;
            14'h29fb 	:	o_val <= 16'b0110110111000010;
            14'h29fc 	:	o_val <= 16'b0110110111000100;
            14'h29fd 	:	o_val <= 16'b0110110111000110;
            14'h29fe 	:	o_val <= 16'b0110110111000111;
            14'h29ff 	:	o_val <= 16'b0110110111001001;
            14'h2a00 	:	o_val <= 16'b0110110111001010;
            14'h2a01 	:	o_val <= 16'b0110110111001100;
            14'h2a02 	:	o_val <= 16'b0110110111001110;
            14'h2a03 	:	o_val <= 16'b0110110111001111;
            14'h2a04 	:	o_val <= 16'b0110110111010001;
            14'h2a05 	:	o_val <= 16'b0110110111010010;
            14'h2a06 	:	o_val <= 16'b0110110111010100;
            14'h2a07 	:	o_val <= 16'b0110110111010110;
            14'h2a08 	:	o_val <= 16'b0110110111010111;
            14'h2a09 	:	o_val <= 16'b0110110111011001;
            14'h2a0a 	:	o_val <= 16'b0110110111011010;
            14'h2a0b 	:	o_val <= 16'b0110110111011100;
            14'h2a0c 	:	o_val <= 16'b0110110111011110;
            14'h2a0d 	:	o_val <= 16'b0110110111011111;
            14'h2a0e 	:	o_val <= 16'b0110110111100001;
            14'h2a0f 	:	o_val <= 16'b0110110111100011;
            14'h2a10 	:	o_val <= 16'b0110110111100100;
            14'h2a11 	:	o_val <= 16'b0110110111100110;
            14'h2a12 	:	o_val <= 16'b0110110111100111;
            14'h2a13 	:	o_val <= 16'b0110110111101001;
            14'h2a14 	:	o_val <= 16'b0110110111101011;
            14'h2a15 	:	o_val <= 16'b0110110111101100;
            14'h2a16 	:	o_val <= 16'b0110110111101110;
            14'h2a17 	:	o_val <= 16'b0110110111101111;
            14'h2a18 	:	o_val <= 16'b0110110111110001;
            14'h2a19 	:	o_val <= 16'b0110110111110011;
            14'h2a1a 	:	o_val <= 16'b0110110111110100;
            14'h2a1b 	:	o_val <= 16'b0110110111110110;
            14'h2a1c 	:	o_val <= 16'b0110110111110111;
            14'h2a1d 	:	o_val <= 16'b0110110111111001;
            14'h2a1e 	:	o_val <= 16'b0110110111111011;
            14'h2a1f 	:	o_val <= 16'b0110110111111100;
            14'h2a20 	:	o_val <= 16'b0110110111111110;
            14'h2a21 	:	o_val <= 16'b0110111000000000;
            14'h2a22 	:	o_val <= 16'b0110111000000001;
            14'h2a23 	:	o_val <= 16'b0110111000000011;
            14'h2a24 	:	o_val <= 16'b0110111000000100;
            14'h2a25 	:	o_val <= 16'b0110111000000110;
            14'h2a26 	:	o_val <= 16'b0110111000001000;
            14'h2a27 	:	o_val <= 16'b0110111000001001;
            14'h2a28 	:	o_val <= 16'b0110111000001011;
            14'h2a29 	:	o_val <= 16'b0110111000001100;
            14'h2a2a 	:	o_val <= 16'b0110111000001110;
            14'h2a2b 	:	o_val <= 16'b0110111000010000;
            14'h2a2c 	:	o_val <= 16'b0110111000010001;
            14'h2a2d 	:	o_val <= 16'b0110111000010011;
            14'h2a2e 	:	o_val <= 16'b0110111000010100;
            14'h2a2f 	:	o_val <= 16'b0110111000010110;
            14'h2a30 	:	o_val <= 16'b0110111000011000;
            14'h2a31 	:	o_val <= 16'b0110111000011001;
            14'h2a32 	:	o_val <= 16'b0110111000011011;
            14'h2a33 	:	o_val <= 16'b0110111000011100;
            14'h2a34 	:	o_val <= 16'b0110111000011110;
            14'h2a35 	:	o_val <= 16'b0110111000100000;
            14'h2a36 	:	o_val <= 16'b0110111000100001;
            14'h2a37 	:	o_val <= 16'b0110111000100011;
            14'h2a38 	:	o_val <= 16'b0110111000100100;
            14'h2a39 	:	o_val <= 16'b0110111000100110;
            14'h2a3a 	:	o_val <= 16'b0110111000101000;
            14'h2a3b 	:	o_val <= 16'b0110111000101001;
            14'h2a3c 	:	o_val <= 16'b0110111000101011;
            14'h2a3d 	:	o_val <= 16'b0110111000101100;
            14'h2a3e 	:	o_val <= 16'b0110111000101110;
            14'h2a3f 	:	o_val <= 16'b0110111000110000;
            14'h2a40 	:	o_val <= 16'b0110111000110001;
            14'h2a41 	:	o_val <= 16'b0110111000110011;
            14'h2a42 	:	o_val <= 16'b0110111000110100;
            14'h2a43 	:	o_val <= 16'b0110111000110110;
            14'h2a44 	:	o_val <= 16'b0110111000111000;
            14'h2a45 	:	o_val <= 16'b0110111000111001;
            14'h2a46 	:	o_val <= 16'b0110111000111011;
            14'h2a47 	:	o_val <= 16'b0110111000111100;
            14'h2a48 	:	o_val <= 16'b0110111000111110;
            14'h2a49 	:	o_val <= 16'b0110111001000000;
            14'h2a4a 	:	o_val <= 16'b0110111001000001;
            14'h2a4b 	:	o_val <= 16'b0110111001000011;
            14'h2a4c 	:	o_val <= 16'b0110111001000100;
            14'h2a4d 	:	o_val <= 16'b0110111001000110;
            14'h2a4e 	:	o_val <= 16'b0110111001001000;
            14'h2a4f 	:	o_val <= 16'b0110111001001001;
            14'h2a50 	:	o_val <= 16'b0110111001001011;
            14'h2a51 	:	o_val <= 16'b0110111001001100;
            14'h2a52 	:	o_val <= 16'b0110111001001110;
            14'h2a53 	:	o_val <= 16'b0110111001010000;
            14'h2a54 	:	o_val <= 16'b0110111001010001;
            14'h2a55 	:	o_val <= 16'b0110111001010011;
            14'h2a56 	:	o_val <= 16'b0110111001010100;
            14'h2a57 	:	o_val <= 16'b0110111001010110;
            14'h2a58 	:	o_val <= 16'b0110111001010111;
            14'h2a59 	:	o_val <= 16'b0110111001011001;
            14'h2a5a 	:	o_val <= 16'b0110111001011011;
            14'h2a5b 	:	o_val <= 16'b0110111001011100;
            14'h2a5c 	:	o_val <= 16'b0110111001011110;
            14'h2a5d 	:	o_val <= 16'b0110111001011111;
            14'h2a5e 	:	o_val <= 16'b0110111001100001;
            14'h2a5f 	:	o_val <= 16'b0110111001100011;
            14'h2a60 	:	o_val <= 16'b0110111001100100;
            14'h2a61 	:	o_val <= 16'b0110111001100110;
            14'h2a62 	:	o_val <= 16'b0110111001100111;
            14'h2a63 	:	o_val <= 16'b0110111001101001;
            14'h2a64 	:	o_val <= 16'b0110111001101011;
            14'h2a65 	:	o_val <= 16'b0110111001101100;
            14'h2a66 	:	o_val <= 16'b0110111001101110;
            14'h2a67 	:	o_val <= 16'b0110111001101111;
            14'h2a68 	:	o_val <= 16'b0110111001110001;
            14'h2a69 	:	o_val <= 16'b0110111001110011;
            14'h2a6a 	:	o_val <= 16'b0110111001110100;
            14'h2a6b 	:	o_val <= 16'b0110111001110110;
            14'h2a6c 	:	o_val <= 16'b0110111001110111;
            14'h2a6d 	:	o_val <= 16'b0110111001111001;
            14'h2a6e 	:	o_val <= 16'b0110111001111010;
            14'h2a6f 	:	o_val <= 16'b0110111001111100;
            14'h2a70 	:	o_val <= 16'b0110111001111110;
            14'h2a71 	:	o_val <= 16'b0110111001111111;
            14'h2a72 	:	o_val <= 16'b0110111010000001;
            14'h2a73 	:	o_val <= 16'b0110111010000010;
            14'h2a74 	:	o_val <= 16'b0110111010000100;
            14'h2a75 	:	o_val <= 16'b0110111010000110;
            14'h2a76 	:	o_val <= 16'b0110111010000111;
            14'h2a77 	:	o_val <= 16'b0110111010001001;
            14'h2a78 	:	o_val <= 16'b0110111010001010;
            14'h2a79 	:	o_val <= 16'b0110111010001100;
            14'h2a7a 	:	o_val <= 16'b0110111010001101;
            14'h2a7b 	:	o_val <= 16'b0110111010001111;
            14'h2a7c 	:	o_val <= 16'b0110111010010001;
            14'h2a7d 	:	o_val <= 16'b0110111010010010;
            14'h2a7e 	:	o_val <= 16'b0110111010010100;
            14'h2a7f 	:	o_val <= 16'b0110111010010101;
            14'h2a80 	:	o_val <= 16'b0110111010010111;
            14'h2a81 	:	o_val <= 16'b0110111010011001;
            14'h2a82 	:	o_val <= 16'b0110111010011010;
            14'h2a83 	:	o_val <= 16'b0110111010011100;
            14'h2a84 	:	o_val <= 16'b0110111010011101;
            14'h2a85 	:	o_val <= 16'b0110111010011111;
            14'h2a86 	:	o_val <= 16'b0110111010100000;
            14'h2a87 	:	o_val <= 16'b0110111010100010;
            14'h2a88 	:	o_val <= 16'b0110111010100100;
            14'h2a89 	:	o_val <= 16'b0110111010100101;
            14'h2a8a 	:	o_val <= 16'b0110111010100111;
            14'h2a8b 	:	o_val <= 16'b0110111010101000;
            14'h2a8c 	:	o_val <= 16'b0110111010101010;
            14'h2a8d 	:	o_val <= 16'b0110111010101011;
            14'h2a8e 	:	o_val <= 16'b0110111010101101;
            14'h2a8f 	:	o_val <= 16'b0110111010101111;
            14'h2a90 	:	o_val <= 16'b0110111010110000;
            14'h2a91 	:	o_val <= 16'b0110111010110010;
            14'h2a92 	:	o_val <= 16'b0110111010110011;
            14'h2a93 	:	o_val <= 16'b0110111010110101;
            14'h2a94 	:	o_val <= 16'b0110111010110111;
            14'h2a95 	:	o_val <= 16'b0110111010111000;
            14'h2a96 	:	o_val <= 16'b0110111010111010;
            14'h2a97 	:	o_val <= 16'b0110111010111011;
            14'h2a98 	:	o_val <= 16'b0110111010111101;
            14'h2a99 	:	o_val <= 16'b0110111010111110;
            14'h2a9a 	:	o_val <= 16'b0110111011000000;
            14'h2a9b 	:	o_val <= 16'b0110111011000010;
            14'h2a9c 	:	o_val <= 16'b0110111011000011;
            14'h2a9d 	:	o_val <= 16'b0110111011000101;
            14'h2a9e 	:	o_val <= 16'b0110111011000110;
            14'h2a9f 	:	o_val <= 16'b0110111011001000;
            14'h2aa0 	:	o_val <= 16'b0110111011001001;
            14'h2aa1 	:	o_val <= 16'b0110111011001011;
            14'h2aa2 	:	o_val <= 16'b0110111011001101;
            14'h2aa3 	:	o_val <= 16'b0110111011001110;
            14'h2aa4 	:	o_val <= 16'b0110111011010000;
            14'h2aa5 	:	o_val <= 16'b0110111011010001;
            14'h2aa6 	:	o_val <= 16'b0110111011010011;
            14'h2aa7 	:	o_val <= 16'b0110111011010100;
            14'h2aa8 	:	o_val <= 16'b0110111011010110;
            14'h2aa9 	:	o_val <= 16'b0110111011011000;
            14'h2aaa 	:	o_val <= 16'b0110111011011001;
            14'h2aab 	:	o_val <= 16'b0110111011011011;
            14'h2aac 	:	o_val <= 16'b0110111011011100;
            14'h2aad 	:	o_val <= 16'b0110111011011110;
            14'h2aae 	:	o_val <= 16'b0110111011011111;
            14'h2aaf 	:	o_val <= 16'b0110111011100001;
            14'h2ab0 	:	o_val <= 16'b0110111011100011;
            14'h2ab1 	:	o_val <= 16'b0110111011100100;
            14'h2ab2 	:	o_val <= 16'b0110111011100110;
            14'h2ab3 	:	o_val <= 16'b0110111011100111;
            14'h2ab4 	:	o_val <= 16'b0110111011101001;
            14'h2ab5 	:	o_val <= 16'b0110111011101010;
            14'h2ab6 	:	o_val <= 16'b0110111011101100;
            14'h2ab7 	:	o_val <= 16'b0110111011101110;
            14'h2ab8 	:	o_val <= 16'b0110111011101111;
            14'h2ab9 	:	o_val <= 16'b0110111011110001;
            14'h2aba 	:	o_val <= 16'b0110111011110010;
            14'h2abb 	:	o_val <= 16'b0110111011110100;
            14'h2abc 	:	o_val <= 16'b0110111011110101;
            14'h2abd 	:	o_val <= 16'b0110111011110111;
            14'h2abe 	:	o_val <= 16'b0110111011111001;
            14'h2abf 	:	o_val <= 16'b0110111011111010;
            14'h2ac0 	:	o_val <= 16'b0110111011111100;
            14'h2ac1 	:	o_val <= 16'b0110111011111101;
            14'h2ac2 	:	o_val <= 16'b0110111011111111;
            14'h2ac3 	:	o_val <= 16'b0110111100000000;
            14'h2ac4 	:	o_val <= 16'b0110111100000010;
            14'h2ac5 	:	o_val <= 16'b0110111100000011;
            14'h2ac6 	:	o_val <= 16'b0110111100000101;
            14'h2ac7 	:	o_val <= 16'b0110111100000111;
            14'h2ac8 	:	o_val <= 16'b0110111100001000;
            14'h2ac9 	:	o_val <= 16'b0110111100001010;
            14'h2aca 	:	o_val <= 16'b0110111100001011;
            14'h2acb 	:	o_val <= 16'b0110111100001101;
            14'h2acc 	:	o_val <= 16'b0110111100001110;
            14'h2acd 	:	o_val <= 16'b0110111100010000;
            14'h2ace 	:	o_val <= 16'b0110111100010010;
            14'h2acf 	:	o_val <= 16'b0110111100010011;
            14'h2ad0 	:	o_val <= 16'b0110111100010101;
            14'h2ad1 	:	o_val <= 16'b0110111100010110;
            14'h2ad2 	:	o_val <= 16'b0110111100011000;
            14'h2ad3 	:	o_val <= 16'b0110111100011001;
            14'h2ad4 	:	o_val <= 16'b0110111100011011;
            14'h2ad5 	:	o_val <= 16'b0110111100011100;
            14'h2ad6 	:	o_val <= 16'b0110111100011110;
            14'h2ad7 	:	o_val <= 16'b0110111100100000;
            14'h2ad8 	:	o_val <= 16'b0110111100100001;
            14'h2ad9 	:	o_val <= 16'b0110111100100011;
            14'h2ada 	:	o_val <= 16'b0110111100100100;
            14'h2adb 	:	o_val <= 16'b0110111100100110;
            14'h2adc 	:	o_val <= 16'b0110111100100111;
            14'h2add 	:	o_val <= 16'b0110111100101001;
            14'h2ade 	:	o_val <= 16'b0110111100101010;
            14'h2adf 	:	o_val <= 16'b0110111100101100;
            14'h2ae0 	:	o_val <= 16'b0110111100101110;
            14'h2ae1 	:	o_val <= 16'b0110111100101111;
            14'h2ae2 	:	o_val <= 16'b0110111100110001;
            14'h2ae3 	:	o_val <= 16'b0110111100110010;
            14'h2ae4 	:	o_val <= 16'b0110111100110100;
            14'h2ae5 	:	o_val <= 16'b0110111100110101;
            14'h2ae6 	:	o_val <= 16'b0110111100110111;
            14'h2ae7 	:	o_val <= 16'b0110111100111000;
            14'h2ae8 	:	o_val <= 16'b0110111100111010;
            14'h2ae9 	:	o_val <= 16'b0110111100111100;
            14'h2aea 	:	o_val <= 16'b0110111100111101;
            14'h2aeb 	:	o_val <= 16'b0110111100111111;
            14'h2aec 	:	o_val <= 16'b0110111101000000;
            14'h2aed 	:	o_val <= 16'b0110111101000010;
            14'h2aee 	:	o_val <= 16'b0110111101000011;
            14'h2aef 	:	o_val <= 16'b0110111101000101;
            14'h2af0 	:	o_val <= 16'b0110111101000110;
            14'h2af1 	:	o_val <= 16'b0110111101001000;
            14'h2af2 	:	o_val <= 16'b0110111101001010;
            14'h2af3 	:	o_val <= 16'b0110111101001011;
            14'h2af4 	:	o_val <= 16'b0110111101001101;
            14'h2af5 	:	o_val <= 16'b0110111101001110;
            14'h2af6 	:	o_val <= 16'b0110111101010000;
            14'h2af7 	:	o_val <= 16'b0110111101010001;
            14'h2af8 	:	o_val <= 16'b0110111101010011;
            14'h2af9 	:	o_val <= 16'b0110111101010100;
            14'h2afa 	:	o_val <= 16'b0110111101010110;
            14'h2afb 	:	o_val <= 16'b0110111101011000;
            14'h2afc 	:	o_val <= 16'b0110111101011001;
            14'h2afd 	:	o_val <= 16'b0110111101011011;
            14'h2afe 	:	o_val <= 16'b0110111101011100;
            14'h2aff 	:	o_val <= 16'b0110111101011110;
            14'h2b00 	:	o_val <= 16'b0110111101011111;
            14'h2b01 	:	o_val <= 16'b0110111101100001;
            14'h2b02 	:	o_val <= 16'b0110111101100010;
            14'h2b03 	:	o_val <= 16'b0110111101100100;
            14'h2b04 	:	o_val <= 16'b0110111101100101;
            14'h2b05 	:	o_val <= 16'b0110111101100111;
            14'h2b06 	:	o_val <= 16'b0110111101101001;
            14'h2b07 	:	o_val <= 16'b0110111101101010;
            14'h2b08 	:	o_val <= 16'b0110111101101100;
            14'h2b09 	:	o_val <= 16'b0110111101101101;
            14'h2b0a 	:	o_val <= 16'b0110111101101111;
            14'h2b0b 	:	o_val <= 16'b0110111101110000;
            14'h2b0c 	:	o_val <= 16'b0110111101110010;
            14'h2b0d 	:	o_val <= 16'b0110111101110011;
            14'h2b0e 	:	o_val <= 16'b0110111101110101;
            14'h2b0f 	:	o_val <= 16'b0110111101110110;
            14'h2b10 	:	o_val <= 16'b0110111101111000;
            14'h2b11 	:	o_val <= 16'b0110111101111010;
            14'h2b12 	:	o_val <= 16'b0110111101111011;
            14'h2b13 	:	o_val <= 16'b0110111101111101;
            14'h2b14 	:	o_val <= 16'b0110111101111110;
            14'h2b15 	:	o_val <= 16'b0110111110000000;
            14'h2b16 	:	o_val <= 16'b0110111110000001;
            14'h2b17 	:	o_val <= 16'b0110111110000011;
            14'h2b18 	:	o_val <= 16'b0110111110000100;
            14'h2b19 	:	o_val <= 16'b0110111110000110;
            14'h2b1a 	:	o_val <= 16'b0110111110000111;
            14'h2b1b 	:	o_val <= 16'b0110111110001001;
            14'h2b1c 	:	o_val <= 16'b0110111110001011;
            14'h2b1d 	:	o_val <= 16'b0110111110001100;
            14'h2b1e 	:	o_val <= 16'b0110111110001110;
            14'h2b1f 	:	o_val <= 16'b0110111110001111;
            14'h2b20 	:	o_val <= 16'b0110111110010001;
            14'h2b21 	:	o_val <= 16'b0110111110010010;
            14'h2b22 	:	o_val <= 16'b0110111110010100;
            14'h2b23 	:	o_val <= 16'b0110111110010101;
            14'h2b24 	:	o_val <= 16'b0110111110010111;
            14'h2b25 	:	o_val <= 16'b0110111110011000;
            14'h2b26 	:	o_val <= 16'b0110111110011010;
            14'h2b27 	:	o_val <= 16'b0110111110011011;
            14'h2b28 	:	o_val <= 16'b0110111110011101;
            14'h2b29 	:	o_val <= 16'b0110111110011111;
            14'h2b2a 	:	o_val <= 16'b0110111110100000;
            14'h2b2b 	:	o_val <= 16'b0110111110100010;
            14'h2b2c 	:	o_val <= 16'b0110111110100011;
            14'h2b2d 	:	o_val <= 16'b0110111110100101;
            14'h2b2e 	:	o_val <= 16'b0110111110100110;
            14'h2b2f 	:	o_val <= 16'b0110111110101000;
            14'h2b30 	:	o_val <= 16'b0110111110101001;
            14'h2b31 	:	o_val <= 16'b0110111110101011;
            14'h2b32 	:	o_val <= 16'b0110111110101100;
            14'h2b33 	:	o_val <= 16'b0110111110101110;
            14'h2b34 	:	o_val <= 16'b0110111110101111;
            14'h2b35 	:	o_val <= 16'b0110111110110001;
            14'h2b36 	:	o_val <= 16'b0110111110110011;
            14'h2b37 	:	o_val <= 16'b0110111110110100;
            14'h2b38 	:	o_val <= 16'b0110111110110110;
            14'h2b39 	:	o_val <= 16'b0110111110110111;
            14'h2b3a 	:	o_val <= 16'b0110111110111001;
            14'h2b3b 	:	o_val <= 16'b0110111110111010;
            14'h2b3c 	:	o_val <= 16'b0110111110111100;
            14'h2b3d 	:	o_val <= 16'b0110111110111101;
            14'h2b3e 	:	o_val <= 16'b0110111110111111;
            14'h2b3f 	:	o_val <= 16'b0110111111000000;
            14'h2b40 	:	o_val <= 16'b0110111111000010;
            14'h2b41 	:	o_val <= 16'b0110111111000011;
            14'h2b42 	:	o_val <= 16'b0110111111000101;
            14'h2b43 	:	o_val <= 16'b0110111111000110;
            14'h2b44 	:	o_val <= 16'b0110111111001000;
            14'h2b45 	:	o_val <= 16'b0110111111001001;
            14'h2b46 	:	o_val <= 16'b0110111111001011;
            14'h2b47 	:	o_val <= 16'b0110111111001101;
            14'h2b48 	:	o_val <= 16'b0110111111001110;
            14'h2b49 	:	o_val <= 16'b0110111111010000;
            14'h2b4a 	:	o_val <= 16'b0110111111010001;
            14'h2b4b 	:	o_val <= 16'b0110111111010011;
            14'h2b4c 	:	o_val <= 16'b0110111111010100;
            14'h2b4d 	:	o_val <= 16'b0110111111010110;
            14'h2b4e 	:	o_val <= 16'b0110111111010111;
            14'h2b4f 	:	o_val <= 16'b0110111111011001;
            14'h2b50 	:	o_val <= 16'b0110111111011010;
            14'h2b51 	:	o_val <= 16'b0110111111011100;
            14'h2b52 	:	o_val <= 16'b0110111111011101;
            14'h2b53 	:	o_val <= 16'b0110111111011111;
            14'h2b54 	:	o_val <= 16'b0110111111100000;
            14'h2b55 	:	o_val <= 16'b0110111111100010;
            14'h2b56 	:	o_val <= 16'b0110111111100011;
            14'h2b57 	:	o_val <= 16'b0110111111100101;
            14'h2b58 	:	o_val <= 16'b0110111111100111;
            14'h2b59 	:	o_val <= 16'b0110111111101000;
            14'h2b5a 	:	o_val <= 16'b0110111111101010;
            14'h2b5b 	:	o_val <= 16'b0110111111101011;
            14'h2b5c 	:	o_val <= 16'b0110111111101101;
            14'h2b5d 	:	o_val <= 16'b0110111111101110;
            14'h2b5e 	:	o_val <= 16'b0110111111110000;
            14'h2b5f 	:	o_val <= 16'b0110111111110001;
            14'h2b60 	:	o_val <= 16'b0110111111110011;
            14'h2b61 	:	o_val <= 16'b0110111111110100;
            14'h2b62 	:	o_val <= 16'b0110111111110110;
            14'h2b63 	:	o_val <= 16'b0110111111110111;
            14'h2b64 	:	o_val <= 16'b0110111111111001;
            14'h2b65 	:	o_val <= 16'b0110111111111010;
            14'h2b66 	:	o_val <= 16'b0110111111111100;
            14'h2b67 	:	o_val <= 16'b0110111111111101;
            14'h2b68 	:	o_val <= 16'b0110111111111111;
            14'h2b69 	:	o_val <= 16'b0111000000000000;
            14'h2b6a 	:	o_val <= 16'b0111000000000010;
            14'h2b6b 	:	o_val <= 16'b0111000000000011;
            14'h2b6c 	:	o_val <= 16'b0111000000000101;
            14'h2b6d 	:	o_val <= 16'b0111000000000110;
            14'h2b6e 	:	o_val <= 16'b0111000000001000;
            14'h2b6f 	:	o_val <= 16'b0111000000001010;
            14'h2b70 	:	o_val <= 16'b0111000000001011;
            14'h2b71 	:	o_val <= 16'b0111000000001101;
            14'h2b72 	:	o_val <= 16'b0111000000001110;
            14'h2b73 	:	o_val <= 16'b0111000000010000;
            14'h2b74 	:	o_val <= 16'b0111000000010001;
            14'h2b75 	:	o_val <= 16'b0111000000010011;
            14'h2b76 	:	o_val <= 16'b0111000000010100;
            14'h2b77 	:	o_val <= 16'b0111000000010110;
            14'h2b78 	:	o_val <= 16'b0111000000010111;
            14'h2b79 	:	o_val <= 16'b0111000000011001;
            14'h2b7a 	:	o_val <= 16'b0111000000011010;
            14'h2b7b 	:	o_val <= 16'b0111000000011100;
            14'h2b7c 	:	o_val <= 16'b0111000000011101;
            14'h2b7d 	:	o_val <= 16'b0111000000011111;
            14'h2b7e 	:	o_val <= 16'b0111000000100000;
            14'h2b7f 	:	o_val <= 16'b0111000000100010;
            14'h2b80 	:	o_val <= 16'b0111000000100011;
            14'h2b81 	:	o_val <= 16'b0111000000100101;
            14'h2b82 	:	o_val <= 16'b0111000000100110;
            14'h2b83 	:	o_val <= 16'b0111000000101000;
            14'h2b84 	:	o_val <= 16'b0111000000101001;
            14'h2b85 	:	o_val <= 16'b0111000000101011;
            14'h2b86 	:	o_val <= 16'b0111000000101100;
            14'h2b87 	:	o_val <= 16'b0111000000101110;
            14'h2b88 	:	o_val <= 16'b0111000000101111;
            14'h2b89 	:	o_val <= 16'b0111000000110001;
            14'h2b8a 	:	o_val <= 16'b0111000000110010;
            14'h2b8b 	:	o_val <= 16'b0111000000110100;
            14'h2b8c 	:	o_val <= 16'b0111000000110101;
            14'h2b8d 	:	o_val <= 16'b0111000000110111;
            14'h2b8e 	:	o_val <= 16'b0111000000111001;
            14'h2b8f 	:	o_val <= 16'b0111000000111010;
            14'h2b90 	:	o_val <= 16'b0111000000111100;
            14'h2b91 	:	o_val <= 16'b0111000000111101;
            14'h2b92 	:	o_val <= 16'b0111000000111111;
            14'h2b93 	:	o_val <= 16'b0111000001000000;
            14'h2b94 	:	o_val <= 16'b0111000001000010;
            14'h2b95 	:	o_val <= 16'b0111000001000011;
            14'h2b96 	:	o_val <= 16'b0111000001000101;
            14'h2b97 	:	o_val <= 16'b0111000001000110;
            14'h2b98 	:	o_val <= 16'b0111000001001000;
            14'h2b99 	:	o_val <= 16'b0111000001001001;
            14'h2b9a 	:	o_val <= 16'b0111000001001011;
            14'h2b9b 	:	o_val <= 16'b0111000001001100;
            14'h2b9c 	:	o_val <= 16'b0111000001001110;
            14'h2b9d 	:	o_val <= 16'b0111000001001111;
            14'h2b9e 	:	o_val <= 16'b0111000001010001;
            14'h2b9f 	:	o_val <= 16'b0111000001010010;
            14'h2ba0 	:	o_val <= 16'b0111000001010100;
            14'h2ba1 	:	o_val <= 16'b0111000001010101;
            14'h2ba2 	:	o_val <= 16'b0111000001010111;
            14'h2ba3 	:	o_val <= 16'b0111000001011000;
            14'h2ba4 	:	o_val <= 16'b0111000001011010;
            14'h2ba5 	:	o_val <= 16'b0111000001011011;
            14'h2ba6 	:	o_val <= 16'b0111000001011101;
            14'h2ba7 	:	o_val <= 16'b0111000001011110;
            14'h2ba8 	:	o_val <= 16'b0111000001100000;
            14'h2ba9 	:	o_val <= 16'b0111000001100001;
            14'h2baa 	:	o_val <= 16'b0111000001100011;
            14'h2bab 	:	o_val <= 16'b0111000001100100;
            14'h2bac 	:	o_val <= 16'b0111000001100110;
            14'h2bad 	:	o_val <= 16'b0111000001100111;
            14'h2bae 	:	o_val <= 16'b0111000001101001;
            14'h2baf 	:	o_val <= 16'b0111000001101010;
            14'h2bb0 	:	o_val <= 16'b0111000001101100;
            14'h2bb1 	:	o_val <= 16'b0111000001101101;
            14'h2bb2 	:	o_val <= 16'b0111000001101111;
            14'h2bb3 	:	o_val <= 16'b0111000001110000;
            14'h2bb4 	:	o_val <= 16'b0111000001110010;
            14'h2bb5 	:	o_val <= 16'b0111000001110011;
            14'h2bb6 	:	o_val <= 16'b0111000001110101;
            14'h2bb7 	:	o_val <= 16'b0111000001110110;
            14'h2bb8 	:	o_val <= 16'b0111000001111000;
            14'h2bb9 	:	o_val <= 16'b0111000001111001;
            14'h2bba 	:	o_val <= 16'b0111000001111011;
            14'h2bbb 	:	o_val <= 16'b0111000001111100;
            14'h2bbc 	:	o_val <= 16'b0111000001111110;
            14'h2bbd 	:	o_val <= 16'b0111000001111111;
            14'h2bbe 	:	o_val <= 16'b0111000010000001;
            14'h2bbf 	:	o_val <= 16'b0111000010000010;
            14'h2bc0 	:	o_val <= 16'b0111000010000100;
            14'h2bc1 	:	o_val <= 16'b0111000010000101;
            14'h2bc2 	:	o_val <= 16'b0111000010000111;
            14'h2bc3 	:	o_val <= 16'b0111000010001000;
            14'h2bc4 	:	o_val <= 16'b0111000010001010;
            14'h2bc5 	:	o_val <= 16'b0111000010001011;
            14'h2bc6 	:	o_val <= 16'b0111000010001101;
            14'h2bc7 	:	o_val <= 16'b0111000010001110;
            14'h2bc8 	:	o_val <= 16'b0111000010010000;
            14'h2bc9 	:	o_val <= 16'b0111000010010001;
            14'h2bca 	:	o_val <= 16'b0111000010010011;
            14'h2bcb 	:	o_val <= 16'b0111000010010100;
            14'h2bcc 	:	o_val <= 16'b0111000010010110;
            14'h2bcd 	:	o_val <= 16'b0111000010010111;
            14'h2bce 	:	o_val <= 16'b0111000010011001;
            14'h2bcf 	:	o_val <= 16'b0111000010011010;
            14'h2bd0 	:	o_val <= 16'b0111000010011100;
            14'h2bd1 	:	o_val <= 16'b0111000010011101;
            14'h2bd2 	:	o_val <= 16'b0111000010011111;
            14'h2bd3 	:	o_val <= 16'b0111000010100000;
            14'h2bd4 	:	o_val <= 16'b0111000010100010;
            14'h2bd5 	:	o_val <= 16'b0111000010100011;
            14'h2bd6 	:	o_val <= 16'b0111000010100101;
            14'h2bd7 	:	o_val <= 16'b0111000010100110;
            14'h2bd8 	:	o_val <= 16'b0111000010101000;
            14'h2bd9 	:	o_val <= 16'b0111000010101001;
            14'h2bda 	:	o_val <= 16'b0111000010101011;
            14'h2bdb 	:	o_val <= 16'b0111000010101100;
            14'h2bdc 	:	o_val <= 16'b0111000010101110;
            14'h2bdd 	:	o_val <= 16'b0111000010101111;
            14'h2bde 	:	o_val <= 16'b0111000010110001;
            14'h2bdf 	:	o_val <= 16'b0111000010110010;
            14'h2be0 	:	o_val <= 16'b0111000010110100;
            14'h2be1 	:	o_val <= 16'b0111000010110101;
            14'h2be2 	:	o_val <= 16'b0111000010110110;
            14'h2be3 	:	o_val <= 16'b0111000010111000;
            14'h2be4 	:	o_val <= 16'b0111000010111001;
            14'h2be5 	:	o_val <= 16'b0111000010111011;
            14'h2be6 	:	o_val <= 16'b0111000010111100;
            14'h2be7 	:	o_val <= 16'b0111000010111110;
            14'h2be8 	:	o_val <= 16'b0111000010111111;
            14'h2be9 	:	o_val <= 16'b0111000011000001;
            14'h2bea 	:	o_val <= 16'b0111000011000010;
            14'h2beb 	:	o_val <= 16'b0111000011000100;
            14'h2bec 	:	o_val <= 16'b0111000011000101;
            14'h2bed 	:	o_val <= 16'b0111000011000111;
            14'h2bee 	:	o_val <= 16'b0111000011001000;
            14'h2bef 	:	o_val <= 16'b0111000011001010;
            14'h2bf0 	:	o_val <= 16'b0111000011001011;
            14'h2bf1 	:	o_val <= 16'b0111000011001101;
            14'h2bf2 	:	o_val <= 16'b0111000011001110;
            14'h2bf3 	:	o_val <= 16'b0111000011010000;
            14'h2bf4 	:	o_val <= 16'b0111000011010001;
            14'h2bf5 	:	o_val <= 16'b0111000011010011;
            14'h2bf6 	:	o_val <= 16'b0111000011010100;
            14'h2bf7 	:	o_val <= 16'b0111000011010110;
            14'h2bf8 	:	o_val <= 16'b0111000011010111;
            14'h2bf9 	:	o_val <= 16'b0111000011011001;
            14'h2bfa 	:	o_val <= 16'b0111000011011010;
            14'h2bfb 	:	o_val <= 16'b0111000011011100;
            14'h2bfc 	:	o_val <= 16'b0111000011011101;
            14'h2bfd 	:	o_val <= 16'b0111000011011111;
            14'h2bfe 	:	o_val <= 16'b0111000011100000;
            14'h2bff 	:	o_val <= 16'b0111000011100010;
            14'h2c00 	:	o_val <= 16'b0111000011100011;
            14'h2c01 	:	o_val <= 16'b0111000011100101;
            14'h2c02 	:	o_val <= 16'b0111000011100110;
            14'h2c03 	:	o_val <= 16'b0111000011100111;
            14'h2c04 	:	o_val <= 16'b0111000011101001;
            14'h2c05 	:	o_val <= 16'b0111000011101010;
            14'h2c06 	:	o_val <= 16'b0111000011101100;
            14'h2c07 	:	o_val <= 16'b0111000011101101;
            14'h2c08 	:	o_val <= 16'b0111000011101111;
            14'h2c09 	:	o_val <= 16'b0111000011110000;
            14'h2c0a 	:	o_val <= 16'b0111000011110010;
            14'h2c0b 	:	o_val <= 16'b0111000011110011;
            14'h2c0c 	:	o_val <= 16'b0111000011110101;
            14'h2c0d 	:	o_val <= 16'b0111000011110110;
            14'h2c0e 	:	o_val <= 16'b0111000011111000;
            14'h2c0f 	:	o_val <= 16'b0111000011111001;
            14'h2c10 	:	o_val <= 16'b0111000011111011;
            14'h2c11 	:	o_val <= 16'b0111000011111100;
            14'h2c12 	:	o_val <= 16'b0111000011111110;
            14'h2c13 	:	o_val <= 16'b0111000011111111;
            14'h2c14 	:	o_val <= 16'b0111000100000001;
            14'h2c15 	:	o_val <= 16'b0111000100000010;
            14'h2c16 	:	o_val <= 16'b0111000100000100;
            14'h2c17 	:	o_val <= 16'b0111000100000101;
            14'h2c18 	:	o_val <= 16'b0111000100000110;
            14'h2c19 	:	o_val <= 16'b0111000100001000;
            14'h2c1a 	:	o_val <= 16'b0111000100001001;
            14'h2c1b 	:	o_val <= 16'b0111000100001011;
            14'h2c1c 	:	o_val <= 16'b0111000100001100;
            14'h2c1d 	:	o_val <= 16'b0111000100001110;
            14'h2c1e 	:	o_val <= 16'b0111000100001111;
            14'h2c1f 	:	o_val <= 16'b0111000100010001;
            14'h2c20 	:	o_val <= 16'b0111000100010010;
            14'h2c21 	:	o_val <= 16'b0111000100010100;
            14'h2c22 	:	o_val <= 16'b0111000100010101;
            14'h2c23 	:	o_val <= 16'b0111000100010111;
            14'h2c24 	:	o_val <= 16'b0111000100011000;
            14'h2c25 	:	o_val <= 16'b0111000100011010;
            14'h2c26 	:	o_val <= 16'b0111000100011011;
            14'h2c27 	:	o_val <= 16'b0111000100011101;
            14'h2c28 	:	o_val <= 16'b0111000100011110;
            14'h2c29 	:	o_val <= 16'b0111000100100000;
            14'h2c2a 	:	o_val <= 16'b0111000100100001;
            14'h2c2b 	:	o_val <= 16'b0111000100100010;
            14'h2c2c 	:	o_val <= 16'b0111000100100100;
            14'h2c2d 	:	o_val <= 16'b0111000100100101;
            14'h2c2e 	:	o_val <= 16'b0111000100100111;
            14'h2c2f 	:	o_val <= 16'b0111000100101000;
            14'h2c30 	:	o_val <= 16'b0111000100101010;
            14'h2c31 	:	o_val <= 16'b0111000100101011;
            14'h2c32 	:	o_val <= 16'b0111000100101101;
            14'h2c33 	:	o_val <= 16'b0111000100101110;
            14'h2c34 	:	o_val <= 16'b0111000100110000;
            14'h2c35 	:	o_val <= 16'b0111000100110001;
            14'h2c36 	:	o_val <= 16'b0111000100110011;
            14'h2c37 	:	o_val <= 16'b0111000100110100;
            14'h2c38 	:	o_val <= 16'b0111000100110110;
            14'h2c39 	:	o_val <= 16'b0111000100110111;
            14'h2c3a 	:	o_val <= 16'b0111000100111000;
            14'h2c3b 	:	o_val <= 16'b0111000100111010;
            14'h2c3c 	:	o_val <= 16'b0111000100111011;
            14'h2c3d 	:	o_val <= 16'b0111000100111101;
            14'h2c3e 	:	o_val <= 16'b0111000100111110;
            14'h2c3f 	:	o_val <= 16'b0111000101000000;
            14'h2c40 	:	o_val <= 16'b0111000101000001;
            14'h2c41 	:	o_val <= 16'b0111000101000011;
            14'h2c42 	:	o_val <= 16'b0111000101000100;
            14'h2c43 	:	o_val <= 16'b0111000101000110;
            14'h2c44 	:	o_val <= 16'b0111000101000111;
            14'h2c45 	:	o_val <= 16'b0111000101001001;
            14'h2c46 	:	o_val <= 16'b0111000101001010;
            14'h2c47 	:	o_val <= 16'b0111000101001100;
            14'h2c48 	:	o_val <= 16'b0111000101001101;
            14'h2c49 	:	o_val <= 16'b0111000101001110;
            14'h2c4a 	:	o_val <= 16'b0111000101010000;
            14'h2c4b 	:	o_val <= 16'b0111000101010001;
            14'h2c4c 	:	o_val <= 16'b0111000101010011;
            14'h2c4d 	:	o_val <= 16'b0111000101010100;
            14'h2c4e 	:	o_val <= 16'b0111000101010110;
            14'h2c4f 	:	o_val <= 16'b0111000101010111;
            14'h2c50 	:	o_val <= 16'b0111000101011001;
            14'h2c51 	:	o_val <= 16'b0111000101011010;
            14'h2c52 	:	o_val <= 16'b0111000101011100;
            14'h2c53 	:	o_val <= 16'b0111000101011101;
            14'h2c54 	:	o_val <= 16'b0111000101011110;
            14'h2c55 	:	o_val <= 16'b0111000101100000;
            14'h2c56 	:	o_val <= 16'b0111000101100001;
            14'h2c57 	:	o_val <= 16'b0111000101100011;
            14'h2c58 	:	o_val <= 16'b0111000101100100;
            14'h2c59 	:	o_val <= 16'b0111000101100110;
            14'h2c5a 	:	o_val <= 16'b0111000101100111;
            14'h2c5b 	:	o_val <= 16'b0111000101101001;
            14'h2c5c 	:	o_val <= 16'b0111000101101010;
            14'h2c5d 	:	o_val <= 16'b0111000101101100;
            14'h2c5e 	:	o_val <= 16'b0111000101101101;
            14'h2c5f 	:	o_val <= 16'b0111000101101111;
            14'h2c60 	:	o_val <= 16'b0111000101110000;
            14'h2c61 	:	o_val <= 16'b0111000101110001;
            14'h2c62 	:	o_val <= 16'b0111000101110011;
            14'h2c63 	:	o_val <= 16'b0111000101110100;
            14'h2c64 	:	o_val <= 16'b0111000101110110;
            14'h2c65 	:	o_val <= 16'b0111000101110111;
            14'h2c66 	:	o_val <= 16'b0111000101111001;
            14'h2c67 	:	o_val <= 16'b0111000101111010;
            14'h2c68 	:	o_val <= 16'b0111000101111100;
            14'h2c69 	:	o_val <= 16'b0111000101111101;
            14'h2c6a 	:	o_val <= 16'b0111000101111111;
            14'h2c6b 	:	o_val <= 16'b0111000110000000;
            14'h2c6c 	:	o_val <= 16'b0111000110000001;
            14'h2c6d 	:	o_val <= 16'b0111000110000011;
            14'h2c6e 	:	o_val <= 16'b0111000110000100;
            14'h2c6f 	:	o_val <= 16'b0111000110000110;
            14'h2c70 	:	o_val <= 16'b0111000110000111;
            14'h2c71 	:	o_val <= 16'b0111000110001001;
            14'h2c72 	:	o_val <= 16'b0111000110001010;
            14'h2c73 	:	o_val <= 16'b0111000110001100;
            14'h2c74 	:	o_val <= 16'b0111000110001101;
            14'h2c75 	:	o_val <= 16'b0111000110001110;
            14'h2c76 	:	o_val <= 16'b0111000110010000;
            14'h2c77 	:	o_val <= 16'b0111000110010001;
            14'h2c78 	:	o_val <= 16'b0111000110010011;
            14'h2c79 	:	o_val <= 16'b0111000110010100;
            14'h2c7a 	:	o_val <= 16'b0111000110010110;
            14'h2c7b 	:	o_val <= 16'b0111000110010111;
            14'h2c7c 	:	o_val <= 16'b0111000110011001;
            14'h2c7d 	:	o_val <= 16'b0111000110011010;
            14'h2c7e 	:	o_val <= 16'b0111000110011100;
            14'h2c7f 	:	o_val <= 16'b0111000110011101;
            14'h2c80 	:	o_val <= 16'b0111000110011110;
            14'h2c81 	:	o_val <= 16'b0111000110100000;
            14'h2c82 	:	o_val <= 16'b0111000110100001;
            14'h2c83 	:	o_val <= 16'b0111000110100011;
            14'h2c84 	:	o_val <= 16'b0111000110100100;
            14'h2c85 	:	o_val <= 16'b0111000110100110;
            14'h2c86 	:	o_val <= 16'b0111000110100111;
            14'h2c87 	:	o_val <= 16'b0111000110101001;
            14'h2c88 	:	o_val <= 16'b0111000110101010;
            14'h2c89 	:	o_val <= 16'b0111000110101011;
            14'h2c8a 	:	o_val <= 16'b0111000110101101;
            14'h2c8b 	:	o_val <= 16'b0111000110101110;
            14'h2c8c 	:	o_val <= 16'b0111000110110000;
            14'h2c8d 	:	o_val <= 16'b0111000110110001;
            14'h2c8e 	:	o_val <= 16'b0111000110110011;
            14'h2c8f 	:	o_val <= 16'b0111000110110100;
            14'h2c90 	:	o_val <= 16'b0111000110110110;
            14'h2c91 	:	o_val <= 16'b0111000110110111;
            14'h2c92 	:	o_val <= 16'b0111000110111000;
            14'h2c93 	:	o_val <= 16'b0111000110111010;
            14'h2c94 	:	o_val <= 16'b0111000110111011;
            14'h2c95 	:	o_val <= 16'b0111000110111101;
            14'h2c96 	:	o_val <= 16'b0111000110111110;
            14'h2c97 	:	o_val <= 16'b0111000111000000;
            14'h2c98 	:	o_val <= 16'b0111000111000001;
            14'h2c99 	:	o_val <= 16'b0111000111000010;
            14'h2c9a 	:	o_val <= 16'b0111000111000100;
            14'h2c9b 	:	o_val <= 16'b0111000111000101;
            14'h2c9c 	:	o_val <= 16'b0111000111000111;
            14'h2c9d 	:	o_val <= 16'b0111000111001000;
            14'h2c9e 	:	o_val <= 16'b0111000111001010;
            14'h2c9f 	:	o_val <= 16'b0111000111001011;
            14'h2ca0 	:	o_val <= 16'b0111000111001101;
            14'h2ca1 	:	o_val <= 16'b0111000111001110;
            14'h2ca2 	:	o_val <= 16'b0111000111001111;
            14'h2ca3 	:	o_val <= 16'b0111000111010001;
            14'h2ca4 	:	o_val <= 16'b0111000111010010;
            14'h2ca5 	:	o_val <= 16'b0111000111010100;
            14'h2ca6 	:	o_val <= 16'b0111000111010101;
            14'h2ca7 	:	o_val <= 16'b0111000111010111;
            14'h2ca8 	:	o_val <= 16'b0111000111011000;
            14'h2ca9 	:	o_val <= 16'b0111000111011001;
            14'h2caa 	:	o_val <= 16'b0111000111011011;
            14'h2cab 	:	o_val <= 16'b0111000111011100;
            14'h2cac 	:	o_val <= 16'b0111000111011110;
            14'h2cad 	:	o_val <= 16'b0111000111011111;
            14'h2cae 	:	o_val <= 16'b0111000111100001;
            14'h2caf 	:	o_val <= 16'b0111000111100010;
            14'h2cb0 	:	o_val <= 16'b0111000111100100;
            14'h2cb1 	:	o_val <= 16'b0111000111100101;
            14'h2cb2 	:	o_val <= 16'b0111000111100110;
            14'h2cb3 	:	o_val <= 16'b0111000111101000;
            14'h2cb4 	:	o_val <= 16'b0111000111101001;
            14'h2cb5 	:	o_val <= 16'b0111000111101011;
            14'h2cb6 	:	o_val <= 16'b0111000111101100;
            14'h2cb7 	:	o_val <= 16'b0111000111101110;
            14'h2cb8 	:	o_val <= 16'b0111000111101111;
            14'h2cb9 	:	o_val <= 16'b0111000111110000;
            14'h2cba 	:	o_val <= 16'b0111000111110010;
            14'h2cbb 	:	o_val <= 16'b0111000111110011;
            14'h2cbc 	:	o_val <= 16'b0111000111110101;
            14'h2cbd 	:	o_val <= 16'b0111000111110110;
            14'h2cbe 	:	o_val <= 16'b0111000111111000;
            14'h2cbf 	:	o_val <= 16'b0111000111111001;
            14'h2cc0 	:	o_val <= 16'b0111000111111010;
            14'h2cc1 	:	o_val <= 16'b0111000111111100;
            14'h2cc2 	:	o_val <= 16'b0111000111111101;
            14'h2cc3 	:	o_val <= 16'b0111000111111111;
            14'h2cc4 	:	o_val <= 16'b0111001000000000;
            14'h2cc5 	:	o_val <= 16'b0111001000000010;
            14'h2cc6 	:	o_val <= 16'b0111001000000011;
            14'h2cc7 	:	o_val <= 16'b0111001000000100;
            14'h2cc8 	:	o_val <= 16'b0111001000000110;
            14'h2cc9 	:	o_val <= 16'b0111001000000111;
            14'h2cca 	:	o_val <= 16'b0111001000001001;
            14'h2ccb 	:	o_val <= 16'b0111001000001010;
            14'h2ccc 	:	o_val <= 16'b0111001000001100;
            14'h2ccd 	:	o_val <= 16'b0111001000001101;
            14'h2cce 	:	o_val <= 16'b0111001000001110;
            14'h2ccf 	:	o_val <= 16'b0111001000010000;
            14'h2cd0 	:	o_val <= 16'b0111001000010001;
            14'h2cd1 	:	o_val <= 16'b0111001000010011;
            14'h2cd2 	:	o_val <= 16'b0111001000010100;
            14'h2cd3 	:	o_val <= 16'b0111001000010110;
            14'h2cd4 	:	o_val <= 16'b0111001000010111;
            14'h2cd5 	:	o_val <= 16'b0111001000011000;
            14'h2cd6 	:	o_val <= 16'b0111001000011010;
            14'h2cd7 	:	o_val <= 16'b0111001000011011;
            14'h2cd8 	:	o_val <= 16'b0111001000011101;
            14'h2cd9 	:	o_val <= 16'b0111001000011110;
            14'h2cda 	:	o_val <= 16'b0111001000100000;
            14'h2cdb 	:	o_val <= 16'b0111001000100001;
            14'h2cdc 	:	o_val <= 16'b0111001000100010;
            14'h2cdd 	:	o_val <= 16'b0111001000100100;
            14'h2cde 	:	o_val <= 16'b0111001000100101;
            14'h2cdf 	:	o_val <= 16'b0111001000100111;
            14'h2ce0 	:	o_val <= 16'b0111001000101000;
            14'h2ce1 	:	o_val <= 16'b0111001000101001;
            14'h2ce2 	:	o_val <= 16'b0111001000101011;
            14'h2ce3 	:	o_val <= 16'b0111001000101100;
            14'h2ce4 	:	o_val <= 16'b0111001000101110;
            14'h2ce5 	:	o_val <= 16'b0111001000101111;
            14'h2ce6 	:	o_val <= 16'b0111001000110001;
            14'h2ce7 	:	o_val <= 16'b0111001000110010;
            14'h2ce8 	:	o_val <= 16'b0111001000110011;
            14'h2ce9 	:	o_val <= 16'b0111001000110101;
            14'h2cea 	:	o_val <= 16'b0111001000110110;
            14'h2ceb 	:	o_val <= 16'b0111001000111000;
            14'h2cec 	:	o_val <= 16'b0111001000111001;
            14'h2ced 	:	o_val <= 16'b0111001000111010;
            14'h2cee 	:	o_val <= 16'b0111001000111100;
            14'h2cef 	:	o_val <= 16'b0111001000111101;
            14'h2cf0 	:	o_val <= 16'b0111001000111111;
            14'h2cf1 	:	o_val <= 16'b0111001001000000;
            14'h2cf2 	:	o_val <= 16'b0111001001000010;
            14'h2cf3 	:	o_val <= 16'b0111001001000011;
            14'h2cf4 	:	o_val <= 16'b0111001001000100;
            14'h2cf5 	:	o_val <= 16'b0111001001000110;
            14'h2cf6 	:	o_val <= 16'b0111001001000111;
            14'h2cf7 	:	o_val <= 16'b0111001001001001;
            14'h2cf8 	:	o_val <= 16'b0111001001001010;
            14'h2cf9 	:	o_val <= 16'b0111001001001011;
            14'h2cfa 	:	o_val <= 16'b0111001001001101;
            14'h2cfb 	:	o_val <= 16'b0111001001001110;
            14'h2cfc 	:	o_val <= 16'b0111001001010000;
            14'h2cfd 	:	o_val <= 16'b0111001001010001;
            14'h2cfe 	:	o_val <= 16'b0111001001010011;
            14'h2cff 	:	o_val <= 16'b0111001001010100;
            14'h2d00 	:	o_val <= 16'b0111001001010101;
            14'h2d01 	:	o_val <= 16'b0111001001010111;
            14'h2d02 	:	o_val <= 16'b0111001001011000;
            14'h2d03 	:	o_val <= 16'b0111001001011010;
            14'h2d04 	:	o_val <= 16'b0111001001011011;
            14'h2d05 	:	o_val <= 16'b0111001001011100;
            14'h2d06 	:	o_val <= 16'b0111001001011110;
            14'h2d07 	:	o_val <= 16'b0111001001011111;
            14'h2d08 	:	o_val <= 16'b0111001001100001;
            14'h2d09 	:	o_val <= 16'b0111001001100010;
            14'h2d0a 	:	o_val <= 16'b0111001001100011;
            14'h2d0b 	:	o_val <= 16'b0111001001100101;
            14'h2d0c 	:	o_val <= 16'b0111001001100110;
            14'h2d0d 	:	o_val <= 16'b0111001001101000;
            14'h2d0e 	:	o_val <= 16'b0111001001101001;
            14'h2d0f 	:	o_val <= 16'b0111001001101011;
            14'h2d10 	:	o_val <= 16'b0111001001101100;
            14'h2d11 	:	o_val <= 16'b0111001001101101;
            14'h2d12 	:	o_val <= 16'b0111001001101111;
            14'h2d13 	:	o_val <= 16'b0111001001110000;
            14'h2d14 	:	o_val <= 16'b0111001001110010;
            14'h2d15 	:	o_val <= 16'b0111001001110011;
            14'h2d16 	:	o_val <= 16'b0111001001110100;
            14'h2d17 	:	o_val <= 16'b0111001001110110;
            14'h2d18 	:	o_val <= 16'b0111001001110111;
            14'h2d19 	:	o_val <= 16'b0111001001111001;
            14'h2d1a 	:	o_val <= 16'b0111001001111010;
            14'h2d1b 	:	o_val <= 16'b0111001001111011;
            14'h2d1c 	:	o_val <= 16'b0111001001111101;
            14'h2d1d 	:	o_val <= 16'b0111001001111110;
            14'h2d1e 	:	o_val <= 16'b0111001010000000;
            14'h2d1f 	:	o_val <= 16'b0111001010000001;
            14'h2d20 	:	o_val <= 16'b0111001010000010;
            14'h2d21 	:	o_val <= 16'b0111001010000100;
            14'h2d22 	:	o_val <= 16'b0111001010000101;
            14'h2d23 	:	o_val <= 16'b0111001010000111;
            14'h2d24 	:	o_val <= 16'b0111001010001000;
            14'h2d25 	:	o_val <= 16'b0111001010001001;
            14'h2d26 	:	o_val <= 16'b0111001010001011;
            14'h2d27 	:	o_val <= 16'b0111001010001100;
            14'h2d28 	:	o_val <= 16'b0111001010001110;
            14'h2d29 	:	o_val <= 16'b0111001010001111;
            14'h2d2a 	:	o_val <= 16'b0111001010010000;
            14'h2d2b 	:	o_val <= 16'b0111001010010010;
            14'h2d2c 	:	o_val <= 16'b0111001010010011;
            14'h2d2d 	:	o_val <= 16'b0111001010010101;
            14'h2d2e 	:	o_val <= 16'b0111001010010110;
            14'h2d2f 	:	o_val <= 16'b0111001010010111;
            14'h2d30 	:	o_val <= 16'b0111001010011001;
            14'h2d31 	:	o_val <= 16'b0111001010011010;
            14'h2d32 	:	o_val <= 16'b0111001010011100;
            14'h2d33 	:	o_val <= 16'b0111001010011101;
            14'h2d34 	:	o_val <= 16'b0111001010011110;
            14'h2d35 	:	o_val <= 16'b0111001010100000;
            14'h2d36 	:	o_val <= 16'b0111001010100001;
            14'h2d37 	:	o_val <= 16'b0111001010100011;
            14'h2d38 	:	o_val <= 16'b0111001010100100;
            14'h2d39 	:	o_val <= 16'b0111001010100101;
            14'h2d3a 	:	o_val <= 16'b0111001010100111;
            14'h2d3b 	:	o_val <= 16'b0111001010101000;
            14'h2d3c 	:	o_val <= 16'b0111001010101010;
            14'h2d3d 	:	o_val <= 16'b0111001010101011;
            14'h2d3e 	:	o_val <= 16'b0111001010101100;
            14'h2d3f 	:	o_val <= 16'b0111001010101110;
            14'h2d40 	:	o_val <= 16'b0111001010101111;
            14'h2d41 	:	o_val <= 16'b0111001010110001;
            14'h2d42 	:	o_val <= 16'b0111001010110010;
            14'h2d43 	:	o_val <= 16'b0111001010110011;
            14'h2d44 	:	o_val <= 16'b0111001010110101;
            14'h2d45 	:	o_val <= 16'b0111001010110110;
            14'h2d46 	:	o_val <= 16'b0111001010111000;
            14'h2d47 	:	o_val <= 16'b0111001010111001;
            14'h2d48 	:	o_val <= 16'b0111001010111010;
            14'h2d49 	:	o_val <= 16'b0111001010111100;
            14'h2d4a 	:	o_val <= 16'b0111001010111101;
            14'h2d4b 	:	o_val <= 16'b0111001010111111;
            14'h2d4c 	:	o_val <= 16'b0111001011000000;
            14'h2d4d 	:	o_val <= 16'b0111001011000001;
            14'h2d4e 	:	o_val <= 16'b0111001011000011;
            14'h2d4f 	:	o_val <= 16'b0111001011000100;
            14'h2d50 	:	o_val <= 16'b0111001011000110;
            14'h2d51 	:	o_val <= 16'b0111001011000111;
            14'h2d52 	:	o_val <= 16'b0111001011001000;
            14'h2d53 	:	o_val <= 16'b0111001011001010;
            14'h2d54 	:	o_val <= 16'b0111001011001011;
            14'h2d55 	:	o_val <= 16'b0111001011001100;
            14'h2d56 	:	o_val <= 16'b0111001011001110;
            14'h2d57 	:	o_val <= 16'b0111001011001111;
            14'h2d58 	:	o_val <= 16'b0111001011010001;
            14'h2d59 	:	o_val <= 16'b0111001011010010;
            14'h2d5a 	:	o_val <= 16'b0111001011010011;
            14'h2d5b 	:	o_val <= 16'b0111001011010101;
            14'h2d5c 	:	o_val <= 16'b0111001011010110;
            14'h2d5d 	:	o_val <= 16'b0111001011011000;
            14'h2d5e 	:	o_val <= 16'b0111001011011001;
            14'h2d5f 	:	o_val <= 16'b0111001011011010;
            14'h2d60 	:	o_val <= 16'b0111001011011100;
            14'h2d61 	:	o_val <= 16'b0111001011011101;
            14'h2d62 	:	o_val <= 16'b0111001011011110;
            14'h2d63 	:	o_val <= 16'b0111001011100000;
            14'h2d64 	:	o_val <= 16'b0111001011100001;
            14'h2d65 	:	o_val <= 16'b0111001011100011;
            14'h2d66 	:	o_val <= 16'b0111001011100100;
            14'h2d67 	:	o_val <= 16'b0111001011100101;
            14'h2d68 	:	o_val <= 16'b0111001011100111;
            14'h2d69 	:	o_val <= 16'b0111001011101000;
            14'h2d6a 	:	o_val <= 16'b0111001011101010;
            14'h2d6b 	:	o_val <= 16'b0111001011101011;
            14'h2d6c 	:	o_val <= 16'b0111001011101100;
            14'h2d6d 	:	o_val <= 16'b0111001011101110;
            14'h2d6e 	:	o_val <= 16'b0111001011101111;
            14'h2d6f 	:	o_val <= 16'b0111001011110000;
            14'h2d70 	:	o_val <= 16'b0111001011110010;
            14'h2d71 	:	o_val <= 16'b0111001011110011;
            14'h2d72 	:	o_val <= 16'b0111001011110101;
            14'h2d73 	:	o_val <= 16'b0111001011110110;
            14'h2d74 	:	o_val <= 16'b0111001011110111;
            14'h2d75 	:	o_val <= 16'b0111001011111001;
            14'h2d76 	:	o_val <= 16'b0111001011111010;
            14'h2d77 	:	o_val <= 16'b0111001011111100;
            14'h2d78 	:	o_val <= 16'b0111001011111101;
            14'h2d79 	:	o_val <= 16'b0111001011111110;
            14'h2d7a 	:	o_val <= 16'b0111001100000000;
            14'h2d7b 	:	o_val <= 16'b0111001100000001;
            14'h2d7c 	:	o_val <= 16'b0111001100000010;
            14'h2d7d 	:	o_val <= 16'b0111001100000100;
            14'h2d7e 	:	o_val <= 16'b0111001100000101;
            14'h2d7f 	:	o_val <= 16'b0111001100000111;
            14'h2d80 	:	o_val <= 16'b0111001100001000;
            14'h2d81 	:	o_val <= 16'b0111001100001001;
            14'h2d82 	:	o_val <= 16'b0111001100001011;
            14'h2d83 	:	o_val <= 16'b0111001100001100;
            14'h2d84 	:	o_val <= 16'b0111001100001101;
            14'h2d85 	:	o_val <= 16'b0111001100001111;
            14'h2d86 	:	o_val <= 16'b0111001100010000;
            14'h2d87 	:	o_val <= 16'b0111001100010010;
            14'h2d88 	:	o_val <= 16'b0111001100010011;
            14'h2d89 	:	o_val <= 16'b0111001100010100;
            14'h2d8a 	:	o_val <= 16'b0111001100010110;
            14'h2d8b 	:	o_val <= 16'b0111001100010111;
            14'h2d8c 	:	o_val <= 16'b0111001100011000;
            14'h2d8d 	:	o_val <= 16'b0111001100011010;
            14'h2d8e 	:	o_val <= 16'b0111001100011011;
            14'h2d8f 	:	o_val <= 16'b0111001100011101;
            14'h2d90 	:	o_val <= 16'b0111001100011110;
            14'h2d91 	:	o_val <= 16'b0111001100011111;
            14'h2d92 	:	o_val <= 16'b0111001100100001;
            14'h2d93 	:	o_val <= 16'b0111001100100010;
            14'h2d94 	:	o_val <= 16'b0111001100100011;
            14'h2d95 	:	o_val <= 16'b0111001100100101;
            14'h2d96 	:	o_val <= 16'b0111001100100110;
            14'h2d97 	:	o_val <= 16'b0111001100101000;
            14'h2d98 	:	o_val <= 16'b0111001100101001;
            14'h2d99 	:	o_val <= 16'b0111001100101010;
            14'h2d9a 	:	o_val <= 16'b0111001100101100;
            14'h2d9b 	:	o_val <= 16'b0111001100101101;
            14'h2d9c 	:	o_val <= 16'b0111001100101110;
            14'h2d9d 	:	o_val <= 16'b0111001100110000;
            14'h2d9e 	:	o_val <= 16'b0111001100110001;
            14'h2d9f 	:	o_val <= 16'b0111001100110011;
            14'h2da0 	:	o_val <= 16'b0111001100110100;
            14'h2da1 	:	o_val <= 16'b0111001100110101;
            14'h2da2 	:	o_val <= 16'b0111001100110111;
            14'h2da3 	:	o_val <= 16'b0111001100111000;
            14'h2da4 	:	o_val <= 16'b0111001100111001;
            14'h2da5 	:	o_val <= 16'b0111001100111011;
            14'h2da6 	:	o_val <= 16'b0111001100111100;
            14'h2da7 	:	o_val <= 16'b0111001100111101;
            14'h2da8 	:	o_val <= 16'b0111001100111111;
            14'h2da9 	:	o_val <= 16'b0111001101000000;
            14'h2daa 	:	o_val <= 16'b0111001101000010;
            14'h2dab 	:	o_val <= 16'b0111001101000011;
            14'h2dac 	:	o_val <= 16'b0111001101000100;
            14'h2dad 	:	o_val <= 16'b0111001101000110;
            14'h2dae 	:	o_val <= 16'b0111001101000111;
            14'h2daf 	:	o_val <= 16'b0111001101001000;
            14'h2db0 	:	o_val <= 16'b0111001101001010;
            14'h2db1 	:	o_val <= 16'b0111001101001011;
            14'h2db2 	:	o_val <= 16'b0111001101001101;
            14'h2db3 	:	o_val <= 16'b0111001101001110;
            14'h2db4 	:	o_val <= 16'b0111001101001111;
            14'h2db5 	:	o_val <= 16'b0111001101010001;
            14'h2db6 	:	o_val <= 16'b0111001101010010;
            14'h2db7 	:	o_val <= 16'b0111001101010011;
            14'h2db8 	:	o_val <= 16'b0111001101010101;
            14'h2db9 	:	o_val <= 16'b0111001101010110;
            14'h2dba 	:	o_val <= 16'b0111001101010111;
            14'h2dbb 	:	o_val <= 16'b0111001101011001;
            14'h2dbc 	:	o_val <= 16'b0111001101011010;
            14'h2dbd 	:	o_val <= 16'b0111001101011011;
            14'h2dbe 	:	o_val <= 16'b0111001101011101;
            14'h2dbf 	:	o_val <= 16'b0111001101011110;
            14'h2dc0 	:	o_val <= 16'b0111001101100000;
            14'h2dc1 	:	o_val <= 16'b0111001101100001;
            14'h2dc2 	:	o_val <= 16'b0111001101100010;
            14'h2dc3 	:	o_val <= 16'b0111001101100100;
            14'h2dc4 	:	o_val <= 16'b0111001101100101;
            14'h2dc5 	:	o_val <= 16'b0111001101100110;
            14'h2dc6 	:	o_val <= 16'b0111001101101000;
            14'h2dc7 	:	o_val <= 16'b0111001101101001;
            14'h2dc8 	:	o_val <= 16'b0111001101101010;
            14'h2dc9 	:	o_val <= 16'b0111001101101100;
            14'h2dca 	:	o_val <= 16'b0111001101101101;
            14'h2dcb 	:	o_val <= 16'b0111001101101111;
            14'h2dcc 	:	o_val <= 16'b0111001101110000;
            14'h2dcd 	:	o_val <= 16'b0111001101110001;
            14'h2dce 	:	o_val <= 16'b0111001101110011;
            14'h2dcf 	:	o_val <= 16'b0111001101110100;
            14'h2dd0 	:	o_val <= 16'b0111001101110101;
            14'h2dd1 	:	o_val <= 16'b0111001101110111;
            14'h2dd2 	:	o_val <= 16'b0111001101111000;
            14'h2dd3 	:	o_val <= 16'b0111001101111001;
            14'h2dd4 	:	o_val <= 16'b0111001101111011;
            14'h2dd5 	:	o_val <= 16'b0111001101111100;
            14'h2dd6 	:	o_val <= 16'b0111001101111101;
            14'h2dd7 	:	o_val <= 16'b0111001101111111;
            14'h2dd8 	:	o_val <= 16'b0111001110000000;
            14'h2dd9 	:	o_val <= 16'b0111001110000010;
            14'h2dda 	:	o_val <= 16'b0111001110000011;
            14'h2ddb 	:	o_val <= 16'b0111001110000100;
            14'h2ddc 	:	o_val <= 16'b0111001110000110;
            14'h2ddd 	:	o_val <= 16'b0111001110000111;
            14'h2dde 	:	o_val <= 16'b0111001110001000;
            14'h2ddf 	:	o_val <= 16'b0111001110001010;
            14'h2de0 	:	o_val <= 16'b0111001110001011;
            14'h2de1 	:	o_val <= 16'b0111001110001100;
            14'h2de2 	:	o_val <= 16'b0111001110001110;
            14'h2de3 	:	o_val <= 16'b0111001110001111;
            14'h2de4 	:	o_val <= 16'b0111001110010000;
            14'h2de5 	:	o_val <= 16'b0111001110010010;
            14'h2de6 	:	o_val <= 16'b0111001110010011;
            14'h2de7 	:	o_val <= 16'b0111001110010100;
            14'h2de8 	:	o_val <= 16'b0111001110010110;
            14'h2de9 	:	o_val <= 16'b0111001110010111;
            14'h2dea 	:	o_val <= 16'b0111001110011000;
            14'h2deb 	:	o_val <= 16'b0111001110011010;
            14'h2dec 	:	o_val <= 16'b0111001110011011;
            14'h2ded 	:	o_val <= 16'b0111001110011101;
            14'h2dee 	:	o_val <= 16'b0111001110011110;
            14'h2def 	:	o_val <= 16'b0111001110011111;
            14'h2df0 	:	o_val <= 16'b0111001110100001;
            14'h2df1 	:	o_val <= 16'b0111001110100010;
            14'h2df2 	:	o_val <= 16'b0111001110100011;
            14'h2df3 	:	o_val <= 16'b0111001110100101;
            14'h2df4 	:	o_val <= 16'b0111001110100110;
            14'h2df5 	:	o_val <= 16'b0111001110100111;
            14'h2df6 	:	o_val <= 16'b0111001110101001;
            14'h2df7 	:	o_val <= 16'b0111001110101010;
            14'h2df8 	:	o_val <= 16'b0111001110101011;
            14'h2df9 	:	o_val <= 16'b0111001110101101;
            14'h2dfa 	:	o_val <= 16'b0111001110101110;
            14'h2dfb 	:	o_val <= 16'b0111001110101111;
            14'h2dfc 	:	o_val <= 16'b0111001110110001;
            14'h2dfd 	:	o_val <= 16'b0111001110110010;
            14'h2dfe 	:	o_val <= 16'b0111001110110011;
            14'h2dff 	:	o_val <= 16'b0111001110110101;
            14'h2e00 	:	o_val <= 16'b0111001110110110;
            14'h2e01 	:	o_val <= 16'b0111001110110111;
            14'h2e02 	:	o_val <= 16'b0111001110111001;
            14'h2e03 	:	o_val <= 16'b0111001110111010;
            14'h2e04 	:	o_val <= 16'b0111001110111011;
            14'h2e05 	:	o_val <= 16'b0111001110111101;
            14'h2e06 	:	o_val <= 16'b0111001110111110;
            14'h2e07 	:	o_val <= 16'b0111001110111111;
            14'h2e08 	:	o_val <= 16'b0111001111000001;
            14'h2e09 	:	o_val <= 16'b0111001111000010;
            14'h2e0a 	:	o_val <= 16'b0111001111000100;
            14'h2e0b 	:	o_val <= 16'b0111001111000101;
            14'h2e0c 	:	o_val <= 16'b0111001111000110;
            14'h2e0d 	:	o_val <= 16'b0111001111001000;
            14'h2e0e 	:	o_val <= 16'b0111001111001001;
            14'h2e0f 	:	o_val <= 16'b0111001111001010;
            14'h2e10 	:	o_val <= 16'b0111001111001100;
            14'h2e11 	:	o_val <= 16'b0111001111001101;
            14'h2e12 	:	o_val <= 16'b0111001111001110;
            14'h2e13 	:	o_val <= 16'b0111001111010000;
            14'h2e14 	:	o_val <= 16'b0111001111010001;
            14'h2e15 	:	o_val <= 16'b0111001111010010;
            14'h2e16 	:	o_val <= 16'b0111001111010100;
            14'h2e17 	:	o_val <= 16'b0111001111010101;
            14'h2e18 	:	o_val <= 16'b0111001111010110;
            14'h2e19 	:	o_val <= 16'b0111001111011000;
            14'h2e1a 	:	o_val <= 16'b0111001111011001;
            14'h2e1b 	:	o_val <= 16'b0111001111011010;
            14'h2e1c 	:	o_val <= 16'b0111001111011100;
            14'h2e1d 	:	o_val <= 16'b0111001111011101;
            14'h2e1e 	:	o_val <= 16'b0111001111011110;
            14'h2e1f 	:	o_val <= 16'b0111001111100000;
            14'h2e20 	:	o_val <= 16'b0111001111100001;
            14'h2e21 	:	o_val <= 16'b0111001111100010;
            14'h2e22 	:	o_val <= 16'b0111001111100100;
            14'h2e23 	:	o_val <= 16'b0111001111100101;
            14'h2e24 	:	o_val <= 16'b0111001111100110;
            14'h2e25 	:	o_val <= 16'b0111001111101000;
            14'h2e26 	:	o_val <= 16'b0111001111101001;
            14'h2e27 	:	o_val <= 16'b0111001111101010;
            14'h2e28 	:	o_val <= 16'b0111001111101100;
            14'h2e29 	:	o_val <= 16'b0111001111101101;
            14'h2e2a 	:	o_val <= 16'b0111001111101110;
            14'h2e2b 	:	o_val <= 16'b0111001111110000;
            14'h2e2c 	:	o_val <= 16'b0111001111110001;
            14'h2e2d 	:	o_val <= 16'b0111001111110010;
            14'h2e2e 	:	o_val <= 16'b0111001111110100;
            14'h2e2f 	:	o_val <= 16'b0111001111110101;
            14'h2e30 	:	o_val <= 16'b0111001111110110;
            14'h2e31 	:	o_val <= 16'b0111001111111000;
            14'h2e32 	:	o_val <= 16'b0111001111111001;
            14'h2e33 	:	o_val <= 16'b0111001111111010;
            14'h2e34 	:	o_val <= 16'b0111001111111100;
            14'h2e35 	:	o_val <= 16'b0111001111111101;
            14'h2e36 	:	o_val <= 16'b0111001111111110;
            14'h2e37 	:	o_val <= 16'b0111010000000000;
            14'h2e38 	:	o_val <= 16'b0111010000000001;
            14'h2e39 	:	o_val <= 16'b0111010000000010;
            14'h2e3a 	:	o_val <= 16'b0111010000000100;
            14'h2e3b 	:	o_val <= 16'b0111010000000101;
            14'h2e3c 	:	o_val <= 16'b0111010000000110;
            14'h2e3d 	:	o_val <= 16'b0111010000001000;
            14'h2e3e 	:	o_val <= 16'b0111010000001001;
            14'h2e3f 	:	o_val <= 16'b0111010000001010;
            14'h2e40 	:	o_val <= 16'b0111010000001011;
            14'h2e41 	:	o_val <= 16'b0111010000001101;
            14'h2e42 	:	o_val <= 16'b0111010000001110;
            14'h2e43 	:	o_val <= 16'b0111010000001111;
            14'h2e44 	:	o_val <= 16'b0111010000010001;
            14'h2e45 	:	o_val <= 16'b0111010000010010;
            14'h2e46 	:	o_val <= 16'b0111010000010011;
            14'h2e47 	:	o_val <= 16'b0111010000010101;
            14'h2e48 	:	o_val <= 16'b0111010000010110;
            14'h2e49 	:	o_val <= 16'b0111010000010111;
            14'h2e4a 	:	o_val <= 16'b0111010000011001;
            14'h2e4b 	:	o_val <= 16'b0111010000011010;
            14'h2e4c 	:	o_val <= 16'b0111010000011011;
            14'h2e4d 	:	o_val <= 16'b0111010000011101;
            14'h2e4e 	:	o_val <= 16'b0111010000011110;
            14'h2e4f 	:	o_val <= 16'b0111010000011111;
            14'h2e50 	:	o_val <= 16'b0111010000100001;
            14'h2e51 	:	o_val <= 16'b0111010000100010;
            14'h2e52 	:	o_val <= 16'b0111010000100011;
            14'h2e53 	:	o_val <= 16'b0111010000100101;
            14'h2e54 	:	o_val <= 16'b0111010000100110;
            14'h2e55 	:	o_val <= 16'b0111010000100111;
            14'h2e56 	:	o_val <= 16'b0111010000101001;
            14'h2e57 	:	o_val <= 16'b0111010000101010;
            14'h2e58 	:	o_val <= 16'b0111010000101011;
            14'h2e59 	:	o_val <= 16'b0111010000101101;
            14'h2e5a 	:	o_val <= 16'b0111010000101110;
            14'h2e5b 	:	o_val <= 16'b0111010000101111;
            14'h2e5c 	:	o_val <= 16'b0111010000110001;
            14'h2e5d 	:	o_val <= 16'b0111010000110010;
            14'h2e5e 	:	o_val <= 16'b0111010000110011;
            14'h2e5f 	:	o_val <= 16'b0111010000110100;
            14'h2e60 	:	o_val <= 16'b0111010000110110;
            14'h2e61 	:	o_val <= 16'b0111010000110111;
            14'h2e62 	:	o_val <= 16'b0111010000111000;
            14'h2e63 	:	o_val <= 16'b0111010000111010;
            14'h2e64 	:	o_val <= 16'b0111010000111011;
            14'h2e65 	:	o_val <= 16'b0111010000111100;
            14'h2e66 	:	o_val <= 16'b0111010000111110;
            14'h2e67 	:	o_val <= 16'b0111010000111111;
            14'h2e68 	:	o_val <= 16'b0111010001000000;
            14'h2e69 	:	o_val <= 16'b0111010001000010;
            14'h2e6a 	:	o_val <= 16'b0111010001000011;
            14'h2e6b 	:	o_val <= 16'b0111010001000100;
            14'h2e6c 	:	o_val <= 16'b0111010001000110;
            14'h2e6d 	:	o_val <= 16'b0111010001000111;
            14'h2e6e 	:	o_val <= 16'b0111010001001000;
            14'h2e6f 	:	o_val <= 16'b0111010001001001;
            14'h2e70 	:	o_val <= 16'b0111010001001011;
            14'h2e71 	:	o_val <= 16'b0111010001001100;
            14'h2e72 	:	o_val <= 16'b0111010001001101;
            14'h2e73 	:	o_val <= 16'b0111010001001111;
            14'h2e74 	:	o_val <= 16'b0111010001010000;
            14'h2e75 	:	o_val <= 16'b0111010001010001;
            14'h2e76 	:	o_val <= 16'b0111010001010011;
            14'h2e77 	:	o_val <= 16'b0111010001010100;
            14'h2e78 	:	o_val <= 16'b0111010001010101;
            14'h2e79 	:	o_val <= 16'b0111010001010111;
            14'h2e7a 	:	o_val <= 16'b0111010001011000;
            14'h2e7b 	:	o_val <= 16'b0111010001011001;
            14'h2e7c 	:	o_val <= 16'b0111010001011011;
            14'h2e7d 	:	o_val <= 16'b0111010001011100;
            14'h2e7e 	:	o_val <= 16'b0111010001011101;
            14'h2e7f 	:	o_val <= 16'b0111010001011110;
            14'h2e80 	:	o_val <= 16'b0111010001100000;
            14'h2e81 	:	o_val <= 16'b0111010001100001;
            14'h2e82 	:	o_val <= 16'b0111010001100010;
            14'h2e83 	:	o_val <= 16'b0111010001100100;
            14'h2e84 	:	o_val <= 16'b0111010001100101;
            14'h2e85 	:	o_val <= 16'b0111010001100110;
            14'h2e86 	:	o_val <= 16'b0111010001101000;
            14'h2e87 	:	o_val <= 16'b0111010001101001;
            14'h2e88 	:	o_val <= 16'b0111010001101010;
            14'h2e89 	:	o_val <= 16'b0111010001101100;
            14'h2e8a 	:	o_val <= 16'b0111010001101101;
            14'h2e8b 	:	o_val <= 16'b0111010001101110;
            14'h2e8c 	:	o_val <= 16'b0111010001101111;
            14'h2e8d 	:	o_val <= 16'b0111010001110001;
            14'h2e8e 	:	o_val <= 16'b0111010001110010;
            14'h2e8f 	:	o_val <= 16'b0111010001110011;
            14'h2e90 	:	o_val <= 16'b0111010001110101;
            14'h2e91 	:	o_val <= 16'b0111010001110110;
            14'h2e92 	:	o_val <= 16'b0111010001110111;
            14'h2e93 	:	o_val <= 16'b0111010001111001;
            14'h2e94 	:	o_val <= 16'b0111010001111010;
            14'h2e95 	:	o_val <= 16'b0111010001111011;
            14'h2e96 	:	o_val <= 16'b0111010001111100;
            14'h2e97 	:	o_val <= 16'b0111010001111110;
            14'h2e98 	:	o_val <= 16'b0111010001111111;
            14'h2e99 	:	o_val <= 16'b0111010010000000;
            14'h2e9a 	:	o_val <= 16'b0111010010000010;
            14'h2e9b 	:	o_val <= 16'b0111010010000011;
            14'h2e9c 	:	o_val <= 16'b0111010010000100;
            14'h2e9d 	:	o_val <= 16'b0111010010000110;
            14'h2e9e 	:	o_val <= 16'b0111010010000111;
            14'h2e9f 	:	o_val <= 16'b0111010010001000;
            14'h2ea0 	:	o_val <= 16'b0111010010001001;
            14'h2ea1 	:	o_val <= 16'b0111010010001011;
            14'h2ea2 	:	o_val <= 16'b0111010010001100;
            14'h2ea3 	:	o_val <= 16'b0111010010001101;
            14'h2ea4 	:	o_val <= 16'b0111010010001111;
            14'h2ea5 	:	o_val <= 16'b0111010010010000;
            14'h2ea6 	:	o_val <= 16'b0111010010010001;
            14'h2ea7 	:	o_val <= 16'b0111010010010011;
            14'h2ea8 	:	o_val <= 16'b0111010010010100;
            14'h2ea9 	:	o_val <= 16'b0111010010010101;
            14'h2eaa 	:	o_val <= 16'b0111010010010110;
            14'h2eab 	:	o_val <= 16'b0111010010011000;
            14'h2eac 	:	o_val <= 16'b0111010010011001;
            14'h2ead 	:	o_val <= 16'b0111010010011010;
            14'h2eae 	:	o_val <= 16'b0111010010011100;
            14'h2eaf 	:	o_val <= 16'b0111010010011101;
            14'h2eb0 	:	o_val <= 16'b0111010010011110;
            14'h2eb1 	:	o_val <= 16'b0111010010100000;
            14'h2eb2 	:	o_val <= 16'b0111010010100001;
            14'h2eb3 	:	o_val <= 16'b0111010010100010;
            14'h2eb4 	:	o_val <= 16'b0111010010100011;
            14'h2eb5 	:	o_val <= 16'b0111010010100101;
            14'h2eb6 	:	o_val <= 16'b0111010010100110;
            14'h2eb7 	:	o_val <= 16'b0111010010100111;
            14'h2eb8 	:	o_val <= 16'b0111010010101001;
            14'h2eb9 	:	o_val <= 16'b0111010010101010;
            14'h2eba 	:	o_val <= 16'b0111010010101011;
            14'h2ebb 	:	o_val <= 16'b0111010010101100;
            14'h2ebc 	:	o_val <= 16'b0111010010101110;
            14'h2ebd 	:	o_val <= 16'b0111010010101111;
            14'h2ebe 	:	o_val <= 16'b0111010010110000;
            14'h2ebf 	:	o_val <= 16'b0111010010110010;
            14'h2ec0 	:	o_val <= 16'b0111010010110011;
            14'h2ec1 	:	o_val <= 16'b0111010010110100;
            14'h2ec2 	:	o_val <= 16'b0111010010110110;
            14'h2ec3 	:	o_val <= 16'b0111010010110111;
            14'h2ec4 	:	o_val <= 16'b0111010010111000;
            14'h2ec5 	:	o_val <= 16'b0111010010111001;
            14'h2ec6 	:	o_val <= 16'b0111010010111011;
            14'h2ec7 	:	o_val <= 16'b0111010010111100;
            14'h2ec8 	:	o_val <= 16'b0111010010111101;
            14'h2ec9 	:	o_val <= 16'b0111010010111111;
            14'h2eca 	:	o_val <= 16'b0111010011000000;
            14'h2ecb 	:	o_val <= 16'b0111010011000001;
            14'h2ecc 	:	o_val <= 16'b0111010011000010;
            14'h2ecd 	:	o_val <= 16'b0111010011000100;
            14'h2ece 	:	o_val <= 16'b0111010011000101;
            14'h2ecf 	:	o_val <= 16'b0111010011000110;
            14'h2ed0 	:	o_val <= 16'b0111010011001000;
            14'h2ed1 	:	o_val <= 16'b0111010011001001;
            14'h2ed2 	:	o_val <= 16'b0111010011001010;
            14'h2ed3 	:	o_val <= 16'b0111010011001011;
            14'h2ed4 	:	o_val <= 16'b0111010011001101;
            14'h2ed5 	:	o_val <= 16'b0111010011001110;
            14'h2ed6 	:	o_val <= 16'b0111010011001111;
            14'h2ed7 	:	o_val <= 16'b0111010011010001;
            14'h2ed8 	:	o_val <= 16'b0111010011010010;
            14'h2ed9 	:	o_val <= 16'b0111010011010011;
            14'h2eda 	:	o_val <= 16'b0111010011010100;
            14'h2edb 	:	o_val <= 16'b0111010011010110;
            14'h2edc 	:	o_val <= 16'b0111010011010111;
            14'h2edd 	:	o_val <= 16'b0111010011011000;
            14'h2ede 	:	o_val <= 16'b0111010011011010;
            14'h2edf 	:	o_val <= 16'b0111010011011011;
            14'h2ee0 	:	o_val <= 16'b0111010011011100;
            14'h2ee1 	:	o_val <= 16'b0111010011011101;
            14'h2ee2 	:	o_val <= 16'b0111010011011111;
            14'h2ee3 	:	o_val <= 16'b0111010011100000;
            14'h2ee4 	:	o_val <= 16'b0111010011100001;
            14'h2ee5 	:	o_val <= 16'b0111010011100010;
            14'h2ee6 	:	o_val <= 16'b0111010011100100;
            14'h2ee7 	:	o_val <= 16'b0111010011100101;
            14'h2ee8 	:	o_val <= 16'b0111010011100110;
            14'h2ee9 	:	o_val <= 16'b0111010011101000;
            14'h2eea 	:	o_val <= 16'b0111010011101001;
            14'h2eeb 	:	o_val <= 16'b0111010011101010;
            14'h2eec 	:	o_val <= 16'b0111010011101011;
            14'h2eed 	:	o_val <= 16'b0111010011101101;
            14'h2eee 	:	o_val <= 16'b0111010011101110;
            14'h2eef 	:	o_val <= 16'b0111010011101111;
            14'h2ef0 	:	o_val <= 16'b0111010011110001;
            14'h2ef1 	:	o_val <= 16'b0111010011110010;
            14'h2ef2 	:	o_val <= 16'b0111010011110011;
            14'h2ef3 	:	o_val <= 16'b0111010011110100;
            14'h2ef4 	:	o_val <= 16'b0111010011110110;
            14'h2ef5 	:	o_val <= 16'b0111010011110111;
            14'h2ef6 	:	o_val <= 16'b0111010011111000;
            14'h2ef7 	:	o_val <= 16'b0111010011111001;
            14'h2ef8 	:	o_val <= 16'b0111010011111011;
            14'h2ef9 	:	o_val <= 16'b0111010011111100;
            14'h2efa 	:	o_val <= 16'b0111010011111101;
            14'h2efb 	:	o_val <= 16'b0111010011111111;
            14'h2efc 	:	o_val <= 16'b0111010100000000;
            14'h2efd 	:	o_val <= 16'b0111010100000001;
            14'h2efe 	:	o_val <= 16'b0111010100000010;
            14'h2eff 	:	o_val <= 16'b0111010100000100;
            14'h2f00 	:	o_val <= 16'b0111010100000101;
            14'h2f01 	:	o_val <= 16'b0111010100000110;
            14'h2f02 	:	o_val <= 16'b0111010100001000;
            14'h2f03 	:	o_val <= 16'b0111010100001001;
            14'h2f04 	:	o_val <= 16'b0111010100001010;
            14'h2f05 	:	o_val <= 16'b0111010100001011;
            14'h2f06 	:	o_val <= 16'b0111010100001101;
            14'h2f07 	:	o_val <= 16'b0111010100001110;
            14'h2f08 	:	o_val <= 16'b0111010100001111;
            14'h2f09 	:	o_val <= 16'b0111010100010000;
            14'h2f0a 	:	o_val <= 16'b0111010100010010;
            14'h2f0b 	:	o_val <= 16'b0111010100010011;
            14'h2f0c 	:	o_val <= 16'b0111010100010100;
            14'h2f0d 	:	o_val <= 16'b0111010100010101;
            14'h2f0e 	:	o_val <= 16'b0111010100010111;
            14'h2f0f 	:	o_val <= 16'b0111010100011000;
            14'h2f10 	:	o_val <= 16'b0111010100011001;
            14'h2f11 	:	o_val <= 16'b0111010100011011;
            14'h2f12 	:	o_val <= 16'b0111010100011100;
            14'h2f13 	:	o_val <= 16'b0111010100011101;
            14'h2f14 	:	o_val <= 16'b0111010100011110;
            14'h2f15 	:	o_val <= 16'b0111010100100000;
            14'h2f16 	:	o_val <= 16'b0111010100100001;
            14'h2f17 	:	o_val <= 16'b0111010100100010;
            14'h2f18 	:	o_val <= 16'b0111010100100011;
            14'h2f19 	:	o_val <= 16'b0111010100100101;
            14'h2f1a 	:	o_val <= 16'b0111010100100110;
            14'h2f1b 	:	o_val <= 16'b0111010100100111;
            14'h2f1c 	:	o_val <= 16'b0111010100101000;
            14'h2f1d 	:	o_val <= 16'b0111010100101010;
            14'h2f1e 	:	o_val <= 16'b0111010100101011;
            14'h2f1f 	:	o_val <= 16'b0111010100101100;
            14'h2f20 	:	o_val <= 16'b0111010100101110;
            14'h2f21 	:	o_val <= 16'b0111010100101111;
            14'h2f22 	:	o_val <= 16'b0111010100110000;
            14'h2f23 	:	o_val <= 16'b0111010100110001;
            14'h2f24 	:	o_val <= 16'b0111010100110011;
            14'h2f25 	:	o_val <= 16'b0111010100110100;
            14'h2f26 	:	o_val <= 16'b0111010100110101;
            14'h2f27 	:	o_val <= 16'b0111010100110110;
            14'h2f28 	:	o_val <= 16'b0111010100111000;
            14'h2f29 	:	o_val <= 16'b0111010100111001;
            14'h2f2a 	:	o_val <= 16'b0111010100111010;
            14'h2f2b 	:	o_val <= 16'b0111010100111011;
            14'h2f2c 	:	o_val <= 16'b0111010100111101;
            14'h2f2d 	:	o_val <= 16'b0111010100111110;
            14'h2f2e 	:	o_val <= 16'b0111010100111111;
            14'h2f2f 	:	o_val <= 16'b0111010101000000;
            14'h2f30 	:	o_val <= 16'b0111010101000010;
            14'h2f31 	:	o_val <= 16'b0111010101000011;
            14'h2f32 	:	o_val <= 16'b0111010101000100;
            14'h2f33 	:	o_val <= 16'b0111010101000110;
            14'h2f34 	:	o_val <= 16'b0111010101000111;
            14'h2f35 	:	o_val <= 16'b0111010101001000;
            14'h2f36 	:	o_val <= 16'b0111010101001001;
            14'h2f37 	:	o_val <= 16'b0111010101001011;
            14'h2f38 	:	o_val <= 16'b0111010101001100;
            14'h2f39 	:	o_val <= 16'b0111010101001101;
            14'h2f3a 	:	o_val <= 16'b0111010101001110;
            14'h2f3b 	:	o_val <= 16'b0111010101010000;
            14'h2f3c 	:	o_val <= 16'b0111010101010001;
            14'h2f3d 	:	o_val <= 16'b0111010101010010;
            14'h2f3e 	:	o_val <= 16'b0111010101010011;
            14'h2f3f 	:	o_val <= 16'b0111010101010101;
            14'h2f40 	:	o_val <= 16'b0111010101010110;
            14'h2f41 	:	o_val <= 16'b0111010101010111;
            14'h2f42 	:	o_val <= 16'b0111010101011000;
            14'h2f43 	:	o_val <= 16'b0111010101011010;
            14'h2f44 	:	o_val <= 16'b0111010101011011;
            14'h2f45 	:	o_val <= 16'b0111010101011100;
            14'h2f46 	:	o_val <= 16'b0111010101011101;
            14'h2f47 	:	o_val <= 16'b0111010101011111;
            14'h2f48 	:	o_val <= 16'b0111010101100000;
            14'h2f49 	:	o_val <= 16'b0111010101100001;
            14'h2f4a 	:	o_val <= 16'b0111010101100010;
            14'h2f4b 	:	o_val <= 16'b0111010101100100;
            14'h2f4c 	:	o_val <= 16'b0111010101100101;
            14'h2f4d 	:	o_val <= 16'b0111010101100110;
            14'h2f4e 	:	o_val <= 16'b0111010101100111;
            14'h2f4f 	:	o_val <= 16'b0111010101101001;
            14'h2f50 	:	o_val <= 16'b0111010101101010;
            14'h2f51 	:	o_val <= 16'b0111010101101011;
            14'h2f52 	:	o_val <= 16'b0111010101101100;
            14'h2f53 	:	o_val <= 16'b0111010101101110;
            14'h2f54 	:	o_val <= 16'b0111010101101111;
            14'h2f55 	:	o_val <= 16'b0111010101110000;
            14'h2f56 	:	o_val <= 16'b0111010101110001;
            14'h2f57 	:	o_val <= 16'b0111010101110011;
            14'h2f58 	:	o_val <= 16'b0111010101110100;
            14'h2f59 	:	o_val <= 16'b0111010101110101;
            14'h2f5a 	:	o_val <= 16'b0111010101110110;
            14'h2f5b 	:	o_val <= 16'b0111010101111000;
            14'h2f5c 	:	o_val <= 16'b0111010101111001;
            14'h2f5d 	:	o_val <= 16'b0111010101111010;
            14'h2f5e 	:	o_val <= 16'b0111010101111011;
            14'h2f5f 	:	o_val <= 16'b0111010101111101;
            14'h2f60 	:	o_val <= 16'b0111010101111110;
            14'h2f61 	:	o_val <= 16'b0111010101111111;
            14'h2f62 	:	o_val <= 16'b0111010110000000;
            14'h2f63 	:	o_val <= 16'b0111010110000010;
            14'h2f64 	:	o_val <= 16'b0111010110000011;
            14'h2f65 	:	o_val <= 16'b0111010110000100;
            14'h2f66 	:	o_val <= 16'b0111010110000101;
            14'h2f67 	:	o_val <= 16'b0111010110000111;
            14'h2f68 	:	o_val <= 16'b0111010110001000;
            14'h2f69 	:	o_val <= 16'b0111010110001001;
            14'h2f6a 	:	o_val <= 16'b0111010110001010;
            14'h2f6b 	:	o_val <= 16'b0111010110001100;
            14'h2f6c 	:	o_val <= 16'b0111010110001101;
            14'h2f6d 	:	o_val <= 16'b0111010110001110;
            14'h2f6e 	:	o_val <= 16'b0111010110001111;
            14'h2f6f 	:	o_val <= 16'b0111010110010001;
            14'h2f70 	:	o_val <= 16'b0111010110010010;
            14'h2f71 	:	o_val <= 16'b0111010110010011;
            14'h2f72 	:	o_val <= 16'b0111010110010100;
            14'h2f73 	:	o_val <= 16'b0111010110010110;
            14'h2f74 	:	o_val <= 16'b0111010110010111;
            14'h2f75 	:	o_val <= 16'b0111010110011000;
            14'h2f76 	:	o_val <= 16'b0111010110011001;
            14'h2f77 	:	o_val <= 16'b0111010110011010;
            14'h2f78 	:	o_val <= 16'b0111010110011100;
            14'h2f79 	:	o_val <= 16'b0111010110011101;
            14'h2f7a 	:	o_val <= 16'b0111010110011110;
            14'h2f7b 	:	o_val <= 16'b0111010110011111;
            14'h2f7c 	:	o_val <= 16'b0111010110100001;
            14'h2f7d 	:	o_val <= 16'b0111010110100010;
            14'h2f7e 	:	o_val <= 16'b0111010110100011;
            14'h2f7f 	:	o_val <= 16'b0111010110100100;
            14'h2f80 	:	o_val <= 16'b0111010110100110;
            14'h2f81 	:	o_val <= 16'b0111010110100111;
            14'h2f82 	:	o_val <= 16'b0111010110101000;
            14'h2f83 	:	o_val <= 16'b0111010110101001;
            14'h2f84 	:	o_val <= 16'b0111010110101011;
            14'h2f85 	:	o_val <= 16'b0111010110101100;
            14'h2f86 	:	o_val <= 16'b0111010110101101;
            14'h2f87 	:	o_val <= 16'b0111010110101110;
            14'h2f88 	:	o_val <= 16'b0111010110110000;
            14'h2f89 	:	o_val <= 16'b0111010110110001;
            14'h2f8a 	:	o_val <= 16'b0111010110110010;
            14'h2f8b 	:	o_val <= 16'b0111010110110011;
            14'h2f8c 	:	o_val <= 16'b0111010110110100;
            14'h2f8d 	:	o_val <= 16'b0111010110110110;
            14'h2f8e 	:	o_val <= 16'b0111010110110111;
            14'h2f8f 	:	o_val <= 16'b0111010110111000;
            14'h2f90 	:	o_val <= 16'b0111010110111001;
            14'h2f91 	:	o_val <= 16'b0111010110111011;
            14'h2f92 	:	o_val <= 16'b0111010110111100;
            14'h2f93 	:	o_val <= 16'b0111010110111101;
            14'h2f94 	:	o_val <= 16'b0111010110111110;
            14'h2f95 	:	o_val <= 16'b0111010111000000;
            14'h2f96 	:	o_val <= 16'b0111010111000001;
            14'h2f97 	:	o_val <= 16'b0111010111000010;
            14'h2f98 	:	o_val <= 16'b0111010111000011;
            14'h2f99 	:	o_val <= 16'b0111010111000100;
            14'h2f9a 	:	o_val <= 16'b0111010111000110;
            14'h2f9b 	:	o_val <= 16'b0111010111000111;
            14'h2f9c 	:	o_val <= 16'b0111010111001000;
            14'h2f9d 	:	o_val <= 16'b0111010111001001;
            14'h2f9e 	:	o_val <= 16'b0111010111001011;
            14'h2f9f 	:	o_val <= 16'b0111010111001100;
            14'h2fa0 	:	o_val <= 16'b0111010111001101;
            14'h2fa1 	:	o_val <= 16'b0111010111001110;
            14'h2fa2 	:	o_val <= 16'b0111010111010000;
            14'h2fa3 	:	o_val <= 16'b0111010111010001;
            14'h2fa4 	:	o_val <= 16'b0111010111010010;
            14'h2fa5 	:	o_val <= 16'b0111010111010011;
            14'h2fa6 	:	o_val <= 16'b0111010111010100;
            14'h2fa7 	:	o_val <= 16'b0111010111010110;
            14'h2fa8 	:	o_val <= 16'b0111010111010111;
            14'h2fa9 	:	o_val <= 16'b0111010111011000;
            14'h2faa 	:	o_val <= 16'b0111010111011001;
            14'h2fab 	:	o_val <= 16'b0111010111011011;
            14'h2fac 	:	o_val <= 16'b0111010111011100;
            14'h2fad 	:	o_val <= 16'b0111010111011101;
            14'h2fae 	:	o_val <= 16'b0111010111011110;
            14'h2faf 	:	o_val <= 16'b0111010111100000;
            14'h2fb0 	:	o_val <= 16'b0111010111100001;
            14'h2fb1 	:	o_val <= 16'b0111010111100010;
            14'h2fb2 	:	o_val <= 16'b0111010111100011;
            14'h2fb3 	:	o_val <= 16'b0111010111100100;
            14'h2fb4 	:	o_val <= 16'b0111010111100110;
            14'h2fb5 	:	o_val <= 16'b0111010111100111;
            14'h2fb6 	:	o_val <= 16'b0111010111101000;
            14'h2fb7 	:	o_val <= 16'b0111010111101001;
            14'h2fb8 	:	o_val <= 16'b0111010111101011;
            14'h2fb9 	:	o_val <= 16'b0111010111101100;
            14'h2fba 	:	o_val <= 16'b0111010111101101;
            14'h2fbb 	:	o_val <= 16'b0111010111101110;
            14'h2fbc 	:	o_val <= 16'b0111010111101111;
            14'h2fbd 	:	o_val <= 16'b0111010111110001;
            14'h2fbe 	:	o_val <= 16'b0111010111110010;
            14'h2fbf 	:	o_val <= 16'b0111010111110011;
            14'h2fc0 	:	o_val <= 16'b0111010111110100;
            14'h2fc1 	:	o_val <= 16'b0111010111110110;
            14'h2fc2 	:	o_val <= 16'b0111010111110111;
            14'h2fc3 	:	o_val <= 16'b0111010111111000;
            14'h2fc4 	:	o_val <= 16'b0111010111111001;
            14'h2fc5 	:	o_val <= 16'b0111010111111010;
            14'h2fc6 	:	o_val <= 16'b0111010111111100;
            14'h2fc7 	:	o_val <= 16'b0111010111111101;
            14'h2fc8 	:	o_val <= 16'b0111010111111110;
            14'h2fc9 	:	o_val <= 16'b0111010111111111;
            14'h2fca 	:	o_val <= 16'b0111011000000000;
            14'h2fcb 	:	o_val <= 16'b0111011000000010;
            14'h2fcc 	:	o_val <= 16'b0111011000000011;
            14'h2fcd 	:	o_val <= 16'b0111011000000100;
            14'h2fce 	:	o_val <= 16'b0111011000000101;
            14'h2fcf 	:	o_val <= 16'b0111011000000111;
            14'h2fd0 	:	o_val <= 16'b0111011000001000;
            14'h2fd1 	:	o_val <= 16'b0111011000001001;
            14'h2fd2 	:	o_val <= 16'b0111011000001010;
            14'h2fd3 	:	o_val <= 16'b0111011000001011;
            14'h2fd4 	:	o_val <= 16'b0111011000001101;
            14'h2fd5 	:	o_val <= 16'b0111011000001110;
            14'h2fd6 	:	o_val <= 16'b0111011000001111;
            14'h2fd7 	:	o_val <= 16'b0111011000010000;
            14'h2fd8 	:	o_val <= 16'b0111011000010001;
            14'h2fd9 	:	o_val <= 16'b0111011000010011;
            14'h2fda 	:	o_val <= 16'b0111011000010100;
            14'h2fdb 	:	o_val <= 16'b0111011000010101;
            14'h2fdc 	:	o_val <= 16'b0111011000010110;
            14'h2fdd 	:	o_val <= 16'b0111011000011000;
            14'h2fde 	:	o_val <= 16'b0111011000011001;
            14'h2fdf 	:	o_val <= 16'b0111011000011010;
            14'h2fe0 	:	o_val <= 16'b0111011000011011;
            14'h2fe1 	:	o_val <= 16'b0111011000011100;
            14'h2fe2 	:	o_val <= 16'b0111011000011110;
            14'h2fe3 	:	o_val <= 16'b0111011000011111;
            14'h2fe4 	:	o_val <= 16'b0111011000100000;
            14'h2fe5 	:	o_val <= 16'b0111011000100001;
            14'h2fe6 	:	o_val <= 16'b0111011000100010;
            14'h2fe7 	:	o_val <= 16'b0111011000100100;
            14'h2fe8 	:	o_val <= 16'b0111011000100101;
            14'h2fe9 	:	o_val <= 16'b0111011000100110;
            14'h2fea 	:	o_val <= 16'b0111011000100111;
            14'h2feb 	:	o_val <= 16'b0111011000101000;
            14'h2fec 	:	o_val <= 16'b0111011000101010;
            14'h2fed 	:	o_val <= 16'b0111011000101011;
            14'h2fee 	:	o_val <= 16'b0111011000101100;
            14'h2fef 	:	o_val <= 16'b0111011000101101;
            14'h2ff0 	:	o_val <= 16'b0111011000101111;
            14'h2ff1 	:	o_val <= 16'b0111011000110000;
            14'h2ff2 	:	o_val <= 16'b0111011000110001;
            14'h2ff3 	:	o_val <= 16'b0111011000110010;
            14'h2ff4 	:	o_val <= 16'b0111011000110011;
            14'h2ff5 	:	o_val <= 16'b0111011000110101;
            14'h2ff6 	:	o_val <= 16'b0111011000110110;
            14'h2ff7 	:	o_val <= 16'b0111011000110111;
            14'h2ff8 	:	o_val <= 16'b0111011000111000;
            14'h2ff9 	:	o_val <= 16'b0111011000111001;
            14'h2ffa 	:	o_val <= 16'b0111011000111011;
            14'h2ffb 	:	o_val <= 16'b0111011000111100;
            14'h2ffc 	:	o_val <= 16'b0111011000111101;
            14'h2ffd 	:	o_val <= 16'b0111011000111110;
            14'h2ffe 	:	o_val <= 16'b0111011000111111;
            14'h2fff 	:	o_val <= 16'b0111011001000001;
            14'h3000 	:	o_val <= 16'b0111011001000010;
            14'h3001 	:	o_val <= 16'b0111011001000011;
            14'h3002 	:	o_val <= 16'b0111011001000100;
            14'h3003 	:	o_val <= 16'b0111011001000101;
            14'h3004 	:	o_val <= 16'b0111011001000111;
            14'h3005 	:	o_val <= 16'b0111011001001000;
            14'h3006 	:	o_val <= 16'b0111011001001001;
            14'h3007 	:	o_val <= 16'b0111011001001010;
            14'h3008 	:	o_val <= 16'b0111011001001011;
            14'h3009 	:	o_val <= 16'b0111011001001101;
            14'h300a 	:	o_val <= 16'b0111011001001110;
            14'h300b 	:	o_val <= 16'b0111011001001111;
            14'h300c 	:	o_val <= 16'b0111011001010000;
            14'h300d 	:	o_val <= 16'b0111011001010001;
            14'h300e 	:	o_val <= 16'b0111011001010011;
            14'h300f 	:	o_val <= 16'b0111011001010100;
            14'h3010 	:	o_val <= 16'b0111011001010101;
            14'h3011 	:	o_val <= 16'b0111011001010110;
            14'h3012 	:	o_val <= 16'b0111011001010111;
            14'h3013 	:	o_val <= 16'b0111011001011001;
            14'h3014 	:	o_val <= 16'b0111011001011010;
            14'h3015 	:	o_val <= 16'b0111011001011011;
            14'h3016 	:	o_val <= 16'b0111011001011100;
            14'h3017 	:	o_val <= 16'b0111011001011101;
            14'h3018 	:	o_val <= 16'b0111011001011111;
            14'h3019 	:	o_val <= 16'b0111011001100000;
            14'h301a 	:	o_val <= 16'b0111011001100001;
            14'h301b 	:	o_val <= 16'b0111011001100010;
            14'h301c 	:	o_val <= 16'b0111011001100011;
            14'h301d 	:	o_val <= 16'b0111011001100101;
            14'h301e 	:	o_val <= 16'b0111011001100110;
            14'h301f 	:	o_val <= 16'b0111011001100111;
            14'h3020 	:	o_val <= 16'b0111011001101000;
            14'h3021 	:	o_val <= 16'b0111011001101001;
            14'h3022 	:	o_val <= 16'b0111011001101010;
            14'h3023 	:	o_val <= 16'b0111011001101100;
            14'h3024 	:	o_val <= 16'b0111011001101101;
            14'h3025 	:	o_val <= 16'b0111011001101110;
            14'h3026 	:	o_val <= 16'b0111011001101111;
            14'h3027 	:	o_val <= 16'b0111011001110000;
            14'h3028 	:	o_val <= 16'b0111011001110010;
            14'h3029 	:	o_val <= 16'b0111011001110011;
            14'h302a 	:	o_val <= 16'b0111011001110100;
            14'h302b 	:	o_val <= 16'b0111011001110101;
            14'h302c 	:	o_val <= 16'b0111011001110110;
            14'h302d 	:	o_val <= 16'b0111011001111000;
            14'h302e 	:	o_val <= 16'b0111011001111001;
            14'h302f 	:	o_val <= 16'b0111011001111010;
            14'h3030 	:	o_val <= 16'b0111011001111011;
            14'h3031 	:	o_val <= 16'b0111011001111100;
            14'h3032 	:	o_val <= 16'b0111011001111110;
            14'h3033 	:	o_val <= 16'b0111011001111111;
            14'h3034 	:	o_val <= 16'b0111011010000000;
            14'h3035 	:	o_val <= 16'b0111011010000001;
            14'h3036 	:	o_val <= 16'b0111011010000010;
            14'h3037 	:	o_val <= 16'b0111011010000011;
            14'h3038 	:	o_val <= 16'b0111011010000101;
            14'h3039 	:	o_val <= 16'b0111011010000110;
            14'h303a 	:	o_val <= 16'b0111011010000111;
            14'h303b 	:	o_val <= 16'b0111011010001000;
            14'h303c 	:	o_val <= 16'b0111011010001001;
            14'h303d 	:	o_val <= 16'b0111011010001011;
            14'h303e 	:	o_val <= 16'b0111011010001100;
            14'h303f 	:	o_val <= 16'b0111011010001101;
            14'h3040 	:	o_val <= 16'b0111011010001110;
            14'h3041 	:	o_val <= 16'b0111011010001111;
            14'h3042 	:	o_val <= 16'b0111011010010001;
            14'h3043 	:	o_val <= 16'b0111011010010010;
            14'h3044 	:	o_val <= 16'b0111011010010011;
            14'h3045 	:	o_val <= 16'b0111011010010100;
            14'h3046 	:	o_val <= 16'b0111011010010101;
            14'h3047 	:	o_val <= 16'b0111011010010110;
            14'h3048 	:	o_val <= 16'b0111011010011000;
            14'h3049 	:	o_val <= 16'b0111011010011001;
            14'h304a 	:	o_val <= 16'b0111011010011010;
            14'h304b 	:	o_val <= 16'b0111011010011011;
            14'h304c 	:	o_val <= 16'b0111011010011100;
            14'h304d 	:	o_val <= 16'b0111011010011110;
            14'h304e 	:	o_val <= 16'b0111011010011111;
            14'h304f 	:	o_val <= 16'b0111011010100000;
            14'h3050 	:	o_val <= 16'b0111011010100001;
            14'h3051 	:	o_val <= 16'b0111011010100010;
            14'h3052 	:	o_val <= 16'b0111011010100011;
            14'h3053 	:	o_val <= 16'b0111011010100101;
            14'h3054 	:	o_val <= 16'b0111011010100110;
            14'h3055 	:	o_val <= 16'b0111011010100111;
            14'h3056 	:	o_val <= 16'b0111011010101000;
            14'h3057 	:	o_val <= 16'b0111011010101001;
            14'h3058 	:	o_val <= 16'b0111011010101010;
            14'h3059 	:	o_val <= 16'b0111011010101100;
            14'h305a 	:	o_val <= 16'b0111011010101101;
            14'h305b 	:	o_val <= 16'b0111011010101110;
            14'h305c 	:	o_val <= 16'b0111011010101111;
            14'h305d 	:	o_val <= 16'b0111011010110000;
            14'h305e 	:	o_val <= 16'b0111011010110010;
            14'h305f 	:	o_val <= 16'b0111011010110011;
            14'h3060 	:	o_val <= 16'b0111011010110100;
            14'h3061 	:	o_val <= 16'b0111011010110101;
            14'h3062 	:	o_val <= 16'b0111011010110110;
            14'h3063 	:	o_val <= 16'b0111011010110111;
            14'h3064 	:	o_val <= 16'b0111011010111001;
            14'h3065 	:	o_val <= 16'b0111011010111010;
            14'h3066 	:	o_val <= 16'b0111011010111011;
            14'h3067 	:	o_val <= 16'b0111011010111100;
            14'h3068 	:	o_val <= 16'b0111011010111101;
            14'h3069 	:	o_val <= 16'b0111011010111110;
            14'h306a 	:	o_val <= 16'b0111011011000000;
            14'h306b 	:	o_val <= 16'b0111011011000001;
            14'h306c 	:	o_val <= 16'b0111011011000010;
            14'h306d 	:	o_val <= 16'b0111011011000011;
            14'h306e 	:	o_val <= 16'b0111011011000100;
            14'h306f 	:	o_val <= 16'b0111011011000110;
            14'h3070 	:	o_val <= 16'b0111011011000111;
            14'h3071 	:	o_val <= 16'b0111011011001000;
            14'h3072 	:	o_val <= 16'b0111011011001001;
            14'h3073 	:	o_val <= 16'b0111011011001010;
            14'h3074 	:	o_val <= 16'b0111011011001011;
            14'h3075 	:	o_val <= 16'b0111011011001101;
            14'h3076 	:	o_val <= 16'b0111011011001110;
            14'h3077 	:	o_val <= 16'b0111011011001111;
            14'h3078 	:	o_val <= 16'b0111011011010000;
            14'h3079 	:	o_val <= 16'b0111011011010001;
            14'h307a 	:	o_val <= 16'b0111011011010010;
            14'h307b 	:	o_val <= 16'b0111011011010100;
            14'h307c 	:	o_val <= 16'b0111011011010101;
            14'h307d 	:	o_val <= 16'b0111011011010110;
            14'h307e 	:	o_val <= 16'b0111011011010111;
            14'h307f 	:	o_val <= 16'b0111011011011000;
            14'h3080 	:	o_val <= 16'b0111011011011001;
            14'h3081 	:	o_val <= 16'b0111011011011011;
            14'h3082 	:	o_val <= 16'b0111011011011100;
            14'h3083 	:	o_val <= 16'b0111011011011101;
            14'h3084 	:	o_val <= 16'b0111011011011110;
            14'h3085 	:	o_val <= 16'b0111011011011111;
            14'h3086 	:	o_val <= 16'b0111011011100000;
            14'h3087 	:	o_val <= 16'b0111011011100010;
            14'h3088 	:	o_val <= 16'b0111011011100011;
            14'h3089 	:	o_val <= 16'b0111011011100100;
            14'h308a 	:	o_val <= 16'b0111011011100101;
            14'h308b 	:	o_val <= 16'b0111011011100110;
            14'h308c 	:	o_val <= 16'b0111011011100111;
            14'h308d 	:	o_val <= 16'b0111011011101001;
            14'h308e 	:	o_val <= 16'b0111011011101010;
            14'h308f 	:	o_val <= 16'b0111011011101011;
            14'h3090 	:	o_val <= 16'b0111011011101100;
            14'h3091 	:	o_val <= 16'b0111011011101101;
            14'h3092 	:	o_val <= 16'b0111011011101110;
            14'h3093 	:	o_val <= 16'b0111011011101111;
            14'h3094 	:	o_val <= 16'b0111011011110001;
            14'h3095 	:	o_val <= 16'b0111011011110010;
            14'h3096 	:	o_val <= 16'b0111011011110011;
            14'h3097 	:	o_val <= 16'b0111011011110100;
            14'h3098 	:	o_val <= 16'b0111011011110101;
            14'h3099 	:	o_val <= 16'b0111011011110110;
            14'h309a 	:	o_val <= 16'b0111011011111000;
            14'h309b 	:	o_val <= 16'b0111011011111001;
            14'h309c 	:	o_val <= 16'b0111011011111010;
            14'h309d 	:	o_val <= 16'b0111011011111011;
            14'h309e 	:	o_val <= 16'b0111011011111100;
            14'h309f 	:	o_val <= 16'b0111011011111101;
            14'h30a0 	:	o_val <= 16'b0111011011111111;
            14'h30a1 	:	o_val <= 16'b0111011100000000;
            14'h30a2 	:	o_val <= 16'b0111011100000001;
            14'h30a3 	:	o_val <= 16'b0111011100000010;
            14'h30a4 	:	o_val <= 16'b0111011100000011;
            14'h30a5 	:	o_val <= 16'b0111011100000100;
            14'h30a6 	:	o_val <= 16'b0111011100000101;
            14'h30a7 	:	o_val <= 16'b0111011100000111;
            14'h30a8 	:	o_val <= 16'b0111011100001000;
            14'h30a9 	:	o_val <= 16'b0111011100001001;
            14'h30aa 	:	o_val <= 16'b0111011100001010;
            14'h30ab 	:	o_val <= 16'b0111011100001011;
            14'h30ac 	:	o_val <= 16'b0111011100001100;
            14'h30ad 	:	o_val <= 16'b0111011100001110;
            14'h30ae 	:	o_val <= 16'b0111011100001111;
            14'h30af 	:	o_val <= 16'b0111011100010000;
            14'h30b0 	:	o_val <= 16'b0111011100010001;
            14'h30b1 	:	o_val <= 16'b0111011100010010;
            14'h30b2 	:	o_val <= 16'b0111011100010011;
            14'h30b3 	:	o_val <= 16'b0111011100010100;
            14'h30b4 	:	o_val <= 16'b0111011100010110;
            14'h30b5 	:	o_val <= 16'b0111011100010111;
            14'h30b6 	:	o_val <= 16'b0111011100011000;
            14'h30b7 	:	o_val <= 16'b0111011100011001;
            14'h30b8 	:	o_val <= 16'b0111011100011010;
            14'h30b9 	:	o_val <= 16'b0111011100011011;
            14'h30ba 	:	o_val <= 16'b0111011100011101;
            14'h30bb 	:	o_val <= 16'b0111011100011110;
            14'h30bc 	:	o_val <= 16'b0111011100011111;
            14'h30bd 	:	o_val <= 16'b0111011100100000;
            14'h30be 	:	o_val <= 16'b0111011100100001;
            14'h30bf 	:	o_val <= 16'b0111011100100010;
            14'h30c0 	:	o_val <= 16'b0111011100100011;
            14'h30c1 	:	o_val <= 16'b0111011100100101;
            14'h30c2 	:	o_val <= 16'b0111011100100110;
            14'h30c3 	:	o_val <= 16'b0111011100100111;
            14'h30c4 	:	o_val <= 16'b0111011100101000;
            14'h30c5 	:	o_val <= 16'b0111011100101001;
            14'h30c6 	:	o_val <= 16'b0111011100101010;
            14'h30c7 	:	o_val <= 16'b0111011100101011;
            14'h30c8 	:	o_val <= 16'b0111011100101101;
            14'h30c9 	:	o_val <= 16'b0111011100101110;
            14'h30ca 	:	o_val <= 16'b0111011100101111;
            14'h30cb 	:	o_val <= 16'b0111011100110000;
            14'h30cc 	:	o_val <= 16'b0111011100110001;
            14'h30cd 	:	o_val <= 16'b0111011100110010;
            14'h30ce 	:	o_val <= 16'b0111011100110011;
            14'h30cf 	:	o_val <= 16'b0111011100110101;
            14'h30d0 	:	o_val <= 16'b0111011100110110;
            14'h30d1 	:	o_val <= 16'b0111011100110111;
            14'h30d2 	:	o_val <= 16'b0111011100111000;
            14'h30d3 	:	o_val <= 16'b0111011100111001;
            14'h30d4 	:	o_val <= 16'b0111011100111010;
            14'h30d5 	:	o_val <= 16'b0111011100111100;
            14'h30d6 	:	o_val <= 16'b0111011100111101;
            14'h30d7 	:	o_val <= 16'b0111011100111110;
            14'h30d8 	:	o_val <= 16'b0111011100111111;
            14'h30d9 	:	o_val <= 16'b0111011101000000;
            14'h30da 	:	o_val <= 16'b0111011101000001;
            14'h30db 	:	o_val <= 16'b0111011101000010;
            14'h30dc 	:	o_val <= 16'b0111011101000011;
            14'h30dd 	:	o_val <= 16'b0111011101000101;
            14'h30de 	:	o_val <= 16'b0111011101000110;
            14'h30df 	:	o_val <= 16'b0111011101000111;
            14'h30e0 	:	o_val <= 16'b0111011101001000;
            14'h30e1 	:	o_val <= 16'b0111011101001001;
            14'h30e2 	:	o_val <= 16'b0111011101001010;
            14'h30e3 	:	o_val <= 16'b0111011101001011;
            14'h30e4 	:	o_val <= 16'b0111011101001101;
            14'h30e5 	:	o_val <= 16'b0111011101001110;
            14'h30e6 	:	o_val <= 16'b0111011101001111;
            14'h30e7 	:	o_val <= 16'b0111011101010000;
            14'h30e8 	:	o_val <= 16'b0111011101010001;
            14'h30e9 	:	o_val <= 16'b0111011101010010;
            14'h30ea 	:	o_val <= 16'b0111011101010011;
            14'h30eb 	:	o_val <= 16'b0111011101010101;
            14'h30ec 	:	o_val <= 16'b0111011101010110;
            14'h30ed 	:	o_val <= 16'b0111011101010111;
            14'h30ee 	:	o_val <= 16'b0111011101011000;
            14'h30ef 	:	o_val <= 16'b0111011101011001;
            14'h30f0 	:	o_val <= 16'b0111011101011010;
            14'h30f1 	:	o_val <= 16'b0111011101011011;
            14'h30f2 	:	o_val <= 16'b0111011101011101;
            14'h30f3 	:	o_val <= 16'b0111011101011110;
            14'h30f4 	:	o_val <= 16'b0111011101011111;
            14'h30f5 	:	o_val <= 16'b0111011101100000;
            14'h30f6 	:	o_val <= 16'b0111011101100001;
            14'h30f7 	:	o_val <= 16'b0111011101100010;
            14'h30f8 	:	o_val <= 16'b0111011101100011;
            14'h30f9 	:	o_val <= 16'b0111011101100100;
            14'h30fa 	:	o_val <= 16'b0111011101100110;
            14'h30fb 	:	o_val <= 16'b0111011101100111;
            14'h30fc 	:	o_val <= 16'b0111011101101000;
            14'h30fd 	:	o_val <= 16'b0111011101101001;
            14'h30fe 	:	o_val <= 16'b0111011101101010;
            14'h30ff 	:	o_val <= 16'b0111011101101011;
            14'h3100 	:	o_val <= 16'b0111011101101100;
            14'h3101 	:	o_val <= 16'b0111011101101110;
            14'h3102 	:	o_val <= 16'b0111011101101111;
            14'h3103 	:	o_val <= 16'b0111011101110000;
            14'h3104 	:	o_val <= 16'b0111011101110001;
            14'h3105 	:	o_val <= 16'b0111011101110010;
            14'h3106 	:	o_val <= 16'b0111011101110011;
            14'h3107 	:	o_val <= 16'b0111011101110100;
            14'h3108 	:	o_val <= 16'b0111011101110101;
            14'h3109 	:	o_val <= 16'b0111011101110111;
            14'h310a 	:	o_val <= 16'b0111011101111000;
            14'h310b 	:	o_val <= 16'b0111011101111001;
            14'h310c 	:	o_val <= 16'b0111011101111010;
            14'h310d 	:	o_val <= 16'b0111011101111011;
            14'h310e 	:	o_val <= 16'b0111011101111100;
            14'h310f 	:	o_val <= 16'b0111011101111101;
            14'h3110 	:	o_val <= 16'b0111011101111110;
            14'h3111 	:	o_val <= 16'b0111011110000000;
            14'h3112 	:	o_val <= 16'b0111011110000001;
            14'h3113 	:	o_val <= 16'b0111011110000010;
            14'h3114 	:	o_val <= 16'b0111011110000011;
            14'h3115 	:	o_val <= 16'b0111011110000100;
            14'h3116 	:	o_val <= 16'b0111011110000101;
            14'h3117 	:	o_val <= 16'b0111011110000110;
            14'h3118 	:	o_val <= 16'b0111011110000111;
            14'h3119 	:	o_val <= 16'b0111011110001001;
            14'h311a 	:	o_val <= 16'b0111011110001010;
            14'h311b 	:	o_val <= 16'b0111011110001011;
            14'h311c 	:	o_val <= 16'b0111011110001100;
            14'h311d 	:	o_val <= 16'b0111011110001101;
            14'h311e 	:	o_val <= 16'b0111011110001110;
            14'h311f 	:	o_val <= 16'b0111011110001111;
            14'h3120 	:	o_val <= 16'b0111011110010000;
            14'h3121 	:	o_val <= 16'b0111011110010010;
            14'h3122 	:	o_val <= 16'b0111011110010011;
            14'h3123 	:	o_val <= 16'b0111011110010100;
            14'h3124 	:	o_val <= 16'b0111011110010101;
            14'h3125 	:	o_val <= 16'b0111011110010110;
            14'h3126 	:	o_val <= 16'b0111011110010111;
            14'h3127 	:	o_val <= 16'b0111011110011000;
            14'h3128 	:	o_val <= 16'b0111011110011001;
            14'h3129 	:	o_val <= 16'b0111011110011010;
            14'h312a 	:	o_val <= 16'b0111011110011100;
            14'h312b 	:	o_val <= 16'b0111011110011101;
            14'h312c 	:	o_val <= 16'b0111011110011110;
            14'h312d 	:	o_val <= 16'b0111011110011111;
            14'h312e 	:	o_val <= 16'b0111011110100000;
            14'h312f 	:	o_val <= 16'b0111011110100001;
            14'h3130 	:	o_val <= 16'b0111011110100010;
            14'h3131 	:	o_val <= 16'b0111011110100011;
            14'h3132 	:	o_val <= 16'b0111011110100101;
            14'h3133 	:	o_val <= 16'b0111011110100110;
            14'h3134 	:	o_val <= 16'b0111011110100111;
            14'h3135 	:	o_val <= 16'b0111011110101000;
            14'h3136 	:	o_val <= 16'b0111011110101001;
            14'h3137 	:	o_val <= 16'b0111011110101010;
            14'h3138 	:	o_val <= 16'b0111011110101011;
            14'h3139 	:	o_val <= 16'b0111011110101100;
            14'h313a 	:	o_val <= 16'b0111011110101101;
            14'h313b 	:	o_val <= 16'b0111011110101111;
            14'h313c 	:	o_val <= 16'b0111011110110000;
            14'h313d 	:	o_val <= 16'b0111011110110001;
            14'h313e 	:	o_val <= 16'b0111011110110010;
            14'h313f 	:	o_val <= 16'b0111011110110011;
            14'h3140 	:	o_val <= 16'b0111011110110100;
            14'h3141 	:	o_val <= 16'b0111011110110101;
            14'h3142 	:	o_val <= 16'b0111011110110110;
            14'h3143 	:	o_val <= 16'b0111011110110111;
            14'h3144 	:	o_val <= 16'b0111011110111001;
            14'h3145 	:	o_val <= 16'b0111011110111010;
            14'h3146 	:	o_val <= 16'b0111011110111011;
            14'h3147 	:	o_val <= 16'b0111011110111100;
            14'h3148 	:	o_val <= 16'b0111011110111101;
            14'h3149 	:	o_val <= 16'b0111011110111110;
            14'h314a 	:	o_val <= 16'b0111011110111111;
            14'h314b 	:	o_val <= 16'b0111011111000000;
            14'h314c 	:	o_val <= 16'b0111011111000001;
            14'h314d 	:	o_val <= 16'b0111011111000011;
            14'h314e 	:	o_val <= 16'b0111011111000100;
            14'h314f 	:	o_val <= 16'b0111011111000101;
            14'h3150 	:	o_val <= 16'b0111011111000110;
            14'h3151 	:	o_val <= 16'b0111011111000111;
            14'h3152 	:	o_val <= 16'b0111011111001000;
            14'h3153 	:	o_val <= 16'b0111011111001001;
            14'h3154 	:	o_val <= 16'b0111011111001010;
            14'h3155 	:	o_val <= 16'b0111011111001011;
            14'h3156 	:	o_val <= 16'b0111011111001101;
            14'h3157 	:	o_val <= 16'b0111011111001110;
            14'h3158 	:	o_val <= 16'b0111011111001111;
            14'h3159 	:	o_val <= 16'b0111011111010000;
            14'h315a 	:	o_val <= 16'b0111011111010001;
            14'h315b 	:	o_val <= 16'b0111011111010010;
            14'h315c 	:	o_val <= 16'b0111011111010011;
            14'h315d 	:	o_val <= 16'b0111011111010100;
            14'h315e 	:	o_val <= 16'b0111011111010101;
            14'h315f 	:	o_val <= 16'b0111011111010111;
            14'h3160 	:	o_val <= 16'b0111011111011000;
            14'h3161 	:	o_val <= 16'b0111011111011001;
            14'h3162 	:	o_val <= 16'b0111011111011010;
            14'h3163 	:	o_val <= 16'b0111011111011011;
            14'h3164 	:	o_val <= 16'b0111011111011100;
            14'h3165 	:	o_val <= 16'b0111011111011101;
            14'h3166 	:	o_val <= 16'b0111011111011110;
            14'h3167 	:	o_val <= 16'b0111011111011111;
            14'h3168 	:	o_val <= 16'b0111011111100000;
            14'h3169 	:	o_val <= 16'b0111011111100010;
            14'h316a 	:	o_val <= 16'b0111011111100011;
            14'h316b 	:	o_val <= 16'b0111011111100100;
            14'h316c 	:	o_val <= 16'b0111011111100101;
            14'h316d 	:	o_val <= 16'b0111011111100110;
            14'h316e 	:	o_val <= 16'b0111011111100111;
            14'h316f 	:	o_val <= 16'b0111011111101000;
            14'h3170 	:	o_val <= 16'b0111011111101001;
            14'h3171 	:	o_val <= 16'b0111011111101010;
            14'h3172 	:	o_val <= 16'b0111011111101011;
            14'h3173 	:	o_val <= 16'b0111011111101101;
            14'h3174 	:	o_val <= 16'b0111011111101110;
            14'h3175 	:	o_val <= 16'b0111011111101111;
            14'h3176 	:	o_val <= 16'b0111011111110000;
            14'h3177 	:	o_val <= 16'b0111011111110001;
            14'h3178 	:	o_val <= 16'b0111011111110010;
            14'h3179 	:	o_val <= 16'b0111011111110011;
            14'h317a 	:	o_val <= 16'b0111011111110100;
            14'h317b 	:	o_val <= 16'b0111011111110101;
            14'h317c 	:	o_val <= 16'b0111011111110110;
            14'h317d 	:	o_val <= 16'b0111011111110111;
            14'h317e 	:	o_val <= 16'b0111011111111001;
            14'h317f 	:	o_val <= 16'b0111011111111010;
            14'h3180 	:	o_val <= 16'b0111011111111011;
            14'h3181 	:	o_val <= 16'b0111011111111100;
            14'h3182 	:	o_val <= 16'b0111011111111101;
            14'h3183 	:	o_val <= 16'b0111011111111110;
            14'h3184 	:	o_val <= 16'b0111011111111111;
            14'h3185 	:	o_val <= 16'b0111100000000000;
            14'h3186 	:	o_val <= 16'b0111100000000001;
            14'h3187 	:	o_val <= 16'b0111100000000010;
            14'h3188 	:	o_val <= 16'b0111100000000100;
            14'h3189 	:	o_val <= 16'b0111100000000101;
            14'h318a 	:	o_val <= 16'b0111100000000110;
            14'h318b 	:	o_val <= 16'b0111100000000111;
            14'h318c 	:	o_val <= 16'b0111100000001000;
            14'h318d 	:	o_val <= 16'b0111100000001001;
            14'h318e 	:	o_val <= 16'b0111100000001010;
            14'h318f 	:	o_val <= 16'b0111100000001011;
            14'h3190 	:	o_val <= 16'b0111100000001100;
            14'h3191 	:	o_val <= 16'b0111100000001101;
            14'h3192 	:	o_val <= 16'b0111100000001110;
            14'h3193 	:	o_val <= 16'b0111100000010000;
            14'h3194 	:	o_val <= 16'b0111100000010001;
            14'h3195 	:	o_val <= 16'b0111100000010010;
            14'h3196 	:	o_val <= 16'b0111100000010011;
            14'h3197 	:	o_val <= 16'b0111100000010100;
            14'h3198 	:	o_val <= 16'b0111100000010101;
            14'h3199 	:	o_val <= 16'b0111100000010110;
            14'h319a 	:	o_val <= 16'b0111100000010111;
            14'h319b 	:	o_val <= 16'b0111100000011000;
            14'h319c 	:	o_val <= 16'b0111100000011001;
            14'h319d 	:	o_val <= 16'b0111100000011010;
            14'h319e 	:	o_val <= 16'b0111100000011011;
            14'h319f 	:	o_val <= 16'b0111100000011101;
            14'h31a0 	:	o_val <= 16'b0111100000011110;
            14'h31a1 	:	o_val <= 16'b0111100000011111;
            14'h31a2 	:	o_val <= 16'b0111100000100000;
            14'h31a3 	:	o_val <= 16'b0111100000100001;
            14'h31a4 	:	o_val <= 16'b0111100000100010;
            14'h31a5 	:	o_val <= 16'b0111100000100011;
            14'h31a6 	:	o_val <= 16'b0111100000100100;
            14'h31a7 	:	o_val <= 16'b0111100000100101;
            14'h31a8 	:	o_val <= 16'b0111100000100110;
            14'h31a9 	:	o_val <= 16'b0111100000100111;
            14'h31aa 	:	o_val <= 16'b0111100000101000;
            14'h31ab 	:	o_val <= 16'b0111100000101010;
            14'h31ac 	:	o_val <= 16'b0111100000101011;
            14'h31ad 	:	o_val <= 16'b0111100000101100;
            14'h31ae 	:	o_val <= 16'b0111100000101101;
            14'h31af 	:	o_val <= 16'b0111100000101110;
            14'h31b0 	:	o_val <= 16'b0111100000101111;
            14'h31b1 	:	o_val <= 16'b0111100000110000;
            14'h31b2 	:	o_val <= 16'b0111100000110001;
            14'h31b3 	:	o_val <= 16'b0111100000110010;
            14'h31b4 	:	o_val <= 16'b0111100000110011;
            14'h31b5 	:	o_val <= 16'b0111100000110100;
            14'h31b6 	:	o_val <= 16'b0111100000110101;
            14'h31b7 	:	o_val <= 16'b0111100000110111;
            14'h31b8 	:	o_val <= 16'b0111100000111000;
            14'h31b9 	:	o_val <= 16'b0111100000111001;
            14'h31ba 	:	o_val <= 16'b0111100000111010;
            14'h31bb 	:	o_val <= 16'b0111100000111011;
            14'h31bc 	:	o_val <= 16'b0111100000111100;
            14'h31bd 	:	o_val <= 16'b0111100000111101;
            14'h31be 	:	o_val <= 16'b0111100000111110;
            14'h31bf 	:	o_val <= 16'b0111100000111111;
            14'h31c0 	:	o_val <= 16'b0111100001000000;
            14'h31c1 	:	o_val <= 16'b0111100001000001;
            14'h31c2 	:	o_val <= 16'b0111100001000010;
            14'h31c3 	:	o_val <= 16'b0111100001000011;
            14'h31c4 	:	o_val <= 16'b0111100001000101;
            14'h31c5 	:	o_val <= 16'b0111100001000110;
            14'h31c6 	:	o_val <= 16'b0111100001000111;
            14'h31c7 	:	o_val <= 16'b0111100001001000;
            14'h31c8 	:	o_val <= 16'b0111100001001001;
            14'h31c9 	:	o_val <= 16'b0111100001001010;
            14'h31ca 	:	o_val <= 16'b0111100001001011;
            14'h31cb 	:	o_val <= 16'b0111100001001100;
            14'h31cc 	:	o_val <= 16'b0111100001001101;
            14'h31cd 	:	o_val <= 16'b0111100001001110;
            14'h31ce 	:	o_val <= 16'b0111100001001111;
            14'h31cf 	:	o_val <= 16'b0111100001010000;
            14'h31d0 	:	o_val <= 16'b0111100001010001;
            14'h31d1 	:	o_val <= 16'b0111100001010010;
            14'h31d2 	:	o_val <= 16'b0111100001010100;
            14'h31d3 	:	o_val <= 16'b0111100001010101;
            14'h31d4 	:	o_val <= 16'b0111100001010110;
            14'h31d5 	:	o_val <= 16'b0111100001010111;
            14'h31d6 	:	o_val <= 16'b0111100001011000;
            14'h31d7 	:	o_val <= 16'b0111100001011001;
            14'h31d8 	:	o_val <= 16'b0111100001011010;
            14'h31d9 	:	o_val <= 16'b0111100001011011;
            14'h31da 	:	o_val <= 16'b0111100001011100;
            14'h31db 	:	o_val <= 16'b0111100001011101;
            14'h31dc 	:	o_val <= 16'b0111100001011110;
            14'h31dd 	:	o_val <= 16'b0111100001011111;
            14'h31de 	:	o_val <= 16'b0111100001100000;
            14'h31df 	:	o_val <= 16'b0111100001100001;
            14'h31e0 	:	o_val <= 16'b0111100001100011;
            14'h31e1 	:	o_val <= 16'b0111100001100100;
            14'h31e2 	:	o_val <= 16'b0111100001100101;
            14'h31e3 	:	o_val <= 16'b0111100001100110;
            14'h31e4 	:	o_val <= 16'b0111100001100111;
            14'h31e5 	:	o_val <= 16'b0111100001101000;
            14'h31e6 	:	o_val <= 16'b0111100001101001;
            14'h31e7 	:	o_val <= 16'b0111100001101010;
            14'h31e8 	:	o_val <= 16'b0111100001101011;
            14'h31e9 	:	o_val <= 16'b0111100001101100;
            14'h31ea 	:	o_val <= 16'b0111100001101101;
            14'h31eb 	:	o_val <= 16'b0111100001101110;
            14'h31ec 	:	o_val <= 16'b0111100001101111;
            14'h31ed 	:	o_val <= 16'b0111100001110000;
            14'h31ee 	:	o_val <= 16'b0111100001110001;
            14'h31ef 	:	o_val <= 16'b0111100001110011;
            14'h31f0 	:	o_val <= 16'b0111100001110100;
            14'h31f1 	:	o_val <= 16'b0111100001110101;
            14'h31f2 	:	o_val <= 16'b0111100001110110;
            14'h31f3 	:	o_val <= 16'b0111100001110111;
            14'h31f4 	:	o_val <= 16'b0111100001111000;
            14'h31f5 	:	o_val <= 16'b0111100001111001;
            14'h31f6 	:	o_val <= 16'b0111100001111010;
            14'h31f7 	:	o_val <= 16'b0111100001111011;
            14'h31f8 	:	o_val <= 16'b0111100001111100;
            14'h31f9 	:	o_val <= 16'b0111100001111101;
            14'h31fa 	:	o_val <= 16'b0111100001111110;
            14'h31fb 	:	o_val <= 16'b0111100001111111;
            14'h31fc 	:	o_val <= 16'b0111100010000000;
            14'h31fd 	:	o_val <= 16'b0111100010000001;
            14'h31fe 	:	o_val <= 16'b0111100010000010;
            14'h31ff 	:	o_val <= 16'b0111100010000011;
            14'h3200 	:	o_val <= 16'b0111100010000101;
            14'h3201 	:	o_val <= 16'b0111100010000110;
            14'h3202 	:	o_val <= 16'b0111100010000111;
            14'h3203 	:	o_val <= 16'b0111100010001000;
            14'h3204 	:	o_val <= 16'b0111100010001001;
            14'h3205 	:	o_val <= 16'b0111100010001010;
            14'h3206 	:	o_val <= 16'b0111100010001011;
            14'h3207 	:	o_val <= 16'b0111100010001100;
            14'h3208 	:	o_val <= 16'b0111100010001101;
            14'h3209 	:	o_val <= 16'b0111100010001110;
            14'h320a 	:	o_val <= 16'b0111100010001111;
            14'h320b 	:	o_val <= 16'b0111100010010000;
            14'h320c 	:	o_val <= 16'b0111100010010001;
            14'h320d 	:	o_val <= 16'b0111100010010010;
            14'h320e 	:	o_val <= 16'b0111100010010011;
            14'h320f 	:	o_val <= 16'b0111100010010100;
            14'h3210 	:	o_val <= 16'b0111100010010101;
            14'h3211 	:	o_val <= 16'b0111100010010110;
            14'h3212 	:	o_val <= 16'b0111100010011000;
            14'h3213 	:	o_val <= 16'b0111100010011001;
            14'h3214 	:	o_val <= 16'b0111100010011010;
            14'h3215 	:	o_val <= 16'b0111100010011011;
            14'h3216 	:	o_val <= 16'b0111100010011100;
            14'h3217 	:	o_val <= 16'b0111100010011101;
            14'h3218 	:	o_val <= 16'b0111100010011110;
            14'h3219 	:	o_val <= 16'b0111100010011111;
            14'h321a 	:	o_val <= 16'b0111100010100000;
            14'h321b 	:	o_val <= 16'b0111100010100001;
            14'h321c 	:	o_val <= 16'b0111100010100010;
            14'h321d 	:	o_val <= 16'b0111100010100011;
            14'h321e 	:	o_val <= 16'b0111100010100100;
            14'h321f 	:	o_val <= 16'b0111100010100101;
            14'h3220 	:	o_val <= 16'b0111100010100110;
            14'h3221 	:	o_val <= 16'b0111100010100111;
            14'h3222 	:	o_val <= 16'b0111100010101000;
            14'h3223 	:	o_val <= 16'b0111100010101001;
            14'h3224 	:	o_val <= 16'b0111100010101010;
            14'h3225 	:	o_val <= 16'b0111100010101100;
            14'h3226 	:	o_val <= 16'b0111100010101101;
            14'h3227 	:	o_val <= 16'b0111100010101110;
            14'h3228 	:	o_val <= 16'b0111100010101111;
            14'h3229 	:	o_val <= 16'b0111100010110000;
            14'h322a 	:	o_val <= 16'b0111100010110001;
            14'h322b 	:	o_val <= 16'b0111100010110010;
            14'h322c 	:	o_val <= 16'b0111100010110011;
            14'h322d 	:	o_val <= 16'b0111100010110100;
            14'h322e 	:	o_val <= 16'b0111100010110101;
            14'h322f 	:	o_val <= 16'b0111100010110110;
            14'h3230 	:	o_val <= 16'b0111100010110111;
            14'h3231 	:	o_val <= 16'b0111100010111000;
            14'h3232 	:	o_val <= 16'b0111100010111001;
            14'h3233 	:	o_val <= 16'b0111100010111010;
            14'h3234 	:	o_val <= 16'b0111100010111011;
            14'h3235 	:	o_val <= 16'b0111100010111100;
            14'h3236 	:	o_val <= 16'b0111100010111101;
            14'h3237 	:	o_val <= 16'b0111100010111110;
            14'h3238 	:	o_val <= 16'b0111100010111111;
            14'h3239 	:	o_val <= 16'b0111100011000000;
            14'h323a 	:	o_val <= 16'b0111100011000001;
            14'h323b 	:	o_val <= 16'b0111100011000010;
            14'h323c 	:	o_val <= 16'b0111100011000100;
            14'h323d 	:	o_val <= 16'b0111100011000101;
            14'h323e 	:	o_val <= 16'b0111100011000110;
            14'h323f 	:	o_val <= 16'b0111100011000111;
            14'h3240 	:	o_val <= 16'b0111100011001000;
            14'h3241 	:	o_val <= 16'b0111100011001001;
            14'h3242 	:	o_val <= 16'b0111100011001010;
            14'h3243 	:	o_val <= 16'b0111100011001011;
            14'h3244 	:	o_val <= 16'b0111100011001100;
            14'h3245 	:	o_val <= 16'b0111100011001101;
            14'h3246 	:	o_val <= 16'b0111100011001110;
            14'h3247 	:	o_val <= 16'b0111100011001111;
            14'h3248 	:	o_val <= 16'b0111100011010000;
            14'h3249 	:	o_val <= 16'b0111100011010001;
            14'h324a 	:	o_val <= 16'b0111100011010010;
            14'h324b 	:	o_val <= 16'b0111100011010011;
            14'h324c 	:	o_val <= 16'b0111100011010100;
            14'h324d 	:	o_val <= 16'b0111100011010101;
            14'h324e 	:	o_val <= 16'b0111100011010110;
            14'h324f 	:	o_val <= 16'b0111100011010111;
            14'h3250 	:	o_val <= 16'b0111100011011000;
            14'h3251 	:	o_val <= 16'b0111100011011001;
            14'h3252 	:	o_val <= 16'b0111100011011010;
            14'h3253 	:	o_val <= 16'b0111100011011011;
            14'h3254 	:	o_val <= 16'b0111100011011100;
            14'h3255 	:	o_val <= 16'b0111100011011101;
            14'h3256 	:	o_val <= 16'b0111100011011111;
            14'h3257 	:	o_val <= 16'b0111100011100000;
            14'h3258 	:	o_val <= 16'b0111100011100001;
            14'h3259 	:	o_val <= 16'b0111100011100010;
            14'h325a 	:	o_val <= 16'b0111100011100011;
            14'h325b 	:	o_val <= 16'b0111100011100100;
            14'h325c 	:	o_val <= 16'b0111100011100101;
            14'h325d 	:	o_val <= 16'b0111100011100110;
            14'h325e 	:	o_val <= 16'b0111100011100111;
            14'h325f 	:	o_val <= 16'b0111100011101000;
            14'h3260 	:	o_val <= 16'b0111100011101001;
            14'h3261 	:	o_val <= 16'b0111100011101010;
            14'h3262 	:	o_val <= 16'b0111100011101011;
            14'h3263 	:	o_val <= 16'b0111100011101100;
            14'h3264 	:	o_val <= 16'b0111100011101101;
            14'h3265 	:	o_val <= 16'b0111100011101110;
            14'h3266 	:	o_val <= 16'b0111100011101111;
            14'h3267 	:	o_val <= 16'b0111100011110000;
            14'h3268 	:	o_val <= 16'b0111100011110001;
            14'h3269 	:	o_val <= 16'b0111100011110010;
            14'h326a 	:	o_val <= 16'b0111100011110011;
            14'h326b 	:	o_val <= 16'b0111100011110100;
            14'h326c 	:	o_val <= 16'b0111100011110101;
            14'h326d 	:	o_val <= 16'b0111100011110110;
            14'h326e 	:	o_val <= 16'b0111100011110111;
            14'h326f 	:	o_val <= 16'b0111100011111000;
            14'h3270 	:	o_val <= 16'b0111100011111001;
            14'h3271 	:	o_val <= 16'b0111100011111010;
            14'h3272 	:	o_val <= 16'b0111100011111011;
            14'h3273 	:	o_val <= 16'b0111100011111100;
            14'h3274 	:	o_val <= 16'b0111100011111101;
            14'h3275 	:	o_val <= 16'b0111100011111110;
            14'h3276 	:	o_val <= 16'b0111100011111111;
            14'h3277 	:	o_val <= 16'b0111100100000000;
            14'h3278 	:	o_val <= 16'b0111100100000001;
            14'h3279 	:	o_val <= 16'b0111100100000011;
            14'h327a 	:	o_val <= 16'b0111100100000100;
            14'h327b 	:	o_val <= 16'b0111100100000101;
            14'h327c 	:	o_val <= 16'b0111100100000110;
            14'h327d 	:	o_val <= 16'b0111100100000111;
            14'h327e 	:	o_val <= 16'b0111100100001000;
            14'h327f 	:	o_val <= 16'b0111100100001001;
            14'h3280 	:	o_val <= 16'b0111100100001010;
            14'h3281 	:	o_val <= 16'b0111100100001011;
            14'h3282 	:	o_val <= 16'b0111100100001100;
            14'h3283 	:	o_val <= 16'b0111100100001101;
            14'h3284 	:	o_val <= 16'b0111100100001110;
            14'h3285 	:	o_val <= 16'b0111100100001111;
            14'h3286 	:	o_val <= 16'b0111100100010000;
            14'h3287 	:	o_val <= 16'b0111100100010001;
            14'h3288 	:	o_val <= 16'b0111100100010010;
            14'h3289 	:	o_val <= 16'b0111100100010011;
            14'h328a 	:	o_val <= 16'b0111100100010100;
            14'h328b 	:	o_val <= 16'b0111100100010101;
            14'h328c 	:	o_val <= 16'b0111100100010110;
            14'h328d 	:	o_val <= 16'b0111100100010111;
            14'h328e 	:	o_val <= 16'b0111100100011000;
            14'h328f 	:	o_val <= 16'b0111100100011001;
            14'h3290 	:	o_val <= 16'b0111100100011010;
            14'h3291 	:	o_val <= 16'b0111100100011011;
            14'h3292 	:	o_val <= 16'b0111100100011100;
            14'h3293 	:	o_val <= 16'b0111100100011101;
            14'h3294 	:	o_val <= 16'b0111100100011110;
            14'h3295 	:	o_val <= 16'b0111100100011111;
            14'h3296 	:	o_val <= 16'b0111100100100000;
            14'h3297 	:	o_val <= 16'b0111100100100001;
            14'h3298 	:	o_val <= 16'b0111100100100010;
            14'h3299 	:	o_val <= 16'b0111100100100011;
            14'h329a 	:	o_val <= 16'b0111100100100100;
            14'h329b 	:	o_val <= 16'b0111100100100101;
            14'h329c 	:	o_val <= 16'b0111100100100110;
            14'h329d 	:	o_val <= 16'b0111100100100111;
            14'h329e 	:	o_val <= 16'b0111100100101000;
            14'h329f 	:	o_val <= 16'b0111100100101001;
            14'h32a0 	:	o_val <= 16'b0111100100101010;
            14'h32a1 	:	o_val <= 16'b0111100100101011;
            14'h32a2 	:	o_val <= 16'b0111100100101100;
            14'h32a3 	:	o_val <= 16'b0111100100101101;
            14'h32a4 	:	o_val <= 16'b0111100100101110;
            14'h32a5 	:	o_val <= 16'b0111100100101111;
            14'h32a6 	:	o_val <= 16'b0111100100110000;
            14'h32a7 	:	o_val <= 16'b0111100100110001;
            14'h32a8 	:	o_val <= 16'b0111100100110010;
            14'h32a9 	:	o_val <= 16'b0111100100110011;
            14'h32aa 	:	o_val <= 16'b0111100100110100;
            14'h32ab 	:	o_val <= 16'b0111100100110101;
            14'h32ac 	:	o_val <= 16'b0111100100110110;
            14'h32ad 	:	o_val <= 16'b0111100100110111;
            14'h32ae 	:	o_val <= 16'b0111100100111000;
            14'h32af 	:	o_val <= 16'b0111100100111001;
            14'h32b0 	:	o_val <= 16'b0111100100111010;
            14'h32b1 	:	o_val <= 16'b0111100100111011;
            14'h32b2 	:	o_val <= 16'b0111100100111100;
            14'h32b3 	:	o_val <= 16'b0111100100111101;
            14'h32b4 	:	o_val <= 16'b0111100100111110;
            14'h32b5 	:	o_val <= 16'b0111100100111111;
            14'h32b6 	:	o_val <= 16'b0111100101000000;
            14'h32b7 	:	o_val <= 16'b0111100101000001;
            14'h32b8 	:	o_val <= 16'b0111100101000010;
            14'h32b9 	:	o_val <= 16'b0111100101000011;
            14'h32ba 	:	o_val <= 16'b0111100101000100;
            14'h32bb 	:	o_val <= 16'b0111100101000101;
            14'h32bc 	:	o_val <= 16'b0111100101000110;
            14'h32bd 	:	o_val <= 16'b0111100101000111;
            14'h32be 	:	o_val <= 16'b0111100101001000;
            14'h32bf 	:	o_val <= 16'b0111100101001001;
            14'h32c0 	:	o_val <= 16'b0111100101001010;
            14'h32c1 	:	o_val <= 16'b0111100101001011;
            14'h32c2 	:	o_val <= 16'b0111100101001100;
            14'h32c3 	:	o_val <= 16'b0111100101001101;
            14'h32c4 	:	o_val <= 16'b0111100101001110;
            14'h32c5 	:	o_val <= 16'b0111100101010000;
            14'h32c6 	:	o_val <= 16'b0111100101010001;
            14'h32c7 	:	o_val <= 16'b0111100101010010;
            14'h32c8 	:	o_val <= 16'b0111100101010011;
            14'h32c9 	:	o_val <= 16'b0111100101010100;
            14'h32ca 	:	o_val <= 16'b0111100101010101;
            14'h32cb 	:	o_val <= 16'b0111100101010110;
            14'h32cc 	:	o_val <= 16'b0111100101010111;
            14'h32cd 	:	o_val <= 16'b0111100101011000;
            14'h32ce 	:	o_val <= 16'b0111100101011001;
            14'h32cf 	:	o_val <= 16'b0111100101011010;
            14'h32d0 	:	o_val <= 16'b0111100101011011;
            14'h32d1 	:	o_val <= 16'b0111100101011100;
            14'h32d2 	:	o_val <= 16'b0111100101011101;
            14'h32d3 	:	o_val <= 16'b0111100101011110;
            14'h32d4 	:	o_val <= 16'b0111100101011111;
            14'h32d5 	:	o_val <= 16'b0111100101011111;
            14'h32d6 	:	o_val <= 16'b0111100101100000;
            14'h32d7 	:	o_val <= 16'b0111100101100001;
            14'h32d8 	:	o_val <= 16'b0111100101100010;
            14'h32d9 	:	o_val <= 16'b0111100101100011;
            14'h32da 	:	o_val <= 16'b0111100101100100;
            14'h32db 	:	o_val <= 16'b0111100101100101;
            14'h32dc 	:	o_val <= 16'b0111100101100110;
            14'h32dd 	:	o_val <= 16'b0111100101100111;
            14'h32de 	:	o_val <= 16'b0111100101101000;
            14'h32df 	:	o_val <= 16'b0111100101101001;
            14'h32e0 	:	o_val <= 16'b0111100101101010;
            14'h32e1 	:	o_val <= 16'b0111100101101011;
            14'h32e2 	:	o_val <= 16'b0111100101101100;
            14'h32e3 	:	o_val <= 16'b0111100101101101;
            14'h32e4 	:	o_val <= 16'b0111100101101110;
            14'h32e5 	:	o_val <= 16'b0111100101101111;
            14'h32e6 	:	o_val <= 16'b0111100101110000;
            14'h32e7 	:	o_val <= 16'b0111100101110001;
            14'h32e8 	:	o_val <= 16'b0111100101110010;
            14'h32e9 	:	o_val <= 16'b0111100101110011;
            14'h32ea 	:	o_val <= 16'b0111100101110100;
            14'h32eb 	:	o_val <= 16'b0111100101110101;
            14'h32ec 	:	o_val <= 16'b0111100101110110;
            14'h32ed 	:	o_val <= 16'b0111100101110111;
            14'h32ee 	:	o_val <= 16'b0111100101111000;
            14'h32ef 	:	o_val <= 16'b0111100101111001;
            14'h32f0 	:	o_val <= 16'b0111100101111010;
            14'h32f1 	:	o_val <= 16'b0111100101111011;
            14'h32f2 	:	o_val <= 16'b0111100101111100;
            14'h32f3 	:	o_val <= 16'b0111100101111101;
            14'h32f4 	:	o_val <= 16'b0111100101111110;
            14'h32f5 	:	o_val <= 16'b0111100101111111;
            14'h32f6 	:	o_val <= 16'b0111100110000000;
            14'h32f7 	:	o_val <= 16'b0111100110000001;
            14'h32f8 	:	o_val <= 16'b0111100110000010;
            14'h32f9 	:	o_val <= 16'b0111100110000011;
            14'h32fa 	:	o_val <= 16'b0111100110000100;
            14'h32fb 	:	o_val <= 16'b0111100110000101;
            14'h32fc 	:	o_val <= 16'b0111100110000110;
            14'h32fd 	:	o_val <= 16'b0111100110000111;
            14'h32fe 	:	o_val <= 16'b0111100110001000;
            14'h32ff 	:	o_val <= 16'b0111100110001001;
            14'h3300 	:	o_val <= 16'b0111100110001010;
            14'h3301 	:	o_val <= 16'b0111100110001011;
            14'h3302 	:	o_val <= 16'b0111100110001100;
            14'h3303 	:	o_val <= 16'b0111100110001101;
            14'h3304 	:	o_val <= 16'b0111100110001110;
            14'h3305 	:	o_val <= 16'b0111100110001111;
            14'h3306 	:	o_val <= 16'b0111100110010000;
            14'h3307 	:	o_val <= 16'b0111100110010001;
            14'h3308 	:	o_val <= 16'b0111100110010010;
            14'h3309 	:	o_val <= 16'b0111100110010011;
            14'h330a 	:	o_val <= 16'b0111100110010100;
            14'h330b 	:	o_val <= 16'b0111100110010101;
            14'h330c 	:	o_val <= 16'b0111100110010110;
            14'h330d 	:	o_val <= 16'b0111100110010111;
            14'h330e 	:	o_val <= 16'b0111100110011000;
            14'h330f 	:	o_val <= 16'b0111100110011001;
            14'h3310 	:	o_val <= 16'b0111100110011010;
            14'h3311 	:	o_val <= 16'b0111100110011011;
            14'h3312 	:	o_val <= 16'b0111100110011100;
            14'h3313 	:	o_val <= 16'b0111100110011101;
            14'h3314 	:	o_val <= 16'b0111100110011110;
            14'h3315 	:	o_val <= 16'b0111100110011111;
            14'h3316 	:	o_val <= 16'b0111100110100000;
            14'h3317 	:	o_val <= 16'b0111100110100001;
            14'h3318 	:	o_val <= 16'b0111100110100010;
            14'h3319 	:	o_val <= 16'b0111100110100011;
            14'h331a 	:	o_val <= 16'b0111100110100100;
            14'h331b 	:	o_val <= 16'b0111100110100101;
            14'h331c 	:	o_val <= 16'b0111100110100110;
            14'h331d 	:	o_val <= 16'b0111100110100111;
            14'h331e 	:	o_val <= 16'b0111100110101000;
            14'h331f 	:	o_val <= 16'b0111100110101001;
            14'h3320 	:	o_val <= 16'b0111100110101010;
            14'h3321 	:	o_val <= 16'b0111100110101010;
            14'h3322 	:	o_val <= 16'b0111100110101011;
            14'h3323 	:	o_val <= 16'b0111100110101100;
            14'h3324 	:	o_val <= 16'b0111100110101101;
            14'h3325 	:	o_val <= 16'b0111100110101110;
            14'h3326 	:	o_val <= 16'b0111100110101111;
            14'h3327 	:	o_val <= 16'b0111100110110000;
            14'h3328 	:	o_val <= 16'b0111100110110001;
            14'h3329 	:	o_val <= 16'b0111100110110010;
            14'h332a 	:	o_val <= 16'b0111100110110011;
            14'h332b 	:	o_val <= 16'b0111100110110100;
            14'h332c 	:	o_val <= 16'b0111100110110101;
            14'h332d 	:	o_val <= 16'b0111100110110110;
            14'h332e 	:	o_val <= 16'b0111100110110111;
            14'h332f 	:	o_val <= 16'b0111100110111000;
            14'h3330 	:	o_val <= 16'b0111100110111001;
            14'h3331 	:	o_val <= 16'b0111100110111010;
            14'h3332 	:	o_val <= 16'b0111100110111011;
            14'h3333 	:	o_val <= 16'b0111100110111100;
            14'h3334 	:	o_val <= 16'b0111100110111101;
            14'h3335 	:	o_val <= 16'b0111100110111110;
            14'h3336 	:	o_val <= 16'b0111100110111111;
            14'h3337 	:	o_val <= 16'b0111100111000000;
            14'h3338 	:	o_val <= 16'b0111100111000001;
            14'h3339 	:	o_val <= 16'b0111100111000010;
            14'h333a 	:	o_val <= 16'b0111100111000011;
            14'h333b 	:	o_val <= 16'b0111100111000100;
            14'h333c 	:	o_val <= 16'b0111100111000101;
            14'h333d 	:	o_val <= 16'b0111100111000110;
            14'h333e 	:	o_val <= 16'b0111100111000111;
            14'h333f 	:	o_val <= 16'b0111100111001000;
            14'h3340 	:	o_val <= 16'b0111100111001001;
            14'h3341 	:	o_val <= 16'b0111100111001010;
            14'h3342 	:	o_val <= 16'b0111100111001011;
            14'h3343 	:	o_val <= 16'b0111100111001100;
            14'h3344 	:	o_val <= 16'b0111100111001100;
            14'h3345 	:	o_val <= 16'b0111100111001101;
            14'h3346 	:	o_val <= 16'b0111100111001110;
            14'h3347 	:	o_val <= 16'b0111100111001111;
            14'h3348 	:	o_val <= 16'b0111100111010000;
            14'h3349 	:	o_val <= 16'b0111100111010001;
            14'h334a 	:	o_val <= 16'b0111100111010010;
            14'h334b 	:	o_val <= 16'b0111100111010011;
            14'h334c 	:	o_val <= 16'b0111100111010100;
            14'h334d 	:	o_val <= 16'b0111100111010101;
            14'h334e 	:	o_val <= 16'b0111100111010110;
            14'h334f 	:	o_val <= 16'b0111100111010111;
            14'h3350 	:	o_val <= 16'b0111100111011000;
            14'h3351 	:	o_val <= 16'b0111100111011001;
            14'h3352 	:	o_val <= 16'b0111100111011010;
            14'h3353 	:	o_val <= 16'b0111100111011011;
            14'h3354 	:	o_val <= 16'b0111100111011100;
            14'h3355 	:	o_val <= 16'b0111100111011101;
            14'h3356 	:	o_val <= 16'b0111100111011110;
            14'h3357 	:	o_val <= 16'b0111100111011111;
            14'h3358 	:	o_val <= 16'b0111100111100000;
            14'h3359 	:	o_val <= 16'b0111100111100001;
            14'h335a 	:	o_val <= 16'b0111100111100010;
            14'h335b 	:	o_val <= 16'b0111100111100011;
            14'h335c 	:	o_val <= 16'b0111100111100100;
            14'h335d 	:	o_val <= 16'b0111100111100101;
            14'h335e 	:	o_val <= 16'b0111100111100101;
            14'h335f 	:	o_val <= 16'b0111100111100110;
            14'h3360 	:	o_val <= 16'b0111100111100111;
            14'h3361 	:	o_val <= 16'b0111100111101000;
            14'h3362 	:	o_val <= 16'b0111100111101001;
            14'h3363 	:	o_val <= 16'b0111100111101010;
            14'h3364 	:	o_val <= 16'b0111100111101011;
            14'h3365 	:	o_val <= 16'b0111100111101100;
            14'h3366 	:	o_val <= 16'b0111100111101101;
            14'h3367 	:	o_val <= 16'b0111100111101110;
            14'h3368 	:	o_val <= 16'b0111100111101111;
            14'h3369 	:	o_val <= 16'b0111100111110000;
            14'h336a 	:	o_val <= 16'b0111100111110001;
            14'h336b 	:	o_val <= 16'b0111100111110010;
            14'h336c 	:	o_val <= 16'b0111100111110011;
            14'h336d 	:	o_val <= 16'b0111100111110100;
            14'h336e 	:	o_val <= 16'b0111100111110101;
            14'h336f 	:	o_val <= 16'b0111100111110110;
            14'h3370 	:	o_val <= 16'b0111100111110111;
            14'h3371 	:	o_val <= 16'b0111100111111000;
            14'h3372 	:	o_val <= 16'b0111100111111001;
            14'h3373 	:	o_val <= 16'b0111100111111010;
            14'h3374 	:	o_val <= 16'b0111100111111011;
            14'h3375 	:	o_val <= 16'b0111100111111011;
            14'h3376 	:	o_val <= 16'b0111100111111100;
            14'h3377 	:	o_val <= 16'b0111100111111101;
            14'h3378 	:	o_val <= 16'b0111100111111110;
            14'h3379 	:	o_val <= 16'b0111100111111111;
            14'h337a 	:	o_val <= 16'b0111101000000000;
            14'h337b 	:	o_val <= 16'b0111101000000001;
            14'h337c 	:	o_val <= 16'b0111101000000010;
            14'h337d 	:	o_val <= 16'b0111101000000011;
            14'h337e 	:	o_val <= 16'b0111101000000100;
            14'h337f 	:	o_val <= 16'b0111101000000101;
            14'h3380 	:	o_val <= 16'b0111101000000110;
            14'h3381 	:	o_val <= 16'b0111101000000111;
            14'h3382 	:	o_val <= 16'b0111101000001000;
            14'h3383 	:	o_val <= 16'b0111101000001001;
            14'h3384 	:	o_val <= 16'b0111101000001010;
            14'h3385 	:	o_val <= 16'b0111101000001011;
            14'h3386 	:	o_val <= 16'b0111101000001100;
            14'h3387 	:	o_val <= 16'b0111101000001101;
            14'h3388 	:	o_val <= 16'b0111101000001101;
            14'h3389 	:	o_val <= 16'b0111101000001110;
            14'h338a 	:	o_val <= 16'b0111101000001111;
            14'h338b 	:	o_val <= 16'b0111101000010000;
            14'h338c 	:	o_val <= 16'b0111101000010001;
            14'h338d 	:	o_val <= 16'b0111101000010010;
            14'h338e 	:	o_val <= 16'b0111101000010011;
            14'h338f 	:	o_val <= 16'b0111101000010100;
            14'h3390 	:	o_val <= 16'b0111101000010101;
            14'h3391 	:	o_val <= 16'b0111101000010110;
            14'h3392 	:	o_val <= 16'b0111101000010111;
            14'h3393 	:	o_val <= 16'b0111101000011000;
            14'h3394 	:	o_val <= 16'b0111101000011001;
            14'h3395 	:	o_val <= 16'b0111101000011010;
            14'h3396 	:	o_val <= 16'b0111101000011011;
            14'h3397 	:	o_val <= 16'b0111101000011100;
            14'h3398 	:	o_val <= 16'b0111101000011101;
            14'h3399 	:	o_val <= 16'b0111101000011110;
            14'h339a 	:	o_val <= 16'b0111101000011110;
            14'h339b 	:	o_val <= 16'b0111101000011111;
            14'h339c 	:	o_val <= 16'b0111101000100000;
            14'h339d 	:	o_val <= 16'b0111101000100001;
            14'h339e 	:	o_val <= 16'b0111101000100010;
            14'h339f 	:	o_val <= 16'b0111101000100011;
            14'h33a0 	:	o_val <= 16'b0111101000100100;
            14'h33a1 	:	o_val <= 16'b0111101000100101;
            14'h33a2 	:	o_val <= 16'b0111101000100110;
            14'h33a3 	:	o_val <= 16'b0111101000100111;
            14'h33a4 	:	o_val <= 16'b0111101000101000;
            14'h33a5 	:	o_val <= 16'b0111101000101001;
            14'h33a6 	:	o_val <= 16'b0111101000101010;
            14'h33a7 	:	o_val <= 16'b0111101000101011;
            14'h33a8 	:	o_val <= 16'b0111101000101100;
            14'h33a9 	:	o_val <= 16'b0111101000101101;
            14'h33aa 	:	o_val <= 16'b0111101000101101;
            14'h33ab 	:	o_val <= 16'b0111101000101110;
            14'h33ac 	:	o_val <= 16'b0111101000101111;
            14'h33ad 	:	o_val <= 16'b0111101000110000;
            14'h33ae 	:	o_val <= 16'b0111101000110001;
            14'h33af 	:	o_val <= 16'b0111101000110010;
            14'h33b0 	:	o_val <= 16'b0111101000110011;
            14'h33b1 	:	o_val <= 16'b0111101000110100;
            14'h33b2 	:	o_val <= 16'b0111101000110101;
            14'h33b3 	:	o_val <= 16'b0111101000110110;
            14'h33b4 	:	o_val <= 16'b0111101000110111;
            14'h33b5 	:	o_val <= 16'b0111101000111000;
            14'h33b6 	:	o_val <= 16'b0111101000111001;
            14'h33b7 	:	o_val <= 16'b0111101000111010;
            14'h33b8 	:	o_val <= 16'b0111101000111011;
            14'h33b9 	:	o_val <= 16'b0111101000111100;
            14'h33ba 	:	o_val <= 16'b0111101000111100;
            14'h33bb 	:	o_val <= 16'b0111101000111101;
            14'h33bc 	:	o_val <= 16'b0111101000111110;
            14'h33bd 	:	o_val <= 16'b0111101000111111;
            14'h33be 	:	o_val <= 16'b0111101001000000;
            14'h33bf 	:	o_val <= 16'b0111101001000001;
            14'h33c0 	:	o_val <= 16'b0111101001000010;
            14'h33c1 	:	o_val <= 16'b0111101001000011;
            14'h33c2 	:	o_val <= 16'b0111101001000100;
            14'h33c3 	:	o_val <= 16'b0111101001000101;
            14'h33c4 	:	o_val <= 16'b0111101001000110;
            14'h33c5 	:	o_val <= 16'b0111101001000111;
            14'h33c6 	:	o_val <= 16'b0111101001001000;
            14'h33c7 	:	o_val <= 16'b0111101001001001;
            14'h33c8 	:	o_val <= 16'b0111101001001001;
            14'h33c9 	:	o_val <= 16'b0111101001001010;
            14'h33ca 	:	o_val <= 16'b0111101001001011;
            14'h33cb 	:	o_val <= 16'b0111101001001100;
            14'h33cc 	:	o_val <= 16'b0111101001001101;
            14'h33cd 	:	o_val <= 16'b0111101001001110;
            14'h33ce 	:	o_val <= 16'b0111101001001111;
            14'h33cf 	:	o_val <= 16'b0111101001010000;
            14'h33d0 	:	o_val <= 16'b0111101001010001;
            14'h33d1 	:	o_val <= 16'b0111101001010010;
            14'h33d2 	:	o_val <= 16'b0111101001010011;
            14'h33d3 	:	o_val <= 16'b0111101001010100;
            14'h33d4 	:	o_val <= 16'b0111101001010101;
            14'h33d5 	:	o_val <= 16'b0111101001010110;
            14'h33d6 	:	o_val <= 16'b0111101001010110;
            14'h33d7 	:	o_val <= 16'b0111101001010111;
            14'h33d8 	:	o_val <= 16'b0111101001011000;
            14'h33d9 	:	o_val <= 16'b0111101001011001;
            14'h33da 	:	o_val <= 16'b0111101001011010;
            14'h33db 	:	o_val <= 16'b0111101001011011;
            14'h33dc 	:	o_val <= 16'b0111101001011100;
            14'h33dd 	:	o_val <= 16'b0111101001011101;
            14'h33de 	:	o_val <= 16'b0111101001011110;
            14'h33df 	:	o_val <= 16'b0111101001011111;
            14'h33e0 	:	o_val <= 16'b0111101001100000;
            14'h33e1 	:	o_val <= 16'b0111101001100001;
            14'h33e2 	:	o_val <= 16'b0111101001100001;
            14'h33e3 	:	o_val <= 16'b0111101001100010;
            14'h33e4 	:	o_val <= 16'b0111101001100011;
            14'h33e5 	:	o_val <= 16'b0111101001100100;
            14'h33e6 	:	o_val <= 16'b0111101001100101;
            14'h33e7 	:	o_val <= 16'b0111101001100110;
            14'h33e8 	:	o_val <= 16'b0111101001100111;
            14'h33e9 	:	o_val <= 16'b0111101001101000;
            14'h33ea 	:	o_val <= 16'b0111101001101001;
            14'h33eb 	:	o_val <= 16'b0111101001101010;
            14'h33ec 	:	o_val <= 16'b0111101001101011;
            14'h33ed 	:	o_val <= 16'b0111101001101100;
            14'h33ee 	:	o_val <= 16'b0111101001101101;
            14'h33ef 	:	o_val <= 16'b0111101001101101;
            14'h33f0 	:	o_val <= 16'b0111101001101110;
            14'h33f1 	:	o_val <= 16'b0111101001101111;
            14'h33f2 	:	o_val <= 16'b0111101001110000;
            14'h33f3 	:	o_val <= 16'b0111101001110001;
            14'h33f4 	:	o_val <= 16'b0111101001110010;
            14'h33f5 	:	o_val <= 16'b0111101001110011;
            14'h33f6 	:	o_val <= 16'b0111101001110100;
            14'h33f7 	:	o_val <= 16'b0111101001110101;
            14'h33f8 	:	o_val <= 16'b0111101001110110;
            14'h33f9 	:	o_val <= 16'b0111101001110111;
            14'h33fa 	:	o_val <= 16'b0111101001111000;
            14'h33fb 	:	o_val <= 16'b0111101001111000;
            14'h33fc 	:	o_val <= 16'b0111101001111001;
            14'h33fd 	:	o_val <= 16'b0111101001111010;
            14'h33fe 	:	o_val <= 16'b0111101001111011;
            14'h33ff 	:	o_val <= 16'b0111101001111100;
            14'h3400 	:	o_val <= 16'b0111101001111101;
            14'h3401 	:	o_val <= 16'b0111101001111110;
            14'h3402 	:	o_val <= 16'b0111101001111111;
            14'h3403 	:	o_val <= 16'b0111101010000000;
            14'h3404 	:	o_val <= 16'b0111101010000001;
            14'h3405 	:	o_val <= 16'b0111101010000010;
            14'h3406 	:	o_val <= 16'b0111101010000010;
            14'h3407 	:	o_val <= 16'b0111101010000011;
            14'h3408 	:	o_val <= 16'b0111101010000100;
            14'h3409 	:	o_val <= 16'b0111101010000101;
            14'h340a 	:	o_val <= 16'b0111101010000110;
            14'h340b 	:	o_val <= 16'b0111101010000111;
            14'h340c 	:	o_val <= 16'b0111101010001000;
            14'h340d 	:	o_val <= 16'b0111101010001001;
            14'h340e 	:	o_val <= 16'b0111101010001010;
            14'h340f 	:	o_val <= 16'b0111101010001011;
            14'h3410 	:	o_val <= 16'b0111101010001100;
            14'h3411 	:	o_val <= 16'b0111101010001100;
            14'h3412 	:	o_val <= 16'b0111101010001101;
            14'h3413 	:	o_val <= 16'b0111101010001110;
            14'h3414 	:	o_val <= 16'b0111101010001111;
            14'h3415 	:	o_val <= 16'b0111101010010000;
            14'h3416 	:	o_val <= 16'b0111101010010001;
            14'h3417 	:	o_val <= 16'b0111101010010010;
            14'h3418 	:	o_val <= 16'b0111101010010011;
            14'h3419 	:	o_val <= 16'b0111101010010100;
            14'h341a 	:	o_val <= 16'b0111101010010101;
            14'h341b 	:	o_val <= 16'b0111101010010101;
            14'h341c 	:	o_val <= 16'b0111101010010110;
            14'h341d 	:	o_val <= 16'b0111101010010111;
            14'h341e 	:	o_val <= 16'b0111101010011000;
            14'h341f 	:	o_val <= 16'b0111101010011001;
            14'h3420 	:	o_val <= 16'b0111101010011010;
            14'h3421 	:	o_val <= 16'b0111101010011011;
            14'h3422 	:	o_val <= 16'b0111101010011100;
            14'h3423 	:	o_val <= 16'b0111101010011101;
            14'h3424 	:	o_val <= 16'b0111101010011110;
            14'h3425 	:	o_val <= 16'b0111101010011111;
            14'h3426 	:	o_val <= 16'b0111101010011111;
            14'h3427 	:	o_val <= 16'b0111101010100000;
            14'h3428 	:	o_val <= 16'b0111101010100001;
            14'h3429 	:	o_val <= 16'b0111101010100010;
            14'h342a 	:	o_val <= 16'b0111101010100011;
            14'h342b 	:	o_val <= 16'b0111101010100100;
            14'h342c 	:	o_val <= 16'b0111101010100101;
            14'h342d 	:	o_val <= 16'b0111101010100110;
            14'h342e 	:	o_val <= 16'b0111101010100111;
            14'h342f 	:	o_val <= 16'b0111101010101000;
            14'h3430 	:	o_val <= 16'b0111101010101000;
            14'h3431 	:	o_val <= 16'b0111101010101001;
            14'h3432 	:	o_val <= 16'b0111101010101010;
            14'h3433 	:	o_val <= 16'b0111101010101011;
            14'h3434 	:	o_val <= 16'b0111101010101100;
            14'h3435 	:	o_val <= 16'b0111101010101101;
            14'h3436 	:	o_val <= 16'b0111101010101110;
            14'h3437 	:	o_val <= 16'b0111101010101111;
            14'h3438 	:	o_val <= 16'b0111101010110000;
            14'h3439 	:	o_val <= 16'b0111101010110000;
            14'h343a 	:	o_val <= 16'b0111101010110001;
            14'h343b 	:	o_val <= 16'b0111101010110010;
            14'h343c 	:	o_val <= 16'b0111101010110011;
            14'h343d 	:	o_val <= 16'b0111101010110100;
            14'h343e 	:	o_val <= 16'b0111101010110101;
            14'h343f 	:	o_val <= 16'b0111101010110110;
            14'h3440 	:	o_val <= 16'b0111101010110111;
            14'h3441 	:	o_val <= 16'b0111101010111000;
            14'h3442 	:	o_val <= 16'b0111101010111001;
            14'h3443 	:	o_val <= 16'b0111101010111001;
            14'h3444 	:	o_val <= 16'b0111101010111010;
            14'h3445 	:	o_val <= 16'b0111101010111011;
            14'h3446 	:	o_val <= 16'b0111101010111100;
            14'h3447 	:	o_val <= 16'b0111101010111101;
            14'h3448 	:	o_val <= 16'b0111101010111110;
            14'h3449 	:	o_val <= 16'b0111101010111111;
            14'h344a 	:	o_val <= 16'b0111101011000000;
            14'h344b 	:	o_val <= 16'b0111101011000001;
            14'h344c 	:	o_val <= 16'b0111101011000001;
            14'h344d 	:	o_val <= 16'b0111101011000010;
            14'h344e 	:	o_val <= 16'b0111101011000011;
            14'h344f 	:	o_val <= 16'b0111101011000100;
            14'h3450 	:	o_val <= 16'b0111101011000101;
            14'h3451 	:	o_val <= 16'b0111101011000110;
            14'h3452 	:	o_val <= 16'b0111101011000111;
            14'h3453 	:	o_val <= 16'b0111101011001000;
            14'h3454 	:	o_val <= 16'b0111101011001001;
            14'h3455 	:	o_val <= 16'b0111101011001001;
            14'h3456 	:	o_val <= 16'b0111101011001010;
            14'h3457 	:	o_val <= 16'b0111101011001011;
            14'h3458 	:	o_val <= 16'b0111101011001100;
            14'h3459 	:	o_val <= 16'b0111101011001101;
            14'h345a 	:	o_val <= 16'b0111101011001110;
            14'h345b 	:	o_val <= 16'b0111101011001111;
            14'h345c 	:	o_val <= 16'b0111101011010000;
            14'h345d 	:	o_val <= 16'b0111101011010001;
            14'h345e 	:	o_val <= 16'b0111101011010001;
            14'h345f 	:	o_val <= 16'b0111101011010010;
            14'h3460 	:	o_val <= 16'b0111101011010011;
            14'h3461 	:	o_val <= 16'b0111101011010100;
            14'h3462 	:	o_val <= 16'b0111101011010101;
            14'h3463 	:	o_val <= 16'b0111101011010110;
            14'h3464 	:	o_val <= 16'b0111101011010111;
            14'h3465 	:	o_val <= 16'b0111101011011000;
            14'h3466 	:	o_val <= 16'b0111101011011000;
            14'h3467 	:	o_val <= 16'b0111101011011001;
            14'h3468 	:	o_val <= 16'b0111101011011010;
            14'h3469 	:	o_val <= 16'b0111101011011011;
            14'h346a 	:	o_val <= 16'b0111101011011100;
            14'h346b 	:	o_val <= 16'b0111101011011101;
            14'h346c 	:	o_val <= 16'b0111101011011110;
            14'h346d 	:	o_val <= 16'b0111101011011111;
            14'h346e 	:	o_val <= 16'b0111101011100000;
            14'h346f 	:	o_val <= 16'b0111101011100000;
            14'h3470 	:	o_val <= 16'b0111101011100001;
            14'h3471 	:	o_val <= 16'b0111101011100010;
            14'h3472 	:	o_val <= 16'b0111101011100011;
            14'h3473 	:	o_val <= 16'b0111101011100100;
            14'h3474 	:	o_val <= 16'b0111101011100101;
            14'h3475 	:	o_val <= 16'b0111101011100110;
            14'h3476 	:	o_val <= 16'b0111101011100111;
            14'h3477 	:	o_val <= 16'b0111101011100111;
            14'h3478 	:	o_val <= 16'b0111101011101000;
            14'h3479 	:	o_val <= 16'b0111101011101001;
            14'h347a 	:	o_val <= 16'b0111101011101010;
            14'h347b 	:	o_val <= 16'b0111101011101011;
            14'h347c 	:	o_val <= 16'b0111101011101100;
            14'h347d 	:	o_val <= 16'b0111101011101101;
            14'h347e 	:	o_val <= 16'b0111101011101110;
            14'h347f 	:	o_val <= 16'b0111101011101110;
            14'h3480 	:	o_val <= 16'b0111101011101111;
            14'h3481 	:	o_val <= 16'b0111101011110000;
            14'h3482 	:	o_val <= 16'b0111101011110001;
            14'h3483 	:	o_val <= 16'b0111101011110010;
            14'h3484 	:	o_val <= 16'b0111101011110011;
            14'h3485 	:	o_val <= 16'b0111101011110100;
            14'h3486 	:	o_val <= 16'b0111101011110101;
            14'h3487 	:	o_val <= 16'b0111101011110101;
            14'h3488 	:	o_val <= 16'b0111101011110110;
            14'h3489 	:	o_val <= 16'b0111101011110111;
            14'h348a 	:	o_val <= 16'b0111101011111000;
            14'h348b 	:	o_val <= 16'b0111101011111001;
            14'h348c 	:	o_val <= 16'b0111101011111010;
            14'h348d 	:	o_val <= 16'b0111101011111011;
            14'h348e 	:	o_val <= 16'b0111101011111100;
            14'h348f 	:	o_val <= 16'b0111101011111100;
            14'h3490 	:	o_val <= 16'b0111101011111101;
            14'h3491 	:	o_val <= 16'b0111101011111110;
            14'h3492 	:	o_val <= 16'b0111101011111111;
            14'h3493 	:	o_val <= 16'b0111101100000000;
            14'h3494 	:	o_val <= 16'b0111101100000001;
            14'h3495 	:	o_val <= 16'b0111101100000010;
            14'h3496 	:	o_val <= 16'b0111101100000011;
            14'h3497 	:	o_val <= 16'b0111101100000011;
            14'h3498 	:	o_val <= 16'b0111101100000100;
            14'h3499 	:	o_val <= 16'b0111101100000101;
            14'h349a 	:	o_val <= 16'b0111101100000110;
            14'h349b 	:	o_val <= 16'b0111101100000111;
            14'h349c 	:	o_val <= 16'b0111101100001000;
            14'h349d 	:	o_val <= 16'b0111101100001001;
            14'h349e 	:	o_val <= 16'b0111101100001001;
            14'h349f 	:	o_val <= 16'b0111101100001010;
            14'h34a0 	:	o_val <= 16'b0111101100001011;
            14'h34a1 	:	o_val <= 16'b0111101100001100;
            14'h34a2 	:	o_val <= 16'b0111101100001101;
            14'h34a3 	:	o_val <= 16'b0111101100001110;
            14'h34a4 	:	o_val <= 16'b0111101100001111;
            14'h34a5 	:	o_val <= 16'b0111101100001111;
            14'h34a6 	:	o_val <= 16'b0111101100010000;
            14'h34a7 	:	o_val <= 16'b0111101100010001;
            14'h34a8 	:	o_val <= 16'b0111101100010010;
            14'h34a9 	:	o_val <= 16'b0111101100010011;
            14'h34aa 	:	o_val <= 16'b0111101100010100;
            14'h34ab 	:	o_val <= 16'b0111101100010101;
            14'h34ac 	:	o_val <= 16'b0111101100010110;
            14'h34ad 	:	o_val <= 16'b0111101100010110;
            14'h34ae 	:	o_val <= 16'b0111101100010111;
            14'h34af 	:	o_val <= 16'b0111101100011000;
            14'h34b0 	:	o_val <= 16'b0111101100011001;
            14'h34b1 	:	o_val <= 16'b0111101100011010;
            14'h34b2 	:	o_val <= 16'b0111101100011011;
            14'h34b3 	:	o_val <= 16'b0111101100011100;
            14'h34b4 	:	o_val <= 16'b0111101100011100;
            14'h34b5 	:	o_val <= 16'b0111101100011101;
            14'h34b6 	:	o_val <= 16'b0111101100011110;
            14'h34b7 	:	o_val <= 16'b0111101100011111;
            14'h34b8 	:	o_val <= 16'b0111101100100000;
            14'h34b9 	:	o_val <= 16'b0111101100100001;
            14'h34ba 	:	o_val <= 16'b0111101100100010;
            14'h34bb 	:	o_val <= 16'b0111101100100010;
            14'h34bc 	:	o_val <= 16'b0111101100100011;
            14'h34bd 	:	o_val <= 16'b0111101100100100;
            14'h34be 	:	o_val <= 16'b0111101100100101;
            14'h34bf 	:	o_val <= 16'b0111101100100110;
            14'h34c0 	:	o_val <= 16'b0111101100100111;
            14'h34c1 	:	o_val <= 16'b0111101100101000;
            14'h34c2 	:	o_val <= 16'b0111101100101000;
            14'h34c3 	:	o_val <= 16'b0111101100101001;
            14'h34c4 	:	o_val <= 16'b0111101100101010;
            14'h34c5 	:	o_val <= 16'b0111101100101011;
            14'h34c6 	:	o_val <= 16'b0111101100101100;
            14'h34c7 	:	o_val <= 16'b0111101100101101;
            14'h34c8 	:	o_val <= 16'b0111101100101110;
            14'h34c9 	:	o_val <= 16'b0111101100101110;
            14'h34ca 	:	o_val <= 16'b0111101100101111;
            14'h34cb 	:	o_val <= 16'b0111101100110000;
            14'h34cc 	:	o_val <= 16'b0111101100110001;
            14'h34cd 	:	o_val <= 16'b0111101100110010;
            14'h34ce 	:	o_val <= 16'b0111101100110011;
            14'h34cf 	:	o_val <= 16'b0111101100110100;
            14'h34d0 	:	o_val <= 16'b0111101100110100;
            14'h34d1 	:	o_val <= 16'b0111101100110101;
            14'h34d2 	:	o_val <= 16'b0111101100110110;
            14'h34d3 	:	o_val <= 16'b0111101100110111;
            14'h34d4 	:	o_val <= 16'b0111101100111000;
            14'h34d5 	:	o_val <= 16'b0111101100111001;
            14'h34d6 	:	o_val <= 16'b0111101100111001;
            14'h34d7 	:	o_val <= 16'b0111101100111010;
            14'h34d8 	:	o_val <= 16'b0111101100111011;
            14'h34d9 	:	o_val <= 16'b0111101100111100;
            14'h34da 	:	o_val <= 16'b0111101100111101;
            14'h34db 	:	o_val <= 16'b0111101100111110;
            14'h34dc 	:	o_val <= 16'b0111101100111111;
            14'h34dd 	:	o_val <= 16'b0111101100111111;
            14'h34de 	:	o_val <= 16'b0111101101000000;
            14'h34df 	:	o_val <= 16'b0111101101000001;
            14'h34e0 	:	o_val <= 16'b0111101101000010;
            14'h34e1 	:	o_val <= 16'b0111101101000011;
            14'h34e2 	:	o_val <= 16'b0111101101000100;
            14'h34e3 	:	o_val <= 16'b0111101101000101;
            14'h34e4 	:	o_val <= 16'b0111101101000101;
            14'h34e5 	:	o_val <= 16'b0111101101000110;
            14'h34e6 	:	o_val <= 16'b0111101101000111;
            14'h34e7 	:	o_val <= 16'b0111101101001000;
            14'h34e8 	:	o_val <= 16'b0111101101001001;
            14'h34e9 	:	o_val <= 16'b0111101101001010;
            14'h34ea 	:	o_val <= 16'b0111101101001010;
            14'h34eb 	:	o_val <= 16'b0111101101001011;
            14'h34ec 	:	o_val <= 16'b0111101101001100;
            14'h34ed 	:	o_val <= 16'b0111101101001101;
            14'h34ee 	:	o_val <= 16'b0111101101001110;
            14'h34ef 	:	o_val <= 16'b0111101101001111;
            14'h34f0 	:	o_val <= 16'b0111101101001111;
            14'h34f1 	:	o_val <= 16'b0111101101010000;
            14'h34f2 	:	o_val <= 16'b0111101101010001;
            14'h34f3 	:	o_val <= 16'b0111101101010010;
            14'h34f4 	:	o_val <= 16'b0111101101010011;
            14'h34f5 	:	o_val <= 16'b0111101101010100;
            14'h34f6 	:	o_val <= 16'b0111101101010101;
            14'h34f7 	:	o_val <= 16'b0111101101010101;
            14'h34f8 	:	o_val <= 16'b0111101101010110;
            14'h34f9 	:	o_val <= 16'b0111101101010111;
            14'h34fa 	:	o_val <= 16'b0111101101011000;
            14'h34fb 	:	o_val <= 16'b0111101101011001;
            14'h34fc 	:	o_val <= 16'b0111101101011010;
            14'h34fd 	:	o_val <= 16'b0111101101011010;
            14'h34fe 	:	o_val <= 16'b0111101101011011;
            14'h34ff 	:	o_val <= 16'b0111101101011100;
            14'h3500 	:	o_val <= 16'b0111101101011101;
            14'h3501 	:	o_val <= 16'b0111101101011110;
            14'h3502 	:	o_val <= 16'b0111101101011111;
            14'h3503 	:	o_val <= 16'b0111101101011111;
            14'h3504 	:	o_val <= 16'b0111101101100000;
            14'h3505 	:	o_val <= 16'b0111101101100001;
            14'h3506 	:	o_val <= 16'b0111101101100010;
            14'h3507 	:	o_val <= 16'b0111101101100011;
            14'h3508 	:	o_val <= 16'b0111101101100100;
            14'h3509 	:	o_val <= 16'b0111101101100100;
            14'h350a 	:	o_val <= 16'b0111101101100101;
            14'h350b 	:	o_val <= 16'b0111101101100110;
            14'h350c 	:	o_val <= 16'b0111101101100111;
            14'h350d 	:	o_val <= 16'b0111101101101000;
            14'h350e 	:	o_val <= 16'b0111101101101001;
            14'h350f 	:	o_val <= 16'b0111101101101001;
            14'h3510 	:	o_val <= 16'b0111101101101010;
            14'h3511 	:	o_val <= 16'b0111101101101011;
            14'h3512 	:	o_val <= 16'b0111101101101100;
            14'h3513 	:	o_val <= 16'b0111101101101101;
            14'h3514 	:	o_val <= 16'b0111101101101110;
            14'h3515 	:	o_val <= 16'b0111101101101110;
            14'h3516 	:	o_val <= 16'b0111101101101111;
            14'h3517 	:	o_val <= 16'b0111101101110000;
            14'h3518 	:	o_val <= 16'b0111101101110001;
            14'h3519 	:	o_val <= 16'b0111101101110010;
            14'h351a 	:	o_val <= 16'b0111101101110011;
            14'h351b 	:	o_val <= 16'b0111101101110011;
            14'h351c 	:	o_val <= 16'b0111101101110100;
            14'h351d 	:	o_val <= 16'b0111101101110101;
            14'h351e 	:	o_val <= 16'b0111101101110110;
            14'h351f 	:	o_val <= 16'b0111101101110111;
            14'h3520 	:	o_val <= 16'b0111101101111000;
            14'h3521 	:	o_val <= 16'b0111101101111000;
            14'h3522 	:	o_val <= 16'b0111101101111001;
            14'h3523 	:	o_val <= 16'b0111101101111010;
            14'h3524 	:	o_val <= 16'b0111101101111011;
            14'h3525 	:	o_val <= 16'b0111101101111100;
            14'h3526 	:	o_val <= 16'b0111101101111101;
            14'h3527 	:	o_val <= 16'b0111101101111101;
            14'h3528 	:	o_val <= 16'b0111101101111110;
            14'h3529 	:	o_val <= 16'b0111101101111111;
            14'h352a 	:	o_val <= 16'b0111101110000000;
            14'h352b 	:	o_val <= 16'b0111101110000001;
            14'h352c 	:	o_val <= 16'b0111101110000010;
            14'h352d 	:	o_val <= 16'b0111101110000010;
            14'h352e 	:	o_val <= 16'b0111101110000011;
            14'h352f 	:	o_val <= 16'b0111101110000100;
            14'h3530 	:	o_val <= 16'b0111101110000101;
            14'h3531 	:	o_val <= 16'b0111101110000110;
            14'h3532 	:	o_val <= 16'b0111101110000110;
            14'h3533 	:	o_val <= 16'b0111101110000111;
            14'h3534 	:	o_val <= 16'b0111101110001000;
            14'h3535 	:	o_val <= 16'b0111101110001001;
            14'h3536 	:	o_val <= 16'b0111101110001010;
            14'h3537 	:	o_val <= 16'b0111101110001011;
            14'h3538 	:	o_val <= 16'b0111101110001011;
            14'h3539 	:	o_val <= 16'b0111101110001100;
            14'h353a 	:	o_val <= 16'b0111101110001101;
            14'h353b 	:	o_val <= 16'b0111101110001110;
            14'h353c 	:	o_val <= 16'b0111101110001111;
            14'h353d 	:	o_val <= 16'b0111101110001111;
            14'h353e 	:	o_val <= 16'b0111101110010000;
            14'h353f 	:	o_val <= 16'b0111101110010001;
            14'h3540 	:	o_val <= 16'b0111101110010010;
            14'h3541 	:	o_val <= 16'b0111101110010011;
            14'h3542 	:	o_val <= 16'b0111101110010100;
            14'h3543 	:	o_val <= 16'b0111101110010100;
            14'h3544 	:	o_val <= 16'b0111101110010101;
            14'h3545 	:	o_val <= 16'b0111101110010110;
            14'h3546 	:	o_val <= 16'b0111101110010111;
            14'h3547 	:	o_val <= 16'b0111101110011000;
            14'h3548 	:	o_val <= 16'b0111101110011000;
            14'h3549 	:	o_val <= 16'b0111101110011001;
            14'h354a 	:	o_val <= 16'b0111101110011010;
            14'h354b 	:	o_val <= 16'b0111101110011011;
            14'h354c 	:	o_val <= 16'b0111101110011100;
            14'h354d 	:	o_val <= 16'b0111101110011101;
            14'h354e 	:	o_val <= 16'b0111101110011101;
            14'h354f 	:	o_val <= 16'b0111101110011110;
            14'h3550 	:	o_val <= 16'b0111101110011111;
            14'h3551 	:	o_val <= 16'b0111101110100000;
            14'h3552 	:	o_val <= 16'b0111101110100001;
            14'h3553 	:	o_val <= 16'b0111101110100001;
            14'h3554 	:	o_val <= 16'b0111101110100010;
            14'h3555 	:	o_val <= 16'b0111101110100011;
            14'h3556 	:	o_val <= 16'b0111101110100100;
            14'h3557 	:	o_val <= 16'b0111101110100101;
            14'h3558 	:	o_val <= 16'b0111101110100110;
            14'h3559 	:	o_val <= 16'b0111101110100110;
            14'h355a 	:	o_val <= 16'b0111101110100111;
            14'h355b 	:	o_val <= 16'b0111101110101000;
            14'h355c 	:	o_val <= 16'b0111101110101001;
            14'h355d 	:	o_val <= 16'b0111101110101010;
            14'h355e 	:	o_val <= 16'b0111101110101010;
            14'h355f 	:	o_val <= 16'b0111101110101011;
            14'h3560 	:	o_val <= 16'b0111101110101100;
            14'h3561 	:	o_val <= 16'b0111101110101101;
            14'h3562 	:	o_val <= 16'b0111101110101110;
            14'h3563 	:	o_val <= 16'b0111101110101110;
            14'h3564 	:	o_val <= 16'b0111101110101111;
            14'h3565 	:	o_val <= 16'b0111101110110000;
            14'h3566 	:	o_val <= 16'b0111101110110001;
            14'h3567 	:	o_val <= 16'b0111101110110010;
            14'h3568 	:	o_val <= 16'b0111101110110010;
            14'h3569 	:	o_val <= 16'b0111101110110011;
            14'h356a 	:	o_val <= 16'b0111101110110100;
            14'h356b 	:	o_val <= 16'b0111101110110101;
            14'h356c 	:	o_val <= 16'b0111101110110110;
            14'h356d 	:	o_val <= 16'b0111101110110111;
            14'h356e 	:	o_val <= 16'b0111101110110111;
            14'h356f 	:	o_val <= 16'b0111101110111000;
            14'h3570 	:	o_val <= 16'b0111101110111001;
            14'h3571 	:	o_val <= 16'b0111101110111010;
            14'h3572 	:	o_val <= 16'b0111101110111011;
            14'h3573 	:	o_val <= 16'b0111101110111011;
            14'h3574 	:	o_val <= 16'b0111101110111100;
            14'h3575 	:	o_val <= 16'b0111101110111101;
            14'h3576 	:	o_val <= 16'b0111101110111110;
            14'h3577 	:	o_val <= 16'b0111101110111111;
            14'h3578 	:	o_val <= 16'b0111101110111111;
            14'h3579 	:	o_val <= 16'b0111101111000000;
            14'h357a 	:	o_val <= 16'b0111101111000001;
            14'h357b 	:	o_val <= 16'b0111101111000010;
            14'h357c 	:	o_val <= 16'b0111101111000011;
            14'h357d 	:	o_val <= 16'b0111101111000011;
            14'h357e 	:	o_val <= 16'b0111101111000100;
            14'h357f 	:	o_val <= 16'b0111101111000101;
            14'h3580 	:	o_val <= 16'b0111101111000110;
            14'h3581 	:	o_val <= 16'b0111101111000111;
            14'h3582 	:	o_val <= 16'b0111101111000111;
            14'h3583 	:	o_val <= 16'b0111101111001000;
            14'h3584 	:	o_val <= 16'b0111101111001001;
            14'h3585 	:	o_val <= 16'b0111101111001010;
            14'h3586 	:	o_val <= 16'b0111101111001011;
            14'h3587 	:	o_val <= 16'b0111101111001011;
            14'h3588 	:	o_val <= 16'b0111101111001100;
            14'h3589 	:	o_val <= 16'b0111101111001101;
            14'h358a 	:	o_val <= 16'b0111101111001110;
            14'h358b 	:	o_val <= 16'b0111101111001111;
            14'h358c 	:	o_val <= 16'b0111101111001111;
            14'h358d 	:	o_val <= 16'b0111101111010000;
            14'h358e 	:	o_val <= 16'b0111101111010001;
            14'h358f 	:	o_val <= 16'b0111101111010010;
            14'h3590 	:	o_val <= 16'b0111101111010011;
            14'h3591 	:	o_val <= 16'b0111101111010011;
            14'h3592 	:	o_val <= 16'b0111101111010100;
            14'h3593 	:	o_val <= 16'b0111101111010101;
            14'h3594 	:	o_val <= 16'b0111101111010110;
            14'h3595 	:	o_val <= 16'b0111101111010111;
            14'h3596 	:	o_val <= 16'b0111101111010111;
            14'h3597 	:	o_val <= 16'b0111101111011000;
            14'h3598 	:	o_val <= 16'b0111101111011001;
            14'h3599 	:	o_val <= 16'b0111101111011010;
            14'h359a 	:	o_val <= 16'b0111101111011011;
            14'h359b 	:	o_val <= 16'b0111101111011011;
            14'h359c 	:	o_val <= 16'b0111101111011100;
            14'h359d 	:	o_val <= 16'b0111101111011101;
            14'h359e 	:	o_val <= 16'b0111101111011110;
            14'h359f 	:	o_val <= 16'b0111101111011110;
            14'h35a0 	:	o_val <= 16'b0111101111011111;
            14'h35a1 	:	o_val <= 16'b0111101111100000;
            14'h35a2 	:	o_val <= 16'b0111101111100001;
            14'h35a3 	:	o_val <= 16'b0111101111100010;
            14'h35a4 	:	o_val <= 16'b0111101111100010;
            14'h35a5 	:	o_val <= 16'b0111101111100011;
            14'h35a6 	:	o_val <= 16'b0111101111100100;
            14'h35a7 	:	o_val <= 16'b0111101111100101;
            14'h35a8 	:	o_val <= 16'b0111101111100110;
            14'h35a9 	:	o_val <= 16'b0111101111100110;
            14'h35aa 	:	o_val <= 16'b0111101111100111;
            14'h35ab 	:	o_val <= 16'b0111101111101000;
            14'h35ac 	:	o_val <= 16'b0111101111101001;
            14'h35ad 	:	o_val <= 16'b0111101111101010;
            14'h35ae 	:	o_val <= 16'b0111101111101010;
            14'h35af 	:	o_val <= 16'b0111101111101011;
            14'h35b0 	:	o_val <= 16'b0111101111101100;
            14'h35b1 	:	o_val <= 16'b0111101111101101;
            14'h35b2 	:	o_val <= 16'b0111101111101101;
            14'h35b3 	:	o_val <= 16'b0111101111101110;
            14'h35b4 	:	o_val <= 16'b0111101111101111;
            14'h35b5 	:	o_val <= 16'b0111101111110000;
            14'h35b6 	:	o_val <= 16'b0111101111110001;
            14'h35b7 	:	o_val <= 16'b0111101111110001;
            14'h35b8 	:	o_val <= 16'b0111101111110010;
            14'h35b9 	:	o_val <= 16'b0111101111110011;
            14'h35ba 	:	o_val <= 16'b0111101111110100;
            14'h35bb 	:	o_val <= 16'b0111101111110101;
            14'h35bc 	:	o_val <= 16'b0111101111110101;
            14'h35bd 	:	o_val <= 16'b0111101111110110;
            14'h35be 	:	o_val <= 16'b0111101111110111;
            14'h35bf 	:	o_val <= 16'b0111101111111000;
            14'h35c0 	:	o_val <= 16'b0111101111111000;
            14'h35c1 	:	o_val <= 16'b0111101111111001;
            14'h35c2 	:	o_val <= 16'b0111101111111010;
            14'h35c3 	:	o_val <= 16'b0111101111111011;
            14'h35c4 	:	o_val <= 16'b0111101111111100;
            14'h35c5 	:	o_val <= 16'b0111101111111100;
            14'h35c6 	:	o_val <= 16'b0111101111111101;
            14'h35c7 	:	o_val <= 16'b0111101111111110;
            14'h35c8 	:	o_val <= 16'b0111101111111111;
            14'h35c9 	:	o_val <= 16'b0111101111111111;
            14'h35ca 	:	o_val <= 16'b0111110000000000;
            14'h35cb 	:	o_val <= 16'b0111110000000001;
            14'h35cc 	:	o_val <= 16'b0111110000000010;
            14'h35cd 	:	o_val <= 16'b0111110000000011;
            14'h35ce 	:	o_val <= 16'b0111110000000011;
            14'h35cf 	:	o_val <= 16'b0111110000000100;
            14'h35d0 	:	o_val <= 16'b0111110000000101;
            14'h35d1 	:	o_val <= 16'b0111110000000110;
            14'h35d2 	:	o_val <= 16'b0111110000000110;
            14'h35d3 	:	o_val <= 16'b0111110000000111;
            14'h35d4 	:	o_val <= 16'b0111110000001000;
            14'h35d5 	:	o_val <= 16'b0111110000001001;
            14'h35d6 	:	o_val <= 16'b0111110000001010;
            14'h35d7 	:	o_val <= 16'b0111110000001010;
            14'h35d8 	:	o_val <= 16'b0111110000001011;
            14'h35d9 	:	o_val <= 16'b0111110000001100;
            14'h35da 	:	o_val <= 16'b0111110000001101;
            14'h35db 	:	o_val <= 16'b0111110000001101;
            14'h35dc 	:	o_val <= 16'b0111110000001110;
            14'h35dd 	:	o_val <= 16'b0111110000001111;
            14'h35de 	:	o_val <= 16'b0111110000010000;
            14'h35df 	:	o_val <= 16'b0111110000010001;
            14'h35e0 	:	o_val <= 16'b0111110000010001;
            14'h35e1 	:	o_val <= 16'b0111110000010010;
            14'h35e2 	:	o_val <= 16'b0111110000010011;
            14'h35e3 	:	o_val <= 16'b0111110000010100;
            14'h35e4 	:	o_val <= 16'b0111110000010100;
            14'h35e5 	:	o_val <= 16'b0111110000010101;
            14'h35e6 	:	o_val <= 16'b0111110000010110;
            14'h35e7 	:	o_val <= 16'b0111110000010111;
            14'h35e8 	:	o_val <= 16'b0111110000010111;
            14'h35e9 	:	o_val <= 16'b0111110000011000;
            14'h35ea 	:	o_val <= 16'b0111110000011001;
            14'h35eb 	:	o_val <= 16'b0111110000011010;
            14'h35ec 	:	o_val <= 16'b0111110000011011;
            14'h35ed 	:	o_val <= 16'b0111110000011011;
            14'h35ee 	:	o_val <= 16'b0111110000011100;
            14'h35ef 	:	o_val <= 16'b0111110000011101;
            14'h35f0 	:	o_val <= 16'b0111110000011110;
            14'h35f1 	:	o_val <= 16'b0111110000011110;
            14'h35f2 	:	o_val <= 16'b0111110000011111;
            14'h35f3 	:	o_val <= 16'b0111110000100000;
            14'h35f4 	:	o_val <= 16'b0111110000100001;
            14'h35f5 	:	o_val <= 16'b0111110000100001;
            14'h35f6 	:	o_val <= 16'b0111110000100010;
            14'h35f7 	:	o_val <= 16'b0111110000100011;
            14'h35f8 	:	o_val <= 16'b0111110000100100;
            14'h35f9 	:	o_val <= 16'b0111110000100101;
            14'h35fa 	:	o_val <= 16'b0111110000100101;
            14'h35fb 	:	o_val <= 16'b0111110000100110;
            14'h35fc 	:	o_val <= 16'b0111110000100111;
            14'h35fd 	:	o_val <= 16'b0111110000101000;
            14'h35fe 	:	o_val <= 16'b0111110000101000;
            14'h35ff 	:	o_val <= 16'b0111110000101001;
            14'h3600 	:	o_val <= 16'b0111110000101010;
            14'h3601 	:	o_val <= 16'b0111110000101011;
            14'h3602 	:	o_val <= 16'b0111110000101011;
            14'h3603 	:	o_val <= 16'b0111110000101100;
            14'h3604 	:	o_val <= 16'b0111110000101101;
            14'h3605 	:	o_val <= 16'b0111110000101110;
            14'h3606 	:	o_val <= 16'b0111110000101110;
            14'h3607 	:	o_val <= 16'b0111110000101111;
            14'h3608 	:	o_val <= 16'b0111110000110000;
            14'h3609 	:	o_val <= 16'b0111110000110001;
            14'h360a 	:	o_val <= 16'b0111110000110001;
            14'h360b 	:	o_val <= 16'b0111110000110010;
            14'h360c 	:	o_val <= 16'b0111110000110011;
            14'h360d 	:	o_val <= 16'b0111110000110100;
            14'h360e 	:	o_val <= 16'b0111110000110101;
            14'h360f 	:	o_val <= 16'b0111110000110101;
            14'h3610 	:	o_val <= 16'b0111110000110110;
            14'h3611 	:	o_val <= 16'b0111110000110111;
            14'h3612 	:	o_val <= 16'b0111110000111000;
            14'h3613 	:	o_val <= 16'b0111110000111000;
            14'h3614 	:	o_val <= 16'b0111110000111001;
            14'h3615 	:	o_val <= 16'b0111110000111010;
            14'h3616 	:	o_val <= 16'b0111110000111011;
            14'h3617 	:	o_val <= 16'b0111110000111011;
            14'h3618 	:	o_val <= 16'b0111110000111100;
            14'h3619 	:	o_val <= 16'b0111110000111101;
            14'h361a 	:	o_val <= 16'b0111110000111110;
            14'h361b 	:	o_val <= 16'b0111110000111110;
            14'h361c 	:	o_val <= 16'b0111110000111111;
            14'h361d 	:	o_val <= 16'b0111110001000000;
            14'h361e 	:	o_val <= 16'b0111110001000001;
            14'h361f 	:	o_val <= 16'b0111110001000001;
            14'h3620 	:	o_val <= 16'b0111110001000010;
            14'h3621 	:	o_val <= 16'b0111110001000011;
            14'h3622 	:	o_val <= 16'b0111110001000100;
            14'h3623 	:	o_val <= 16'b0111110001000100;
            14'h3624 	:	o_val <= 16'b0111110001000101;
            14'h3625 	:	o_val <= 16'b0111110001000110;
            14'h3626 	:	o_val <= 16'b0111110001000111;
            14'h3627 	:	o_val <= 16'b0111110001000111;
            14'h3628 	:	o_val <= 16'b0111110001001000;
            14'h3629 	:	o_val <= 16'b0111110001001001;
            14'h362a 	:	o_val <= 16'b0111110001001010;
            14'h362b 	:	o_val <= 16'b0111110001001010;
            14'h362c 	:	o_val <= 16'b0111110001001011;
            14'h362d 	:	o_val <= 16'b0111110001001100;
            14'h362e 	:	o_val <= 16'b0111110001001101;
            14'h362f 	:	o_val <= 16'b0111110001001101;
            14'h3630 	:	o_val <= 16'b0111110001001110;
            14'h3631 	:	o_val <= 16'b0111110001001111;
            14'h3632 	:	o_val <= 16'b0111110001010000;
            14'h3633 	:	o_val <= 16'b0111110001010000;
            14'h3634 	:	o_val <= 16'b0111110001010001;
            14'h3635 	:	o_val <= 16'b0111110001010010;
            14'h3636 	:	o_val <= 16'b0111110001010011;
            14'h3637 	:	o_val <= 16'b0111110001010011;
            14'h3638 	:	o_val <= 16'b0111110001010100;
            14'h3639 	:	o_val <= 16'b0111110001010101;
            14'h363a 	:	o_val <= 16'b0111110001010110;
            14'h363b 	:	o_val <= 16'b0111110001010110;
            14'h363c 	:	o_val <= 16'b0111110001010111;
            14'h363d 	:	o_val <= 16'b0111110001011000;
            14'h363e 	:	o_val <= 16'b0111110001011001;
            14'h363f 	:	o_val <= 16'b0111110001011001;
            14'h3640 	:	o_val <= 16'b0111110001011010;
            14'h3641 	:	o_val <= 16'b0111110001011011;
            14'h3642 	:	o_val <= 16'b0111110001011100;
            14'h3643 	:	o_val <= 16'b0111110001011100;
            14'h3644 	:	o_val <= 16'b0111110001011101;
            14'h3645 	:	o_val <= 16'b0111110001011110;
            14'h3646 	:	o_val <= 16'b0111110001011111;
            14'h3647 	:	o_val <= 16'b0111110001011111;
            14'h3648 	:	o_val <= 16'b0111110001100000;
            14'h3649 	:	o_val <= 16'b0111110001100001;
            14'h364a 	:	o_val <= 16'b0111110001100010;
            14'h364b 	:	o_val <= 16'b0111110001100010;
            14'h364c 	:	o_val <= 16'b0111110001100011;
            14'h364d 	:	o_val <= 16'b0111110001100100;
            14'h364e 	:	o_val <= 16'b0111110001100101;
            14'h364f 	:	o_val <= 16'b0111110001100101;
            14'h3650 	:	o_val <= 16'b0111110001100110;
            14'h3651 	:	o_val <= 16'b0111110001100111;
            14'h3652 	:	o_val <= 16'b0111110001100111;
            14'h3653 	:	o_val <= 16'b0111110001101000;
            14'h3654 	:	o_val <= 16'b0111110001101001;
            14'h3655 	:	o_val <= 16'b0111110001101010;
            14'h3656 	:	o_val <= 16'b0111110001101010;
            14'h3657 	:	o_val <= 16'b0111110001101011;
            14'h3658 	:	o_val <= 16'b0111110001101100;
            14'h3659 	:	o_val <= 16'b0111110001101101;
            14'h365a 	:	o_val <= 16'b0111110001101101;
            14'h365b 	:	o_val <= 16'b0111110001101110;
            14'h365c 	:	o_val <= 16'b0111110001101111;
            14'h365d 	:	o_val <= 16'b0111110001110000;
            14'h365e 	:	o_val <= 16'b0111110001110000;
            14'h365f 	:	o_val <= 16'b0111110001110001;
            14'h3660 	:	o_val <= 16'b0111110001110010;
            14'h3661 	:	o_val <= 16'b0111110001110011;
            14'h3662 	:	o_val <= 16'b0111110001110011;
            14'h3663 	:	o_val <= 16'b0111110001110100;
            14'h3664 	:	o_val <= 16'b0111110001110101;
            14'h3665 	:	o_val <= 16'b0111110001110101;
            14'h3666 	:	o_val <= 16'b0111110001110110;
            14'h3667 	:	o_val <= 16'b0111110001110111;
            14'h3668 	:	o_val <= 16'b0111110001111000;
            14'h3669 	:	o_val <= 16'b0111110001111000;
            14'h366a 	:	o_val <= 16'b0111110001111001;
            14'h366b 	:	o_val <= 16'b0111110001111010;
            14'h366c 	:	o_val <= 16'b0111110001111011;
            14'h366d 	:	o_val <= 16'b0111110001111011;
            14'h366e 	:	o_val <= 16'b0111110001111100;
            14'h366f 	:	o_val <= 16'b0111110001111101;
            14'h3670 	:	o_val <= 16'b0111110001111110;
            14'h3671 	:	o_val <= 16'b0111110001111110;
            14'h3672 	:	o_val <= 16'b0111110001111111;
            14'h3673 	:	o_val <= 16'b0111110010000000;
            14'h3674 	:	o_val <= 16'b0111110010000000;
            14'h3675 	:	o_val <= 16'b0111110010000001;
            14'h3676 	:	o_val <= 16'b0111110010000010;
            14'h3677 	:	o_val <= 16'b0111110010000011;
            14'h3678 	:	o_val <= 16'b0111110010000011;
            14'h3679 	:	o_val <= 16'b0111110010000100;
            14'h367a 	:	o_val <= 16'b0111110010000101;
            14'h367b 	:	o_val <= 16'b0111110010000110;
            14'h367c 	:	o_val <= 16'b0111110010000110;
            14'h367d 	:	o_val <= 16'b0111110010000111;
            14'h367e 	:	o_val <= 16'b0111110010001000;
            14'h367f 	:	o_val <= 16'b0111110010001000;
            14'h3680 	:	o_val <= 16'b0111110010001001;
            14'h3681 	:	o_val <= 16'b0111110010001010;
            14'h3682 	:	o_val <= 16'b0111110010001011;
            14'h3683 	:	o_val <= 16'b0111110010001011;
            14'h3684 	:	o_val <= 16'b0111110010001100;
            14'h3685 	:	o_val <= 16'b0111110010001101;
            14'h3686 	:	o_val <= 16'b0111110010001110;
            14'h3687 	:	o_val <= 16'b0111110010001110;
            14'h3688 	:	o_val <= 16'b0111110010001111;
            14'h3689 	:	o_val <= 16'b0111110010010000;
            14'h368a 	:	o_val <= 16'b0111110010010000;
            14'h368b 	:	o_val <= 16'b0111110010010001;
            14'h368c 	:	o_val <= 16'b0111110010010010;
            14'h368d 	:	o_val <= 16'b0111110010010011;
            14'h368e 	:	o_val <= 16'b0111110010010011;
            14'h368f 	:	o_val <= 16'b0111110010010100;
            14'h3690 	:	o_val <= 16'b0111110010010101;
            14'h3691 	:	o_val <= 16'b0111110010010101;
            14'h3692 	:	o_val <= 16'b0111110010010110;
            14'h3693 	:	o_val <= 16'b0111110010010111;
            14'h3694 	:	o_val <= 16'b0111110010011000;
            14'h3695 	:	o_val <= 16'b0111110010011000;
            14'h3696 	:	o_val <= 16'b0111110010011001;
            14'h3697 	:	o_val <= 16'b0111110010011010;
            14'h3698 	:	o_val <= 16'b0111110010011010;
            14'h3699 	:	o_val <= 16'b0111110010011011;
            14'h369a 	:	o_val <= 16'b0111110010011100;
            14'h369b 	:	o_val <= 16'b0111110010011101;
            14'h369c 	:	o_val <= 16'b0111110010011101;
            14'h369d 	:	o_val <= 16'b0111110010011110;
            14'h369e 	:	o_val <= 16'b0111110010011111;
            14'h369f 	:	o_val <= 16'b0111110010100000;
            14'h36a0 	:	o_val <= 16'b0111110010100000;
            14'h36a1 	:	o_val <= 16'b0111110010100001;
            14'h36a2 	:	o_val <= 16'b0111110010100010;
            14'h36a3 	:	o_val <= 16'b0111110010100010;
            14'h36a4 	:	o_val <= 16'b0111110010100011;
            14'h36a5 	:	o_val <= 16'b0111110010100100;
            14'h36a6 	:	o_val <= 16'b0111110010100101;
            14'h36a7 	:	o_val <= 16'b0111110010100101;
            14'h36a8 	:	o_val <= 16'b0111110010100110;
            14'h36a9 	:	o_val <= 16'b0111110010100111;
            14'h36aa 	:	o_val <= 16'b0111110010100111;
            14'h36ab 	:	o_val <= 16'b0111110010101000;
            14'h36ac 	:	o_val <= 16'b0111110010101001;
            14'h36ad 	:	o_val <= 16'b0111110010101010;
            14'h36ae 	:	o_val <= 16'b0111110010101010;
            14'h36af 	:	o_val <= 16'b0111110010101011;
            14'h36b0 	:	o_val <= 16'b0111110010101100;
            14'h36b1 	:	o_val <= 16'b0111110010101100;
            14'h36b2 	:	o_val <= 16'b0111110010101101;
            14'h36b3 	:	o_val <= 16'b0111110010101110;
            14'h36b4 	:	o_val <= 16'b0111110010101111;
            14'h36b5 	:	o_val <= 16'b0111110010101111;
            14'h36b6 	:	o_val <= 16'b0111110010110000;
            14'h36b7 	:	o_val <= 16'b0111110010110001;
            14'h36b8 	:	o_val <= 16'b0111110010110001;
            14'h36b9 	:	o_val <= 16'b0111110010110010;
            14'h36ba 	:	o_val <= 16'b0111110010110011;
            14'h36bb 	:	o_val <= 16'b0111110010110011;
            14'h36bc 	:	o_val <= 16'b0111110010110100;
            14'h36bd 	:	o_val <= 16'b0111110010110101;
            14'h36be 	:	o_val <= 16'b0111110010110110;
            14'h36bf 	:	o_val <= 16'b0111110010110110;
            14'h36c0 	:	o_val <= 16'b0111110010110111;
            14'h36c1 	:	o_val <= 16'b0111110010111000;
            14'h36c2 	:	o_val <= 16'b0111110010111000;
            14'h36c3 	:	o_val <= 16'b0111110010111001;
            14'h36c4 	:	o_val <= 16'b0111110010111010;
            14'h36c5 	:	o_val <= 16'b0111110010111011;
            14'h36c6 	:	o_val <= 16'b0111110010111011;
            14'h36c7 	:	o_val <= 16'b0111110010111100;
            14'h36c8 	:	o_val <= 16'b0111110010111101;
            14'h36c9 	:	o_val <= 16'b0111110010111101;
            14'h36ca 	:	o_val <= 16'b0111110010111110;
            14'h36cb 	:	o_val <= 16'b0111110010111111;
            14'h36cc 	:	o_val <= 16'b0111110010111111;
            14'h36cd 	:	o_val <= 16'b0111110011000000;
            14'h36ce 	:	o_val <= 16'b0111110011000001;
            14'h36cf 	:	o_val <= 16'b0111110011000010;
            14'h36d0 	:	o_val <= 16'b0111110011000010;
            14'h36d1 	:	o_val <= 16'b0111110011000011;
            14'h36d2 	:	o_val <= 16'b0111110011000100;
            14'h36d3 	:	o_val <= 16'b0111110011000100;
            14'h36d4 	:	o_val <= 16'b0111110011000101;
            14'h36d5 	:	o_val <= 16'b0111110011000110;
            14'h36d6 	:	o_val <= 16'b0111110011000110;
            14'h36d7 	:	o_val <= 16'b0111110011000111;
            14'h36d8 	:	o_val <= 16'b0111110011001000;
            14'h36d9 	:	o_val <= 16'b0111110011001001;
            14'h36da 	:	o_val <= 16'b0111110011001001;
            14'h36db 	:	o_val <= 16'b0111110011001010;
            14'h36dc 	:	o_val <= 16'b0111110011001011;
            14'h36dd 	:	o_val <= 16'b0111110011001011;
            14'h36de 	:	o_val <= 16'b0111110011001100;
            14'h36df 	:	o_val <= 16'b0111110011001101;
            14'h36e0 	:	o_val <= 16'b0111110011001101;
            14'h36e1 	:	o_val <= 16'b0111110011001110;
            14'h36e2 	:	o_val <= 16'b0111110011001111;
            14'h36e3 	:	o_val <= 16'b0111110011010000;
            14'h36e4 	:	o_val <= 16'b0111110011010000;
            14'h36e5 	:	o_val <= 16'b0111110011010001;
            14'h36e6 	:	o_val <= 16'b0111110011010010;
            14'h36e7 	:	o_val <= 16'b0111110011010010;
            14'h36e8 	:	o_val <= 16'b0111110011010011;
            14'h36e9 	:	o_val <= 16'b0111110011010100;
            14'h36ea 	:	o_val <= 16'b0111110011010100;
            14'h36eb 	:	o_val <= 16'b0111110011010101;
            14'h36ec 	:	o_val <= 16'b0111110011010110;
            14'h36ed 	:	o_val <= 16'b0111110011010111;
            14'h36ee 	:	o_val <= 16'b0111110011010111;
            14'h36ef 	:	o_val <= 16'b0111110011011000;
            14'h36f0 	:	o_val <= 16'b0111110011011001;
            14'h36f1 	:	o_val <= 16'b0111110011011001;
            14'h36f2 	:	o_val <= 16'b0111110011011010;
            14'h36f3 	:	o_val <= 16'b0111110011011011;
            14'h36f4 	:	o_val <= 16'b0111110011011011;
            14'h36f5 	:	o_val <= 16'b0111110011011100;
            14'h36f6 	:	o_val <= 16'b0111110011011101;
            14'h36f7 	:	o_val <= 16'b0111110011011101;
            14'h36f8 	:	o_val <= 16'b0111110011011110;
            14'h36f9 	:	o_val <= 16'b0111110011011111;
            14'h36fa 	:	o_val <= 16'b0111110011100000;
            14'h36fb 	:	o_val <= 16'b0111110011100000;
            14'h36fc 	:	o_val <= 16'b0111110011100001;
            14'h36fd 	:	o_val <= 16'b0111110011100010;
            14'h36fe 	:	o_val <= 16'b0111110011100010;
            14'h36ff 	:	o_val <= 16'b0111110011100011;
            14'h3700 	:	o_val <= 16'b0111110011100100;
            14'h3701 	:	o_val <= 16'b0111110011100100;
            14'h3702 	:	o_val <= 16'b0111110011100101;
            14'h3703 	:	o_val <= 16'b0111110011100110;
            14'h3704 	:	o_val <= 16'b0111110011100110;
            14'h3705 	:	o_val <= 16'b0111110011100111;
            14'h3706 	:	o_val <= 16'b0111110011101000;
            14'h3707 	:	o_val <= 16'b0111110011101000;
            14'h3708 	:	o_val <= 16'b0111110011101001;
            14'h3709 	:	o_val <= 16'b0111110011101010;
            14'h370a 	:	o_val <= 16'b0111110011101011;
            14'h370b 	:	o_val <= 16'b0111110011101011;
            14'h370c 	:	o_val <= 16'b0111110011101100;
            14'h370d 	:	o_val <= 16'b0111110011101101;
            14'h370e 	:	o_val <= 16'b0111110011101101;
            14'h370f 	:	o_val <= 16'b0111110011101110;
            14'h3710 	:	o_val <= 16'b0111110011101111;
            14'h3711 	:	o_val <= 16'b0111110011101111;
            14'h3712 	:	o_val <= 16'b0111110011110000;
            14'h3713 	:	o_val <= 16'b0111110011110001;
            14'h3714 	:	o_val <= 16'b0111110011110001;
            14'h3715 	:	o_val <= 16'b0111110011110010;
            14'h3716 	:	o_val <= 16'b0111110011110011;
            14'h3717 	:	o_val <= 16'b0111110011110011;
            14'h3718 	:	o_val <= 16'b0111110011110100;
            14'h3719 	:	o_val <= 16'b0111110011110101;
            14'h371a 	:	o_val <= 16'b0111110011110101;
            14'h371b 	:	o_val <= 16'b0111110011110110;
            14'h371c 	:	o_val <= 16'b0111110011110111;
            14'h371d 	:	o_val <= 16'b0111110011110111;
            14'h371e 	:	o_val <= 16'b0111110011111000;
            14'h371f 	:	o_val <= 16'b0111110011111001;
            14'h3720 	:	o_val <= 16'b0111110011111010;
            14'h3721 	:	o_val <= 16'b0111110011111010;
            14'h3722 	:	o_val <= 16'b0111110011111011;
            14'h3723 	:	o_val <= 16'b0111110011111100;
            14'h3724 	:	o_val <= 16'b0111110011111100;
            14'h3725 	:	o_val <= 16'b0111110011111101;
            14'h3726 	:	o_val <= 16'b0111110011111110;
            14'h3727 	:	o_val <= 16'b0111110011111110;
            14'h3728 	:	o_val <= 16'b0111110011111111;
            14'h3729 	:	o_val <= 16'b0111110100000000;
            14'h372a 	:	o_val <= 16'b0111110100000000;
            14'h372b 	:	o_val <= 16'b0111110100000001;
            14'h372c 	:	o_val <= 16'b0111110100000010;
            14'h372d 	:	o_val <= 16'b0111110100000010;
            14'h372e 	:	o_val <= 16'b0111110100000011;
            14'h372f 	:	o_val <= 16'b0111110100000100;
            14'h3730 	:	o_val <= 16'b0111110100000100;
            14'h3731 	:	o_val <= 16'b0111110100000101;
            14'h3732 	:	o_val <= 16'b0111110100000110;
            14'h3733 	:	o_val <= 16'b0111110100000110;
            14'h3734 	:	o_val <= 16'b0111110100000111;
            14'h3735 	:	o_val <= 16'b0111110100001000;
            14'h3736 	:	o_val <= 16'b0111110100001000;
            14'h3737 	:	o_val <= 16'b0111110100001001;
            14'h3738 	:	o_val <= 16'b0111110100001010;
            14'h3739 	:	o_val <= 16'b0111110100001010;
            14'h373a 	:	o_val <= 16'b0111110100001011;
            14'h373b 	:	o_val <= 16'b0111110100001100;
            14'h373c 	:	o_val <= 16'b0111110100001100;
            14'h373d 	:	o_val <= 16'b0111110100001101;
            14'h373e 	:	o_val <= 16'b0111110100001110;
            14'h373f 	:	o_val <= 16'b0111110100001110;
            14'h3740 	:	o_val <= 16'b0111110100001111;
            14'h3741 	:	o_val <= 16'b0111110100010000;
            14'h3742 	:	o_val <= 16'b0111110100010000;
            14'h3743 	:	o_val <= 16'b0111110100010001;
            14'h3744 	:	o_val <= 16'b0111110100010010;
            14'h3745 	:	o_val <= 16'b0111110100010010;
            14'h3746 	:	o_val <= 16'b0111110100010011;
            14'h3747 	:	o_val <= 16'b0111110100010100;
            14'h3748 	:	o_val <= 16'b0111110100010100;
            14'h3749 	:	o_val <= 16'b0111110100010101;
            14'h374a 	:	o_val <= 16'b0111110100010110;
            14'h374b 	:	o_val <= 16'b0111110100010110;
            14'h374c 	:	o_val <= 16'b0111110100010111;
            14'h374d 	:	o_val <= 16'b0111110100011000;
            14'h374e 	:	o_val <= 16'b0111110100011000;
            14'h374f 	:	o_val <= 16'b0111110100011001;
            14'h3750 	:	o_val <= 16'b0111110100011010;
            14'h3751 	:	o_val <= 16'b0111110100011010;
            14'h3752 	:	o_val <= 16'b0111110100011011;
            14'h3753 	:	o_val <= 16'b0111110100011100;
            14'h3754 	:	o_val <= 16'b0111110100011100;
            14'h3755 	:	o_val <= 16'b0111110100011101;
            14'h3756 	:	o_val <= 16'b0111110100011110;
            14'h3757 	:	o_val <= 16'b0111110100011110;
            14'h3758 	:	o_val <= 16'b0111110100011111;
            14'h3759 	:	o_val <= 16'b0111110100100000;
            14'h375a 	:	o_val <= 16'b0111110100100000;
            14'h375b 	:	o_val <= 16'b0111110100100001;
            14'h375c 	:	o_val <= 16'b0111110100100010;
            14'h375d 	:	o_val <= 16'b0111110100100010;
            14'h375e 	:	o_val <= 16'b0111110100100011;
            14'h375f 	:	o_val <= 16'b0111110100100100;
            14'h3760 	:	o_val <= 16'b0111110100100100;
            14'h3761 	:	o_val <= 16'b0111110100100101;
            14'h3762 	:	o_val <= 16'b0111110100100110;
            14'h3763 	:	o_val <= 16'b0111110100100110;
            14'h3764 	:	o_val <= 16'b0111110100100111;
            14'h3765 	:	o_val <= 16'b0111110100101000;
            14'h3766 	:	o_val <= 16'b0111110100101000;
            14'h3767 	:	o_val <= 16'b0111110100101001;
            14'h3768 	:	o_val <= 16'b0111110100101010;
            14'h3769 	:	o_val <= 16'b0111110100101010;
            14'h376a 	:	o_val <= 16'b0111110100101011;
            14'h376b 	:	o_val <= 16'b0111110100101100;
            14'h376c 	:	o_val <= 16'b0111110100101100;
            14'h376d 	:	o_val <= 16'b0111110100101101;
            14'h376e 	:	o_val <= 16'b0111110100101110;
            14'h376f 	:	o_val <= 16'b0111110100101110;
            14'h3770 	:	o_val <= 16'b0111110100101111;
            14'h3771 	:	o_val <= 16'b0111110100110000;
            14'h3772 	:	o_val <= 16'b0111110100110000;
            14'h3773 	:	o_val <= 16'b0111110100110001;
            14'h3774 	:	o_val <= 16'b0111110100110010;
            14'h3775 	:	o_val <= 16'b0111110100110010;
            14'h3776 	:	o_val <= 16'b0111110100110011;
            14'h3777 	:	o_val <= 16'b0111110100110011;
            14'h3778 	:	o_val <= 16'b0111110100110100;
            14'h3779 	:	o_val <= 16'b0111110100110101;
            14'h377a 	:	o_val <= 16'b0111110100110101;
            14'h377b 	:	o_val <= 16'b0111110100110110;
            14'h377c 	:	o_val <= 16'b0111110100110111;
            14'h377d 	:	o_val <= 16'b0111110100110111;
            14'h377e 	:	o_val <= 16'b0111110100111000;
            14'h377f 	:	o_val <= 16'b0111110100111001;
            14'h3780 	:	o_val <= 16'b0111110100111001;
            14'h3781 	:	o_val <= 16'b0111110100111010;
            14'h3782 	:	o_val <= 16'b0111110100111011;
            14'h3783 	:	o_val <= 16'b0111110100111011;
            14'h3784 	:	o_val <= 16'b0111110100111100;
            14'h3785 	:	o_val <= 16'b0111110100111101;
            14'h3786 	:	o_val <= 16'b0111110100111101;
            14'h3787 	:	o_val <= 16'b0111110100111110;
            14'h3788 	:	o_val <= 16'b0111110100111111;
            14'h3789 	:	o_val <= 16'b0111110100111111;
            14'h378a 	:	o_val <= 16'b0111110101000000;
            14'h378b 	:	o_val <= 16'b0111110101000000;
            14'h378c 	:	o_val <= 16'b0111110101000001;
            14'h378d 	:	o_val <= 16'b0111110101000010;
            14'h378e 	:	o_val <= 16'b0111110101000010;
            14'h378f 	:	o_val <= 16'b0111110101000011;
            14'h3790 	:	o_val <= 16'b0111110101000100;
            14'h3791 	:	o_val <= 16'b0111110101000100;
            14'h3792 	:	o_val <= 16'b0111110101000101;
            14'h3793 	:	o_val <= 16'b0111110101000110;
            14'h3794 	:	o_val <= 16'b0111110101000110;
            14'h3795 	:	o_val <= 16'b0111110101000111;
            14'h3796 	:	o_val <= 16'b0111110101001000;
            14'h3797 	:	o_val <= 16'b0111110101001000;
            14'h3798 	:	o_val <= 16'b0111110101001001;
            14'h3799 	:	o_val <= 16'b0111110101001001;
            14'h379a 	:	o_val <= 16'b0111110101001010;
            14'h379b 	:	o_val <= 16'b0111110101001011;
            14'h379c 	:	o_val <= 16'b0111110101001011;
            14'h379d 	:	o_val <= 16'b0111110101001100;
            14'h379e 	:	o_val <= 16'b0111110101001101;
            14'h379f 	:	o_val <= 16'b0111110101001101;
            14'h37a0 	:	o_val <= 16'b0111110101001110;
            14'h37a1 	:	o_val <= 16'b0111110101001111;
            14'h37a2 	:	o_val <= 16'b0111110101001111;
            14'h37a3 	:	o_val <= 16'b0111110101010000;
            14'h37a4 	:	o_val <= 16'b0111110101010001;
            14'h37a5 	:	o_val <= 16'b0111110101010001;
            14'h37a6 	:	o_val <= 16'b0111110101010010;
            14'h37a7 	:	o_val <= 16'b0111110101010010;
            14'h37a8 	:	o_val <= 16'b0111110101010011;
            14'h37a9 	:	o_val <= 16'b0111110101010100;
            14'h37aa 	:	o_val <= 16'b0111110101010100;
            14'h37ab 	:	o_val <= 16'b0111110101010101;
            14'h37ac 	:	o_val <= 16'b0111110101010110;
            14'h37ad 	:	o_val <= 16'b0111110101010110;
            14'h37ae 	:	o_val <= 16'b0111110101010111;
            14'h37af 	:	o_val <= 16'b0111110101011000;
            14'h37b0 	:	o_val <= 16'b0111110101011000;
            14'h37b1 	:	o_val <= 16'b0111110101011001;
            14'h37b2 	:	o_val <= 16'b0111110101011001;
            14'h37b3 	:	o_val <= 16'b0111110101011010;
            14'h37b4 	:	o_val <= 16'b0111110101011011;
            14'h37b5 	:	o_val <= 16'b0111110101011011;
            14'h37b6 	:	o_val <= 16'b0111110101011100;
            14'h37b7 	:	o_val <= 16'b0111110101011101;
            14'h37b8 	:	o_val <= 16'b0111110101011101;
            14'h37b9 	:	o_val <= 16'b0111110101011110;
            14'h37ba 	:	o_val <= 16'b0111110101011111;
            14'h37bb 	:	o_val <= 16'b0111110101011111;
            14'h37bc 	:	o_val <= 16'b0111110101100000;
            14'h37bd 	:	o_val <= 16'b0111110101100000;
            14'h37be 	:	o_val <= 16'b0111110101100001;
            14'h37bf 	:	o_val <= 16'b0111110101100010;
            14'h37c0 	:	o_val <= 16'b0111110101100010;
            14'h37c1 	:	o_val <= 16'b0111110101100011;
            14'h37c2 	:	o_val <= 16'b0111110101100100;
            14'h37c3 	:	o_val <= 16'b0111110101100100;
            14'h37c4 	:	o_val <= 16'b0111110101100101;
            14'h37c5 	:	o_val <= 16'b0111110101100110;
            14'h37c6 	:	o_val <= 16'b0111110101100110;
            14'h37c7 	:	o_val <= 16'b0111110101100111;
            14'h37c8 	:	o_val <= 16'b0111110101100111;
            14'h37c9 	:	o_val <= 16'b0111110101101000;
            14'h37ca 	:	o_val <= 16'b0111110101101001;
            14'h37cb 	:	o_val <= 16'b0111110101101001;
            14'h37cc 	:	o_val <= 16'b0111110101101010;
            14'h37cd 	:	o_val <= 16'b0111110101101011;
            14'h37ce 	:	o_val <= 16'b0111110101101011;
            14'h37cf 	:	o_val <= 16'b0111110101101100;
            14'h37d0 	:	o_val <= 16'b0111110101101100;
            14'h37d1 	:	o_val <= 16'b0111110101101101;
            14'h37d2 	:	o_val <= 16'b0111110101101110;
            14'h37d3 	:	o_val <= 16'b0111110101101110;
            14'h37d4 	:	o_val <= 16'b0111110101101111;
            14'h37d5 	:	o_val <= 16'b0111110101110000;
            14'h37d6 	:	o_val <= 16'b0111110101110000;
            14'h37d7 	:	o_val <= 16'b0111110101110001;
            14'h37d8 	:	o_val <= 16'b0111110101110001;
            14'h37d9 	:	o_val <= 16'b0111110101110010;
            14'h37da 	:	o_val <= 16'b0111110101110011;
            14'h37db 	:	o_val <= 16'b0111110101110011;
            14'h37dc 	:	o_val <= 16'b0111110101110100;
            14'h37dd 	:	o_val <= 16'b0111110101110101;
            14'h37de 	:	o_val <= 16'b0111110101110101;
            14'h37df 	:	o_val <= 16'b0111110101110110;
            14'h37e0 	:	o_val <= 16'b0111110101110110;
            14'h37e1 	:	o_val <= 16'b0111110101110111;
            14'h37e2 	:	o_val <= 16'b0111110101111000;
            14'h37e3 	:	o_val <= 16'b0111110101111000;
            14'h37e4 	:	o_val <= 16'b0111110101111001;
            14'h37e5 	:	o_val <= 16'b0111110101111010;
            14'h37e6 	:	o_val <= 16'b0111110101111010;
            14'h37e7 	:	o_val <= 16'b0111110101111011;
            14'h37e8 	:	o_val <= 16'b0111110101111011;
            14'h37e9 	:	o_val <= 16'b0111110101111100;
            14'h37ea 	:	o_val <= 16'b0111110101111101;
            14'h37eb 	:	o_val <= 16'b0111110101111101;
            14'h37ec 	:	o_val <= 16'b0111110101111110;
            14'h37ed 	:	o_val <= 16'b0111110101111110;
            14'h37ee 	:	o_val <= 16'b0111110101111111;
            14'h37ef 	:	o_val <= 16'b0111110110000000;
            14'h37f0 	:	o_val <= 16'b0111110110000000;
            14'h37f1 	:	o_val <= 16'b0111110110000001;
            14'h37f2 	:	o_val <= 16'b0111110110000010;
            14'h37f3 	:	o_val <= 16'b0111110110000010;
            14'h37f4 	:	o_val <= 16'b0111110110000011;
            14'h37f5 	:	o_val <= 16'b0111110110000011;
            14'h37f6 	:	o_val <= 16'b0111110110000100;
            14'h37f7 	:	o_val <= 16'b0111110110000101;
            14'h37f8 	:	o_val <= 16'b0111110110000101;
            14'h37f9 	:	o_val <= 16'b0111110110000110;
            14'h37fa 	:	o_val <= 16'b0111110110000110;
            14'h37fb 	:	o_val <= 16'b0111110110000111;
            14'h37fc 	:	o_val <= 16'b0111110110001000;
            14'h37fd 	:	o_val <= 16'b0111110110001000;
            14'h37fe 	:	o_val <= 16'b0111110110001001;
            14'h37ff 	:	o_val <= 16'b0111110110001010;
            14'h3800 	:	o_val <= 16'b0111110110001010;
            14'h3801 	:	o_val <= 16'b0111110110001011;
            14'h3802 	:	o_val <= 16'b0111110110001011;
            14'h3803 	:	o_val <= 16'b0111110110001100;
            14'h3804 	:	o_val <= 16'b0111110110001101;
            14'h3805 	:	o_val <= 16'b0111110110001101;
            14'h3806 	:	o_val <= 16'b0111110110001110;
            14'h3807 	:	o_val <= 16'b0111110110001110;
            14'h3808 	:	o_val <= 16'b0111110110001111;
            14'h3809 	:	o_val <= 16'b0111110110010000;
            14'h380a 	:	o_val <= 16'b0111110110010000;
            14'h380b 	:	o_val <= 16'b0111110110010001;
            14'h380c 	:	o_val <= 16'b0111110110010010;
            14'h380d 	:	o_val <= 16'b0111110110010010;
            14'h380e 	:	o_val <= 16'b0111110110010011;
            14'h380f 	:	o_val <= 16'b0111110110010011;
            14'h3810 	:	o_val <= 16'b0111110110010100;
            14'h3811 	:	o_val <= 16'b0111110110010101;
            14'h3812 	:	o_val <= 16'b0111110110010101;
            14'h3813 	:	o_val <= 16'b0111110110010110;
            14'h3814 	:	o_val <= 16'b0111110110010110;
            14'h3815 	:	o_val <= 16'b0111110110010111;
            14'h3816 	:	o_val <= 16'b0111110110011000;
            14'h3817 	:	o_val <= 16'b0111110110011000;
            14'h3818 	:	o_val <= 16'b0111110110011001;
            14'h3819 	:	o_val <= 16'b0111110110011001;
            14'h381a 	:	o_val <= 16'b0111110110011010;
            14'h381b 	:	o_val <= 16'b0111110110011011;
            14'h381c 	:	o_val <= 16'b0111110110011011;
            14'h381d 	:	o_val <= 16'b0111110110011100;
            14'h381e 	:	o_val <= 16'b0111110110011100;
            14'h381f 	:	o_val <= 16'b0111110110011101;
            14'h3820 	:	o_val <= 16'b0111110110011110;
            14'h3821 	:	o_val <= 16'b0111110110011110;
            14'h3822 	:	o_val <= 16'b0111110110011111;
            14'h3823 	:	o_val <= 16'b0111110110011111;
            14'h3824 	:	o_val <= 16'b0111110110100000;
            14'h3825 	:	o_val <= 16'b0111110110100001;
            14'h3826 	:	o_val <= 16'b0111110110100001;
            14'h3827 	:	o_val <= 16'b0111110110100010;
            14'h3828 	:	o_val <= 16'b0111110110100010;
            14'h3829 	:	o_val <= 16'b0111110110100011;
            14'h382a 	:	o_val <= 16'b0111110110100100;
            14'h382b 	:	o_val <= 16'b0111110110100100;
            14'h382c 	:	o_val <= 16'b0111110110100101;
            14'h382d 	:	o_val <= 16'b0111110110100101;
            14'h382e 	:	o_val <= 16'b0111110110100110;
            14'h382f 	:	o_val <= 16'b0111110110100111;
            14'h3830 	:	o_val <= 16'b0111110110100111;
            14'h3831 	:	o_val <= 16'b0111110110101000;
            14'h3832 	:	o_val <= 16'b0111110110101000;
            14'h3833 	:	o_val <= 16'b0111110110101001;
            14'h3834 	:	o_val <= 16'b0111110110101010;
            14'h3835 	:	o_val <= 16'b0111110110101010;
            14'h3836 	:	o_val <= 16'b0111110110101011;
            14'h3837 	:	o_val <= 16'b0111110110101011;
            14'h3838 	:	o_val <= 16'b0111110110101100;
            14'h3839 	:	o_val <= 16'b0111110110101101;
            14'h383a 	:	o_val <= 16'b0111110110101101;
            14'h383b 	:	o_val <= 16'b0111110110101110;
            14'h383c 	:	o_val <= 16'b0111110110101110;
            14'h383d 	:	o_val <= 16'b0111110110101111;
            14'h383e 	:	o_val <= 16'b0111110110110000;
            14'h383f 	:	o_val <= 16'b0111110110110000;
            14'h3840 	:	o_val <= 16'b0111110110110001;
            14'h3841 	:	o_val <= 16'b0111110110110001;
            14'h3842 	:	o_val <= 16'b0111110110110010;
            14'h3843 	:	o_val <= 16'b0111110110110011;
            14'h3844 	:	o_val <= 16'b0111110110110011;
            14'h3845 	:	o_val <= 16'b0111110110110100;
            14'h3846 	:	o_val <= 16'b0111110110110100;
            14'h3847 	:	o_val <= 16'b0111110110110101;
            14'h3848 	:	o_val <= 16'b0111110110110110;
            14'h3849 	:	o_val <= 16'b0111110110110110;
            14'h384a 	:	o_val <= 16'b0111110110110111;
            14'h384b 	:	o_val <= 16'b0111110110110111;
            14'h384c 	:	o_val <= 16'b0111110110111000;
            14'h384d 	:	o_val <= 16'b0111110110111000;
            14'h384e 	:	o_val <= 16'b0111110110111001;
            14'h384f 	:	o_val <= 16'b0111110110111010;
            14'h3850 	:	o_val <= 16'b0111110110111010;
            14'h3851 	:	o_val <= 16'b0111110110111011;
            14'h3852 	:	o_val <= 16'b0111110110111011;
            14'h3853 	:	o_val <= 16'b0111110110111100;
            14'h3854 	:	o_val <= 16'b0111110110111101;
            14'h3855 	:	o_val <= 16'b0111110110111101;
            14'h3856 	:	o_val <= 16'b0111110110111110;
            14'h3857 	:	o_val <= 16'b0111110110111110;
            14'h3858 	:	o_val <= 16'b0111110110111111;
            14'h3859 	:	o_val <= 16'b0111110111000000;
            14'h385a 	:	o_val <= 16'b0111110111000000;
            14'h385b 	:	o_val <= 16'b0111110111000001;
            14'h385c 	:	o_val <= 16'b0111110111000001;
            14'h385d 	:	o_val <= 16'b0111110111000010;
            14'h385e 	:	o_val <= 16'b0111110111000010;
            14'h385f 	:	o_val <= 16'b0111110111000011;
            14'h3860 	:	o_val <= 16'b0111110111000100;
            14'h3861 	:	o_val <= 16'b0111110111000100;
            14'h3862 	:	o_val <= 16'b0111110111000101;
            14'h3863 	:	o_val <= 16'b0111110111000101;
            14'h3864 	:	o_val <= 16'b0111110111000110;
            14'h3865 	:	o_val <= 16'b0111110111000111;
            14'h3866 	:	o_val <= 16'b0111110111000111;
            14'h3867 	:	o_val <= 16'b0111110111001000;
            14'h3868 	:	o_val <= 16'b0111110111001000;
            14'h3869 	:	o_val <= 16'b0111110111001001;
            14'h386a 	:	o_val <= 16'b0111110111001001;
            14'h386b 	:	o_val <= 16'b0111110111001010;
            14'h386c 	:	o_val <= 16'b0111110111001011;
            14'h386d 	:	o_val <= 16'b0111110111001011;
            14'h386e 	:	o_val <= 16'b0111110111001100;
            14'h386f 	:	o_val <= 16'b0111110111001100;
            14'h3870 	:	o_val <= 16'b0111110111001101;
            14'h3871 	:	o_val <= 16'b0111110111001110;
            14'h3872 	:	o_val <= 16'b0111110111001110;
            14'h3873 	:	o_val <= 16'b0111110111001111;
            14'h3874 	:	o_val <= 16'b0111110111001111;
            14'h3875 	:	o_val <= 16'b0111110111010000;
            14'h3876 	:	o_val <= 16'b0111110111010000;
            14'h3877 	:	o_val <= 16'b0111110111010001;
            14'h3878 	:	o_val <= 16'b0111110111010010;
            14'h3879 	:	o_val <= 16'b0111110111010010;
            14'h387a 	:	o_val <= 16'b0111110111010011;
            14'h387b 	:	o_val <= 16'b0111110111010011;
            14'h387c 	:	o_val <= 16'b0111110111010100;
            14'h387d 	:	o_val <= 16'b0111110111010100;
            14'h387e 	:	o_val <= 16'b0111110111010101;
            14'h387f 	:	o_val <= 16'b0111110111010110;
            14'h3880 	:	o_val <= 16'b0111110111010110;
            14'h3881 	:	o_val <= 16'b0111110111010111;
            14'h3882 	:	o_val <= 16'b0111110111010111;
            14'h3883 	:	o_val <= 16'b0111110111011000;
            14'h3884 	:	o_val <= 16'b0111110111011000;
            14'h3885 	:	o_val <= 16'b0111110111011001;
            14'h3886 	:	o_val <= 16'b0111110111011010;
            14'h3887 	:	o_val <= 16'b0111110111011010;
            14'h3888 	:	o_val <= 16'b0111110111011011;
            14'h3889 	:	o_val <= 16'b0111110111011011;
            14'h388a 	:	o_val <= 16'b0111110111011100;
            14'h388b 	:	o_val <= 16'b0111110111011100;
            14'h388c 	:	o_val <= 16'b0111110111011101;
            14'h388d 	:	o_val <= 16'b0111110111011110;
            14'h388e 	:	o_val <= 16'b0111110111011110;
            14'h388f 	:	o_val <= 16'b0111110111011111;
            14'h3890 	:	o_val <= 16'b0111110111011111;
            14'h3891 	:	o_val <= 16'b0111110111100000;
            14'h3892 	:	o_val <= 16'b0111110111100000;
            14'h3893 	:	o_val <= 16'b0111110111100001;
            14'h3894 	:	o_val <= 16'b0111110111100010;
            14'h3895 	:	o_val <= 16'b0111110111100010;
            14'h3896 	:	o_val <= 16'b0111110111100011;
            14'h3897 	:	o_val <= 16'b0111110111100011;
            14'h3898 	:	o_val <= 16'b0111110111100100;
            14'h3899 	:	o_val <= 16'b0111110111100100;
            14'h389a 	:	o_val <= 16'b0111110111100101;
            14'h389b 	:	o_val <= 16'b0111110111100110;
            14'h389c 	:	o_val <= 16'b0111110111100110;
            14'h389d 	:	o_val <= 16'b0111110111100111;
            14'h389e 	:	o_val <= 16'b0111110111100111;
            14'h389f 	:	o_val <= 16'b0111110111101000;
            14'h38a0 	:	o_val <= 16'b0111110111101000;
            14'h38a1 	:	o_val <= 16'b0111110111101001;
            14'h38a2 	:	o_val <= 16'b0111110111101010;
            14'h38a3 	:	o_val <= 16'b0111110111101010;
            14'h38a4 	:	o_val <= 16'b0111110111101011;
            14'h38a5 	:	o_val <= 16'b0111110111101011;
            14'h38a6 	:	o_val <= 16'b0111110111101100;
            14'h38a7 	:	o_val <= 16'b0111110111101100;
            14'h38a8 	:	o_val <= 16'b0111110111101101;
            14'h38a9 	:	o_val <= 16'b0111110111101110;
            14'h38aa 	:	o_val <= 16'b0111110111101110;
            14'h38ab 	:	o_val <= 16'b0111110111101111;
            14'h38ac 	:	o_val <= 16'b0111110111101111;
            14'h38ad 	:	o_val <= 16'b0111110111110000;
            14'h38ae 	:	o_val <= 16'b0111110111110000;
            14'h38af 	:	o_val <= 16'b0111110111110001;
            14'h38b0 	:	o_val <= 16'b0111110111110001;
            14'h38b1 	:	o_val <= 16'b0111110111110010;
            14'h38b2 	:	o_val <= 16'b0111110111110011;
            14'h38b3 	:	o_val <= 16'b0111110111110011;
            14'h38b4 	:	o_val <= 16'b0111110111110100;
            14'h38b5 	:	o_val <= 16'b0111110111110100;
            14'h38b6 	:	o_val <= 16'b0111110111110101;
            14'h38b7 	:	o_val <= 16'b0111110111110101;
            14'h38b8 	:	o_val <= 16'b0111110111110110;
            14'h38b9 	:	o_val <= 16'b0111110111110110;
            14'h38ba 	:	o_val <= 16'b0111110111110111;
            14'h38bb 	:	o_val <= 16'b0111110111111000;
            14'h38bc 	:	o_val <= 16'b0111110111111000;
            14'h38bd 	:	o_val <= 16'b0111110111111001;
            14'h38be 	:	o_val <= 16'b0111110111111001;
            14'h38bf 	:	o_val <= 16'b0111110111111010;
            14'h38c0 	:	o_val <= 16'b0111110111111010;
            14'h38c1 	:	o_val <= 16'b0111110111111011;
            14'h38c2 	:	o_val <= 16'b0111110111111011;
            14'h38c3 	:	o_val <= 16'b0111110111111100;
            14'h38c4 	:	o_val <= 16'b0111110111111101;
            14'h38c5 	:	o_val <= 16'b0111110111111101;
            14'h38c6 	:	o_val <= 16'b0111110111111110;
            14'h38c7 	:	o_val <= 16'b0111110111111110;
            14'h38c8 	:	o_val <= 16'b0111110111111111;
            14'h38c9 	:	o_val <= 16'b0111110111111111;
            14'h38ca 	:	o_val <= 16'b0111111000000000;
            14'h38cb 	:	o_val <= 16'b0111111000000000;
            14'h38cc 	:	o_val <= 16'b0111111000000001;
            14'h38cd 	:	o_val <= 16'b0111111000000010;
            14'h38ce 	:	o_val <= 16'b0111111000000010;
            14'h38cf 	:	o_val <= 16'b0111111000000011;
            14'h38d0 	:	o_val <= 16'b0111111000000011;
            14'h38d1 	:	o_val <= 16'b0111111000000100;
            14'h38d2 	:	o_val <= 16'b0111111000000100;
            14'h38d3 	:	o_val <= 16'b0111111000000101;
            14'h38d4 	:	o_val <= 16'b0111111000000101;
            14'h38d5 	:	o_val <= 16'b0111111000000110;
            14'h38d6 	:	o_val <= 16'b0111111000000111;
            14'h38d7 	:	o_val <= 16'b0111111000000111;
            14'h38d8 	:	o_val <= 16'b0111111000001000;
            14'h38d9 	:	o_val <= 16'b0111111000001000;
            14'h38da 	:	o_val <= 16'b0111111000001001;
            14'h38db 	:	o_val <= 16'b0111111000001001;
            14'h38dc 	:	o_val <= 16'b0111111000001010;
            14'h38dd 	:	o_val <= 16'b0111111000001010;
            14'h38de 	:	o_val <= 16'b0111111000001011;
            14'h38df 	:	o_val <= 16'b0111111000001011;
            14'h38e0 	:	o_val <= 16'b0111111000001100;
            14'h38e1 	:	o_val <= 16'b0111111000001101;
            14'h38e2 	:	o_val <= 16'b0111111000001101;
            14'h38e3 	:	o_val <= 16'b0111111000001110;
            14'h38e4 	:	o_val <= 16'b0111111000001110;
            14'h38e5 	:	o_val <= 16'b0111111000001111;
            14'h38e6 	:	o_val <= 16'b0111111000001111;
            14'h38e7 	:	o_val <= 16'b0111111000010000;
            14'h38e8 	:	o_val <= 16'b0111111000010000;
            14'h38e9 	:	o_val <= 16'b0111111000010001;
            14'h38ea 	:	o_val <= 16'b0111111000010001;
            14'h38eb 	:	o_val <= 16'b0111111000010010;
            14'h38ec 	:	o_val <= 16'b0111111000010011;
            14'h38ed 	:	o_val <= 16'b0111111000010011;
            14'h38ee 	:	o_val <= 16'b0111111000010100;
            14'h38ef 	:	o_val <= 16'b0111111000010100;
            14'h38f0 	:	o_val <= 16'b0111111000010101;
            14'h38f1 	:	o_val <= 16'b0111111000010101;
            14'h38f2 	:	o_val <= 16'b0111111000010110;
            14'h38f3 	:	o_val <= 16'b0111111000010110;
            14'h38f4 	:	o_val <= 16'b0111111000010111;
            14'h38f5 	:	o_val <= 16'b0111111000010111;
            14'h38f6 	:	o_val <= 16'b0111111000011000;
            14'h38f7 	:	o_val <= 16'b0111111000011001;
            14'h38f8 	:	o_val <= 16'b0111111000011001;
            14'h38f9 	:	o_val <= 16'b0111111000011010;
            14'h38fa 	:	o_val <= 16'b0111111000011010;
            14'h38fb 	:	o_val <= 16'b0111111000011011;
            14'h38fc 	:	o_val <= 16'b0111111000011011;
            14'h38fd 	:	o_val <= 16'b0111111000011100;
            14'h38fe 	:	o_val <= 16'b0111111000011100;
            14'h38ff 	:	o_val <= 16'b0111111000011101;
            14'h3900 	:	o_val <= 16'b0111111000011101;
            14'h3901 	:	o_val <= 16'b0111111000011110;
            14'h3902 	:	o_val <= 16'b0111111000011110;
            14'h3903 	:	o_val <= 16'b0111111000011111;
            14'h3904 	:	o_val <= 16'b0111111000011111;
            14'h3905 	:	o_val <= 16'b0111111000100000;
            14'h3906 	:	o_val <= 16'b0111111000100001;
            14'h3907 	:	o_val <= 16'b0111111000100001;
            14'h3908 	:	o_val <= 16'b0111111000100010;
            14'h3909 	:	o_val <= 16'b0111111000100010;
            14'h390a 	:	o_val <= 16'b0111111000100011;
            14'h390b 	:	o_val <= 16'b0111111000100011;
            14'h390c 	:	o_val <= 16'b0111111000100100;
            14'h390d 	:	o_val <= 16'b0111111000100100;
            14'h390e 	:	o_val <= 16'b0111111000100101;
            14'h390f 	:	o_val <= 16'b0111111000100101;
            14'h3910 	:	o_val <= 16'b0111111000100110;
            14'h3911 	:	o_val <= 16'b0111111000100110;
            14'h3912 	:	o_val <= 16'b0111111000100111;
            14'h3913 	:	o_val <= 16'b0111111000100111;
            14'h3914 	:	o_val <= 16'b0111111000101000;
            14'h3915 	:	o_val <= 16'b0111111000101001;
            14'h3916 	:	o_val <= 16'b0111111000101001;
            14'h3917 	:	o_val <= 16'b0111111000101010;
            14'h3918 	:	o_val <= 16'b0111111000101010;
            14'h3919 	:	o_val <= 16'b0111111000101011;
            14'h391a 	:	o_val <= 16'b0111111000101011;
            14'h391b 	:	o_val <= 16'b0111111000101100;
            14'h391c 	:	o_val <= 16'b0111111000101100;
            14'h391d 	:	o_val <= 16'b0111111000101101;
            14'h391e 	:	o_val <= 16'b0111111000101101;
            14'h391f 	:	o_val <= 16'b0111111000101110;
            14'h3920 	:	o_val <= 16'b0111111000101110;
            14'h3921 	:	o_val <= 16'b0111111000101111;
            14'h3922 	:	o_val <= 16'b0111111000101111;
            14'h3923 	:	o_val <= 16'b0111111000110000;
            14'h3924 	:	o_val <= 16'b0111111000110000;
            14'h3925 	:	o_val <= 16'b0111111000110001;
            14'h3926 	:	o_val <= 16'b0111111000110010;
            14'h3927 	:	o_val <= 16'b0111111000110010;
            14'h3928 	:	o_val <= 16'b0111111000110011;
            14'h3929 	:	o_val <= 16'b0111111000110011;
            14'h392a 	:	o_val <= 16'b0111111000110100;
            14'h392b 	:	o_val <= 16'b0111111000110100;
            14'h392c 	:	o_val <= 16'b0111111000110101;
            14'h392d 	:	o_val <= 16'b0111111000110101;
            14'h392e 	:	o_val <= 16'b0111111000110110;
            14'h392f 	:	o_val <= 16'b0111111000110110;
            14'h3930 	:	o_val <= 16'b0111111000110111;
            14'h3931 	:	o_val <= 16'b0111111000110111;
            14'h3932 	:	o_val <= 16'b0111111000111000;
            14'h3933 	:	o_val <= 16'b0111111000111000;
            14'h3934 	:	o_val <= 16'b0111111000111001;
            14'h3935 	:	o_val <= 16'b0111111000111001;
            14'h3936 	:	o_val <= 16'b0111111000111010;
            14'h3937 	:	o_val <= 16'b0111111000111010;
            14'h3938 	:	o_val <= 16'b0111111000111011;
            14'h3939 	:	o_val <= 16'b0111111000111011;
            14'h393a 	:	o_val <= 16'b0111111000111100;
            14'h393b 	:	o_val <= 16'b0111111000111101;
            14'h393c 	:	o_val <= 16'b0111111000111101;
            14'h393d 	:	o_val <= 16'b0111111000111110;
            14'h393e 	:	o_val <= 16'b0111111000111110;
            14'h393f 	:	o_val <= 16'b0111111000111111;
            14'h3940 	:	o_val <= 16'b0111111000111111;
            14'h3941 	:	o_val <= 16'b0111111001000000;
            14'h3942 	:	o_val <= 16'b0111111001000000;
            14'h3943 	:	o_val <= 16'b0111111001000001;
            14'h3944 	:	o_val <= 16'b0111111001000001;
            14'h3945 	:	o_val <= 16'b0111111001000010;
            14'h3946 	:	o_val <= 16'b0111111001000010;
            14'h3947 	:	o_val <= 16'b0111111001000011;
            14'h3948 	:	o_val <= 16'b0111111001000011;
            14'h3949 	:	o_val <= 16'b0111111001000100;
            14'h394a 	:	o_val <= 16'b0111111001000100;
            14'h394b 	:	o_val <= 16'b0111111001000101;
            14'h394c 	:	o_val <= 16'b0111111001000101;
            14'h394d 	:	o_val <= 16'b0111111001000110;
            14'h394e 	:	o_val <= 16'b0111111001000110;
            14'h394f 	:	o_val <= 16'b0111111001000111;
            14'h3950 	:	o_val <= 16'b0111111001000111;
            14'h3951 	:	o_val <= 16'b0111111001001000;
            14'h3952 	:	o_val <= 16'b0111111001001000;
            14'h3953 	:	o_val <= 16'b0111111001001001;
            14'h3954 	:	o_val <= 16'b0111111001001001;
            14'h3955 	:	o_val <= 16'b0111111001001010;
            14'h3956 	:	o_val <= 16'b0111111001001010;
            14'h3957 	:	o_val <= 16'b0111111001001011;
            14'h3958 	:	o_val <= 16'b0111111001001011;
            14'h3959 	:	o_val <= 16'b0111111001001100;
            14'h395a 	:	o_val <= 16'b0111111001001100;
            14'h395b 	:	o_val <= 16'b0111111001001101;
            14'h395c 	:	o_val <= 16'b0111111001001101;
            14'h395d 	:	o_val <= 16'b0111111001001110;
            14'h395e 	:	o_val <= 16'b0111111001001111;
            14'h395f 	:	o_val <= 16'b0111111001001111;
            14'h3960 	:	o_val <= 16'b0111111001010000;
            14'h3961 	:	o_val <= 16'b0111111001010000;
            14'h3962 	:	o_val <= 16'b0111111001010001;
            14'h3963 	:	o_val <= 16'b0111111001010001;
            14'h3964 	:	o_val <= 16'b0111111001010010;
            14'h3965 	:	o_val <= 16'b0111111001010010;
            14'h3966 	:	o_val <= 16'b0111111001010011;
            14'h3967 	:	o_val <= 16'b0111111001010011;
            14'h3968 	:	o_val <= 16'b0111111001010100;
            14'h3969 	:	o_val <= 16'b0111111001010100;
            14'h396a 	:	o_val <= 16'b0111111001010101;
            14'h396b 	:	o_val <= 16'b0111111001010101;
            14'h396c 	:	o_val <= 16'b0111111001010110;
            14'h396d 	:	o_val <= 16'b0111111001010110;
            14'h396e 	:	o_val <= 16'b0111111001010111;
            14'h396f 	:	o_val <= 16'b0111111001010111;
            14'h3970 	:	o_val <= 16'b0111111001011000;
            14'h3971 	:	o_val <= 16'b0111111001011000;
            14'h3972 	:	o_val <= 16'b0111111001011001;
            14'h3973 	:	o_val <= 16'b0111111001011001;
            14'h3974 	:	o_val <= 16'b0111111001011010;
            14'h3975 	:	o_val <= 16'b0111111001011010;
            14'h3976 	:	o_val <= 16'b0111111001011011;
            14'h3977 	:	o_val <= 16'b0111111001011011;
            14'h3978 	:	o_val <= 16'b0111111001011100;
            14'h3979 	:	o_val <= 16'b0111111001011100;
            14'h397a 	:	o_val <= 16'b0111111001011101;
            14'h397b 	:	o_val <= 16'b0111111001011101;
            14'h397c 	:	o_val <= 16'b0111111001011110;
            14'h397d 	:	o_val <= 16'b0111111001011110;
            14'h397e 	:	o_val <= 16'b0111111001011111;
            14'h397f 	:	o_val <= 16'b0111111001011111;
            14'h3980 	:	o_val <= 16'b0111111001100000;
            14'h3981 	:	o_val <= 16'b0111111001100000;
            14'h3982 	:	o_val <= 16'b0111111001100001;
            14'h3983 	:	o_val <= 16'b0111111001100001;
            14'h3984 	:	o_val <= 16'b0111111001100010;
            14'h3985 	:	o_val <= 16'b0111111001100010;
            14'h3986 	:	o_val <= 16'b0111111001100011;
            14'h3987 	:	o_val <= 16'b0111111001100011;
            14'h3988 	:	o_val <= 16'b0111111001100100;
            14'h3989 	:	o_val <= 16'b0111111001100100;
            14'h398a 	:	o_val <= 16'b0111111001100101;
            14'h398b 	:	o_val <= 16'b0111111001100101;
            14'h398c 	:	o_val <= 16'b0111111001100110;
            14'h398d 	:	o_val <= 16'b0111111001100110;
            14'h398e 	:	o_val <= 16'b0111111001100111;
            14'h398f 	:	o_val <= 16'b0111111001100111;
            14'h3990 	:	o_val <= 16'b0111111001101000;
            14'h3991 	:	o_val <= 16'b0111111001101000;
            14'h3992 	:	o_val <= 16'b0111111001101001;
            14'h3993 	:	o_val <= 16'b0111111001101001;
            14'h3994 	:	o_val <= 16'b0111111001101010;
            14'h3995 	:	o_val <= 16'b0111111001101010;
            14'h3996 	:	o_val <= 16'b0111111001101011;
            14'h3997 	:	o_val <= 16'b0111111001101011;
            14'h3998 	:	o_val <= 16'b0111111001101100;
            14'h3999 	:	o_val <= 16'b0111111001101100;
            14'h399a 	:	o_val <= 16'b0111111001101101;
            14'h399b 	:	o_val <= 16'b0111111001101101;
            14'h399c 	:	o_val <= 16'b0111111001101101;
            14'h399d 	:	o_val <= 16'b0111111001101110;
            14'h399e 	:	o_val <= 16'b0111111001101110;
            14'h399f 	:	o_val <= 16'b0111111001101111;
            14'h39a0 	:	o_val <= 16'b0111111001101111;
            14'h39a1 	:	o_val <= 16'b0111111001110000;
            14'h39a2 	:	o_val <= 16'b0111111001110000;
            14'h39a3 	:	o_val <= 16'b0111111001110001;
            14'h39a4 	:	o_val <= 16'b0111111001110001;
            14'h39a5 	:	o_val <= 16'b0111111001110010;
            14'h39a6 	:	o_val <= 16'b0111111001110010;
            14'h39a7 	:	o_val <= 16'b0111111001110011;
            14'h39a8 	:	o_val <= 16'b0111111001110011;
            14'h39a9 	:	o_val <= 16'b0111111001110100;
            14'h39aa 	:	o_val <= 16'b0111111001110100;
            14'h39ab 	:	o_val <= 16'b0111111001110101;
            14'h39ac 	:	o_val <= 16'b0111111001110101;
            14'h39ad 	:	o_val <= 16'b0111111001110110;
            14'h39ae 	:	o_val <= 16'b0111111001110110;
            14'h39af 	:	o_val <= 16'b0111111001110111;
            14'h39b0 	:	o_val <= 16'b0111111001110111;
            14'h39b1 	:	o_val <= 16'b0111111001111000;
            14'h39b2 	:	o_val <= 16'b0111111001111000;
            14'h39b3 	:	o_val <= 16'b0111111001111001;
            14'h39b4 	:	o_val <= 16'b0111111001111001;
            14'h39b5 	:	o_val <= 16'b0111111001111010;
            14'h39b6 	:	o_val <= 16'b0111111001111010;
            14'h39b7 	:	o_val <= 16'b0111111001111011;
            14'h39b8 	:	o_val <= 16'b0111111001111011;
            14'h39b9 	:	o_val <= 16'b0111111001111100;
            14'h39ba 	:	o_val <= 16'b0111111001111100;
            14'h39bb 	:	o_val <= 16'b0111111001111101;
            14'h39bc 	:	o_val <= 16'b0111111001111101;
            14'h39bd 	:	o_val <= 16'b0111111001111110;
            14'h39be 	:	o_val <= 16'b0111111001111110;
            14'h39bf 	:	o_val <= 16'b0111111001111110;
            14'h39c0 	:	o_val <= 16'b0111111001111111;
            14'h39c1 	:	o_val <= 16'b0111111001111111;
            14'h39c2 	:	o_val <= 16'b0111111010000000;
            14'h39c3 	:	o_val <= 16'b0111111010000000;
            14'h39c4 	:	o_val <= 16'b0111111010000001;
            14'h39c5 	:	o_val <= 16'b0111111010000001;
            14'h39c6 	:	o_val <= 16'b0111111010000010;
            14'h39c7 	:	o_val <= 16'b0111111010000010;
            14'h39c8 	:	o_val <= 16'b0111111010000011;
            14'h39c9 	:	o_val <= 16'b0111111010000011;
            14'h39ca 	:	o_val <= 16'b0111111010000100;
            14'h39cb 	:	o_val <= 16'b0111111010000100;
            14'h39cc 	:	o_val <= 16'b0111111010000101;
            14'h39cd 	:	o_val <= 16'b0111111010000101;
            14'h39ce 	:	o_val <= 16'b0111111010000110;
            14'h39cf 	:	o_val <= 16'b0111111010000110;
            14'h39d0 	:	o_val <= 16'b0111111010000111;
            14'h39d1 	:	o_val <= 16'b0111111010000111;
            14'h39d2 	:	o_val <= 16'b0111111010001000;
            14'h39d3 	:	o_val <= 16'b0111111010001000;
            14'h39d4 	:	o_val <= 16'b0111111010001001;
            14'h39d5 	:	o_val <= 16'b0111111010001001;
            14'h39d6 	:	o_val <= 16'b0111111010001001;
            14'h39d7 	:	o_val <= 16'b0111111010001010;
            14'h39d8 	:	o_val <= 16'b0111111010001010;
            14'h39d9 	:	o_val <= 16'b0111111010001011;
            14'h39da 	:	o_val <= 16'b0111111010001011;
            14'h39db 	:	o_val <= 16'b0111111010001100;
            14'h39dc 	:	o_val <= 16'b0111111010001100;
            14'h39dd 	:	o_val <= 16'b0111111010001101;
            14'h39de 	:	o_val <= 16'b0111111010001101;
            14'h39df 	:	o_val <= 16'b0111111010001110;
            14'h39e0 	:	o_val <= 16'b0111111010001110;
            14'h39e1 	:	o_val <= 16'b0111111010001111;
            14'h39e2 	:	o_val <= 16'b0111111010001111;
            14'h39e3 	:	o_val <= 16'b0111111010010000;
            14'h39e4 	:	o_val <= 16'b0111111010010000;
            14'h39e5 	:	o_val <= 16'b0111111010010001;
            14'h39e6 	:	o_val <= 16'b0111111010010001;
            14'h39e7 	:	o_val <= 16'b0111111010010001;
            14'h39e8 	:	o_val <= 16'b0111111010010010;
            14'h39e9 	:	o_val <= 16'b0111111010010010;
            14'h39ea 	:	o_val <= 16'b0111111010010011;
            14'h39eb 	:	o_val <= 16'b0111111010010011;
            14'h39ec 	:	o_val <= 16'b0111111010010100;
            14'h39ed 	:	o_val <= 16'b0111111010010100;
            14'h39ee 	:	o_val <= 16'b0111111010010101;
            14'h39ef 	:	o_val <= 16'b0111111010010101;
            14'h39f0 	:	o_val <= 16'b0111111010010110;
            14'h39f1 	:	o_val <= 16'b0111111010010110;
            14'h39f2 	:	o_val <= 16'b0111111010010111;
            14'h39f3 	:	o_val <= 16'b0111111010010111;
            14'h39f4 	:	o_val <= 16'b0111111010011000;
            14'h39f5 	:	o_val <= 16'b0111111010011000;
            14'h39f6 	:	o_val <= 16'b0111111010011000;
            14'h39f7 	:	o_val <= 16'b0111111010011001;
            14'h39f8 	:	o_val <= 16'b0111111010011001;
            14'h39f9 	:	o_val <= 16'b0111111010011010;
            14'h39fa 	:	o_val <= 16'b0111111010011010;
            14'h39fb 	:	o_val <= 16'b0111111010011011;
            14'h39fc 	:	o_val <= 16'b0111111010011011;
            14'h39fd 	:	o_val <= 16'b0111111010011100;
            14'h39fe 	:	o_val <= 16'b0111111010011100;
            14'h39ff 	:	o_val <= 16'b0111111010011101;
            14'h3a00 	:	o_val <= 16'b0111111010011101;
            14'h3a01 	:	o_val <= 16'b0111111010011110;
            14'h3a02 	:	o_val <= 16'b0111111010011110;
            14'h3a03 	:	o_val <= 16'b0111111010011110;
            14'h3a04 	:	o_val <= 16'b0111111010011111;
            14'h3a05 	:	o_val <= 16'b0111111010011111;
            14'h3a06 	:	o_val <= 16'b0111111010100000;
            14'h3a07 	:	o_val <= 16'b0111111010100000;
            14'h3a08 	:	o_val <= 16'b0111111010100001;
            14'h3a09 	:	o_val <= 16'b0111111010100001;
            14'h3a0a 	:	o_val <= 16'b0111111010100010;
            14'h3a0b 	:	o_val <= 16'b0111111010100010;
            14'h3a0c 	:	o_val <= 16'b0111111010100011;
            14'h3a0d 	:	o_val <= 16'b0111111010100011;
            14'h3a0e 	:	o_val <= 16'b0111111010100011;
            14'h3a0f 	:	o_val <= 16'b0111111010100100;
            14'h3a10 	:	o_val <= 16'b0111111010100100;
            14'h3a11 	:	o_val <= 16'b0111111010100101;
            14'h3a12 	:	o_val <= 16'b0111111010100101;
            14'h3a13 	:	o_val <= 16'b0111111010100110;
            14'h3a14 	:	o_val <= 16'b0111111010100110;
            14'h3a15 	:	o_val <= 16'b0111111010100111;
            14'h3a16 	:	o_val <= 16'b0111111010100111;
            14'h3a17 	:	o_val <= 16'b0111111010101000;
            14'h3a18 	:	o_val <= 16'b0111111010101000;
            14'h3a19 	:	o_val <= 16'b0111111010101000;
            14'h3a1a 	:	o_val <= 16'b0111111010101001;
            14'h3a1b 	:	o_val <= 16'b0111111010101001;
            14'h3a1c 	:	o_val <= 16'b0111111010101010;
            14'h3a1d 	:	o_val <= 16'b0111111010101010;
            14'h3a1e 	:	o_val <= 16'b0111111010101011;
            14'h3a1f 	:	o_val <= 16'b0111111010101011;
            14'h3a20 	:	o_val <= 16'b0111111010101100;
            14'h3a21 	:	o_val <= 16'b0111111010101100;
            14'h3a22 	:	o_val <= 16'b0111111010101101;
            14'h3a23 	:	o_val <= 16'b0111111010101101;
            14'h3a24 	:	o_val <= 16'b0111111010101101;
            14'h3a25 	:	o_val <= 16'b0111111010101110;
            14'h3a26 	:	o_val <= 16'b0111111010101110;
            14'h3a27 	:	o_val <= 16'b0111111010101111;
            14'h3a28 	:	o_val <= 16'b0111111010101111;
            14'h3a29 	:	o_val <= 16'b0111111010110000;
            14'h3a2a 	:	o_val <= 16'b0111111010110000;
            14'h3a2b 	:	o_val <= 16'b0111111010110001;
            14'h3a2c 	:	o_val <= 16'b0111111010110001;
            14'h3a2d 	:	o_val <= 16'b0111111010110010;
            14'h3a2e 	:	o_val <= 16'b0111111010110010;
            14'h3a2f 	:	o_val <= 16'b0111111010110010;
            14'h3a30 	:	o_val <= 16'b0111111010110011;
            14'h3a31 	:	o_val <= 16'b0111111010110011;
            14'h3a32 	:	o_val <= 16'b0111111010110100;
            14'h3a33 	:	o_val <= 16'b0111111010110100;
            14'h3a34 	:	o_val <= 16'b0111111010110101;
            14'h3a35 	:	o_val <= 16'b0111111010110101;
            14'h3a36 	:	o_val <= 16'b0111111010110110;
            14'h3a37 	:	o_val <= 16'b0111111010110110;
            14'h3a38 	:	o_val <= 16'b0111111010110110;
            14'h3a39 	:	o_val <= 16'b0111111010110111;
            14'h3a3a 	:	o_val <= 16'b0111111010110111;
            14'h3a3b 	:	o_val <= 16'b0111111010111000;
            14'h3a3c 	:	o_val <= 16'b0111111010111000;
            14'h3a3d 	:	o_val <= 16'b0111111010111001;
            14'h3a3e 	:	o_val <= 16'b0111111010111001;
            14'h3a3f 	:	o_val <= 16'b0111111010111010;
            14'h3a40 	:	o_val <= 16'b0111111010111010;
            14'h3a41 	:	o_val <= 16'b0111111010111010;
            14'h3a42 	:	o_val <= 16'b0111111010111011;
            14'h3a43 	:	o_val <= 16'b0111111010111011;
            14'h3a44 	:	o_val <= 16'b0111111010111100;
            14'h3a45 	:	o_val <= 16'b0111111010111100;
            14'h3a46 	:	o_val <= 16'b0111111010111101;
            14'h3a47 	:	o_val <= 16'b0111111010111101;
            14'h3a48 	:	o_val <= 16'b0111111010111101;
            14'h3a49 	:	o_val <= 16'b0111111010111110;
            14'h3a4a 	:	o_val <= 16'b0111111010111110;
            14'h3a4b 	:	o_val <= 16'b0111111010111111;
            14'h3a4c 	:	o_val <= 16'b0111111010111111;
            14'h3a4d 	:	o_val <= 16'b0111111011000000;
            14'h3a4e 	:	o_val <= 16'b0111111011000000;
            14'h3a4f 	:	o_val <= 16'b0111111011000001;
            14'h3a50 	:	o_val <= 16'b0111111011000001;
            14'h3a51 	:	o_val <= 16'b0111111011000001;
            14'h3a52 	:	o_val <= 16'b0111111011000010;
            14'h3a53 	:	o_val <= 16'b0111111011000010;
            14'h3a54 	:	o_val <= 16'b0111111011000011;
            14'h3a55 	:	o_val <= 16'b0111111011000011;
            14'h3a56 	:	o_val <= 16'b0111111011000100;
            14'h3a57 	:	o_val <= 16'b0111111011000100;
            14'h3a58 	:	o_val <= 16'b0111111011000100;
            14'h3a59 	:	o_val <= 16'b0111111011000101;
            14'h3a5a 	:	o_val <= 16'b0111111011000101;
            14'h3a5b 	:	o_val <= 16'b0111111011000110;
            14'h3a5c 	:	o_val <= 16'b0111111011000110;
            14'h3a5d 	:	o_val <= 16'b0111111011000111;
            14'h3a5e 	:	o_val <= 16'b0111111011000111;
            14'h3a5f 	:	o_val <= 16'b0111111011000111;
            14'h3a60 	:	o_val <= 16'b0111111011001000;
            14'h3a61 	:	o_val <= 16'b0111111011001000;
            14'h3a62 	:	o_val <= 16'b0111111011001001;
            14'h3a63 	:	o_val <= 16'b0111111011001001;
            14'h3a64 	:	o_val <= 16'b0111111011001010;
            14'h3a65 	:	o_val <= 16'b0111111011001010;
            14'h3a66 	:	o_val <= 16'b0111111011001011;
            14'h3a67 	:	o_val <= 16'b0111111011001011;
            14'h3a68 	:	o_val <= 16'b0111111011001011;
            14'h3a69 	:	o_val <= 16'b0111111011001100;
            14'h3a6a 	:	o_val <= 16'b0111111011001100;
            14'h3a6b 	:	o_val <= 16'b0111111011001101;
            14'h3a6c 	:	o_val <= 16'b0111111011001101;
            14'h3a6d 	:	o_val <= 16'b0111111011001110;
            14'h3a6e 	:	o_val <= 16'b0111111011001110;
            14'h3a6f 	:	o_val <= 16'b0111111011001110;
            14'h3a70 	:	o_val <= 16'b0111111011001111;
            14'h3a71 	:	o_val <= 16'b0111111011001111;
            14'h3a72 	:	o_val <= 16'b0111111011010000;
            14'h3a73 	:	o_val <= 16'b0111111011010000;
            14'h3a74 	:	o_val <= 16'b0111111011010001;
            14'h3a75 	:	o_val <= 16'b0111111011010001;
            14'h3a76 	:	o_val <= 16'b0111111011010001;
            14'h3a77 	:	o_val <= 16'b0111111011010010;
            14'h3a78 	:	o_val <= 16'b0111111011010010;
            14'h3a79 	:	o_val <= 16'b0111111011010011;
            14'h3a7a 	:	o_val <= 16'b0111111011010011;
            14'h3a7b 	:	o_val <= 16'b0111111011010011;
            14'h3a7c 	:	o_val <= 16'b0111111011010100;
            14'h3a7d 	:	o_val <= 16'b0111111011010100;
            14'h3a7e 	:	o_val <= 16'b0111111011010101;
            14'h3a7f 	:	o_val <= 16'b0111111011010101;
            14'h3a80 	:	o_val <= 16'b0111111011010110;
            14'h3a81 	:	o_val <= 16'b0111111011010110;
            14'h3a82 	:	o_val <= 16'b0111111011010110;
            14'h3a83 	:	o_val <= 16'b0111111011010111;
            14'h3a84 	:	o_val <= 16'b0111111011010111;
            14'h3a85 	:	o_val <= 16'b0111111011011000;
            14'h3a86 	:	o_val <= 16'b0111111011011000;
            14'h3a87 	:	o_val <= 16'b0111111011011001;
            14'h3a88 	:	o_val <= 16'b0111111011011001;
            14'h3a89 	:	o_val <= 16'b0111111011011001;
            14'h3a8a 	:	o_val <= 16'b0111111011011010;
            14'h3a8b 	:	o_val <= 16'b0111111011011010;
            14'h3a8c 	:	o_val <= 16'b0111111011011011;
            14'h3a8d 	:	o_val <= 16'b0111111011011011;
            14'h3a8e 	:	o_val <= 16'b0111111011011011;
            14'h3a8f 	:	o_val <= 16'b0111111011011100;
            14'h3a90 	:	o_val <= 16'b0111111011011100;
            14'h3a91 	:	o_val <= 16'b0111111011011101;
            14'h3a92 	:	o_val <= 16'b0111111011011101;
            14'h3a93 	:	o_val <= 16'b0111111011011110;
            14'h3a94 	:	o_val <= 16'b0111111011011110;
            14'h3a95 	:	o_val <= 16'b0111111011011110;
            14'h3a96 	:	o_val <= 16'b0111111011011111;
            14'h3a97 	:	o_val <= 16'b0111111011011111;
            14'h3a98 	:	o_val <= 16'b0111111011100000;
            14'h3a99 	:	o_val <= 16'b0111111011100000;
            14'h3a9a 	:	o_val <= 16'b0111111011100000;
            14'h3a9b 	:	o_val <= 16'b0111111011100001;
            14'h3a9c 	:	o_val <= 16'b0111111011100001;
            14'h3a9d 	:	o_val <= 16'b0111111011100010;
            14'h3a9e 	:	o_val <= 16'b0111111011100010;
            14'h3a9f 	:	o_val <= 16'b0111111011100011;
            14'h3aa0 	:	o_val <= 16'b0111111011100011;
            14'h3aa1 	:	o_val <= 16'b0111111011100011;
            14'h3aa2 	:	o_val <= 16'b0111111011100100;
            14'h3aa3 	:	o_val <= 16'b0111111011100100;
            14'h3aa4 	:	o_val <= 16'b0111111011100101;
            14'h3aa5 	:	o_val <= 16'b0111111011100101;
            14'h3aa6 	:	o_val <= 16'b0111111011100101;
            14'h3aa7 	:	o_val <= 16'b0111111011100110;
            14'h3aa8 	:	o_val <= 16'b0111111011100110;
            14'h3aa9 	:	o_val <= 16'b0111111011100111;
            14'h3aaa 	:	o_val <= 16'b0111111011100111;
            14'h3aab 	:	o_val <= 16'b0111111011101000;
            14'h3aac 	:	o_val <= 16'b0111111011101000;
            14'h3aad 	:	o_val <= 16'b0111111011101000;
            14'h3aae 	:	o_val <= 16'b0111111011101001;
            14'h3aaf 	:	o_val <= 16'b0111111011101001;
            14'h3ab0 	:	o_val <= 16'b0111111011101010;
            14'h3ab1 	:	o_val <= 16'b0111111011101010;
            14'h3ab2 	:	o_val <= 16'b0111111011101010;
            14'h3ab3 	:	o_val <= 16'b0111111011101011;
            14'h3ab4 	:	o_val <= 16'b0111111011101011;
            14'h3ab5 	:	o_val <= 16'b0111111011101100;
            14'h3ab6 	:	o_val <= 16'b0111111011101100;
            14'h3ab7 	:	o_val <= 16'b0111111011101100;
            14'h3ab8 	:	o_val <= 16'b0111111011101101;
            14'h3ab9 	:	o_val <= 16'b0111111011101101;
            14'h3aba 	:	o_val <= 16'b0111111011101110;
            14'h3abb 	:	o_val <= 16'b0111111011101110;
            14'h3abc 	:	o_val <= 16'b0111111011101110;
            14'h3abd 	:	o_val <= 16'b0111111011101111;
            14'h3abe 	:	o_val <= 16'b0111111011101111;
            14'h3abf 	:	o_val <= 16'b0111111011110000;
            14'h3ac0 	:	o_val <= 16'b0111111011110000;
            14'h3ac1 	:	o_val <= 16'b0111111011110000;
            14'h3ac2 	:	o_val <= 16'b0111111011110001;
            14'h3ac3 	:	o_val <= 16'b0111111011110001;
            14'h3ac4 	:	o_val <= 16'b0111111011110010;
            14'h3ac5 	:	o_val <= 16'b0111111011110010;
            14'h3ac6 	:	o_val <= 16'b0111111011110010;
            14'h3ac7 	:	o_val <= 16'b0111111011110011;
            14'h3ac8 	:	o_val <= 16'b0111111011110011;
            14'h3ac9 	:	o_val <= 16'b0111111011110100;
            14'h3aca 	:	o_val <= 16'b0111111011110100;
            14'h3acb 	:	o_val <= 16'b0111111011110100;
            14'h3acc 	:	o_val <= 16'b0111111011110101;
            14'h3acd 	:	o_val <= 16'b0111111011110101;
            14'h3ace 	:	o_val <= 16'b0111111011110110;
            14'h3acf 	:	o_val <= 16'b0111111011110110;
            14'h3ad0 	:	o_val <= 16'b0111111011110110;
            14'h3ad1 	:	o_val <= 16'b0111111011110111;
            14'h3ad2 	:	o_val <= 16'b0111111011110111;
            14'h3ad3 	:	o_val <= 16'b0111111011111000;
            14'h3ad4 	:	o_val <= 16'b0111111011111000;
            14'h3ad5 	:	o_val <= 16'b0111111011111000;
            14'h3ad6 	:	o_val <= 16'b0111111011111001;
            14'h3ad7 	:	o_val <= 16'b0111111011111001;
            14'h3ad8 	:	o_val <= 16'b0111111011111010;
            14'h3ad9 	:	o_val <= 16'b0111111011111010;
            14'h3ada 	:	o_val <= 16'b0111111011111010;
            14'h3adb 	:	o_val <= 16'b0111111011111011;
            14'h3adc 	:	o_val <= 16'b0111111011111011;
            14'h3add 	:	o_val <= 16'b0111111011111100;
            14'h3ade 	:	o_val <= 16'b0111111011111100;
            14'h3adf 	:	o_val <= 16'b0111111011111100;
            14'h3ae0 	:	o_val <= 16'b0111111011111101;
            14'h3ae1 	:	o_val <= 16'b0111111011111101;
            14'h3ae2 	:	o_val <= 16'b0111111011111110;
            14'h3ae3 	:	o_val <= 16'b0111111011111110;
            14'h3ae4 	:	o_val <= 16'b0111111011111110;
            14'h3ae5 	:	o_val <= 16'b0111111011111111;
            14'h3ae6 	:	o_val <= 16'b0111111011111111;
            14'h3ae7 	:	o_val <= 16'b0111111100000000;
            14'h3ae8 	:	o_val <= 16'b0111111100000000;
            14'h3ae9 	:	o_val <= 16'b0111111100000000;
            14'h3aea 	:	o_val <= 16'b0111111100000001;
            14'h3aeb 	:	o_val <= 16'b0111111100000001;
            14'h3aec 	:	o_val <= 16'b0111111100000010;
            14'h3aed 	:	o_val <= 16'b0111111100000010;
            14'h3aee 	:	o_val <= 16'b0111111100000010;
            14'h3aef 	:	o_val <= 16'b0111111100000011;
            14'h3af0 	:	o_val <= 16'b0111111100000011;
            14'h3af1 	:	o_val <= 16'b0111111100000011;
            14'h3af2 	:	o_val <= 16'b0111111100000100;
            14'h3af3 	:	o_val <= 16'b0111111100000100;
            14'h3af4 	:	o_val <= 16'b0111111100000101;
            14'h3af5 	:	o_val <= 16'b0111111100000101;
            14'h3af6 	:	o_val <= 16'b0111111100000101;
            14'h3af7 	:	o_val <= 16'b0111111100000110;
            14'h3af8 	:	o_val <= 16'b0111111100000110;
            14'h3af9 	:	o_val <= 16'b0111111100000111;
            14'h3afa 	:	o_val <= 16'b0111111100000111;
            14'h3afb 	:	o_val <= 16'b0111111100000111;
            14'h3afc 	:	o_val <= 16'b0111111100001000;
            14'h3afd 	:	o_val <= 16'b0111111100001000;
            14'h3afe 	:	o_val <= 16'b0111111100001000;
            14'h3aff 	:	o_val <= 16'b0111111100001001;
            14'h3b00 	:	o_val <= 16'b0111111100001001;
            14'h3b01 	:	o_val <= 16'b0111111100001010;
            14'h3b02 	:	o_val <= 16'b0111111100001010;
            14'h3b03 	:	o_val <= 16'b0111111100001010;
            14'h3b04 	:	o_val <= 16'b0111111100001011;
            14'h3b05 	:	o_val <= 16'b0111111100001011;
            14'h3b06 	:	o_val <= 16'b0111111100001100;
            14'h3b07 	:	o_val <= 16'b0111111100001100;
            14'h3b08 	:	o_val <= 16'b0111111100001100;
            14'h3b09 	:	o_val <= 16'b0111111100001101;
            14'h3b0a 	:	o_val <= 16'b0111111100001101;
            14'h3b0b 	:	o_val <= 16'b0111111100001101;
            14'h3b0c 	:	o_val <= 16'b0111111100001110;
            14'h3b0d 	:	o_val <= 16'b0111111100001110;
            14'h3b0e 	:	o_val <= 16'b0111111100001111;
            14'h3b0f 	:	o_val <= 16'b0111111100001111;
            14'h3b10 	:	o_val <= 16'b0111111100001111;
            14'h3b11 	:	o_val <= 16'b0111111100010000;
            14'h3b12 	:	o_val <= 16'b0111111100010000;
            14'h3b13 	:	o_val <= 16'b0111111100010001;
            14'h3b14 	:	o_val <= 16'b0111111100010001;
            14'h3b15 	:	o_val <= 16'b0111111100010001;
            14'h3b16 	:	o_val <= 16'b0111111100010010;
            14'h3b17 	:	o_val <= 16'b0111111100010010;
            14'h3b18 	:	o_val <= 16'b0111111100010010;
            14'h3b19 	:	o_val <= 16'b0111111100010011;
            14'h3b1a 	:	o_val <= 16'b0111111100010011;
            14'h3b1b 	:	o_val <= 16'b0111111100010100;
            14'h3b1c 	:	o_val <= 16'b0111111100010100;
            14'h3b1d 	:	o_val <= 16'b0111111100010100;
            14'h3b1e 	:	o_val <= 16'b0111111100010101;
            14'h3b1f 	:	o_val <= 16'b0111111100010101;
            14'h3b20 	:	o_val <= 16'b0111111100010101;
            14'h3b21 	:	o_val <= 16'b0111111100010110;
            14'h3b22 	:	o_val <= 16'b0111111100010110;
            14'h3b23 	:	o_val <= 16'b0111111100010111;
            14'h3b24 	:	o_val <= 16'b0111111100010111;
            14'h3b25 	:	o_val <= 16'b0111111100010111;
            14'h3b26 	:	o_val <= 16'b0111111100011000;
            14'h3b27 	:	o_val <= 16'b0111111100011000;
            14'h3b28 	:	o_val <= 16'b0111111100011000;
            14'h3b29 	:	o_val <= 16'b0111111100011001;
            14'h3b2a 	:	o_val <= 16'b0111111100011001;
            14'h3b2b 	:	o_val <= 16'b0111111100011010;
            14'h3b2c 	:	o_val <= 16'b0111111100011010;
            14'h3b2d 	:	o_val <= 16'b0111111100011010;
            14'h3b2e 	:	o_val <= 16'b0111111100011011;
            14'h3b2f 	:	o_val <= 16'b0111111100011011;
            14'h3b30 	:	o_val <= 16'b0111111100011011;
            14'h3b31 	:	o_val <= 16'b0111111100011100;
            14'h3b32 	:	o_val <= 16'b0111111100011100;
            14'h3b33 	:	o_val <= 16'b0111111100011100;
            14'h3b34 	:	o_val <= 16'b0111111100011101;
            14'h3b35 	:	o_val <= 16'b0111111100011101;
            14'h3b36 	:	o_val <= 16'b0111111100011110;
            14'h3b37 	:	o_val <= 16'b0111111100011110;
            14'h3b38 	:	o_val <= 16'b0111111100011110;
            14'h3b39 	:	o_val <= 16'b0111111100011111;
            14'h3b3a 	:	o_val <= 16'b0111111100011111;
            14'h3b3b 	:	o_val <= 16'b0111111100011111;
            14'h3b3c 	:	o_val <= 16'b0111111100100000;
            14'h3b3d 	:	o_val <= 16'b0111111100100000;
            14'h3b3e 	:	o_val <= 16'b0111111100100001;
            14'h3b3f 	:	o_val <= 16'b0111111100100001;
            14'h3b40 	:	o_val <= 16'b0111111100100001;
            14'h3b41 	:	o_val <= 16'b0111111100100010;
            14'h3b42 	:	o_val <= 16'b0111111100100010;
            14'h3b43 	:	o_val <= 16'b0111111100100010;
            14'h3b44 	:	o_val <= 16'b0111111100100011;
            14'h3b45 	:	o_val <= 16'b0111111100100011;
            14'h3b46 	:	o_val <= 16'b0111111100100011;
            14'h3b47 	:	o_val <= 16'b0111111100100100;
            14'h3b48 	:	o_val <= 16'b0111111100100100;
            14'h3b49 	:	o_val <= 16'b0111111100100101;
            14'h3b4a 	:	o_val <= 16'b0111111100100101;
            14'h3b4b 	:	o_val <= 16'b0111111100100101;
            14'h3b4c 	:	o_val <= 16'b0111111100100110;
            14'h3b4d 	:	o_val <= 16'b0111111100100110;
            14'h3b4e 	:	o_val <= 16'b0111111100100110;
            14'h3b4f 	:	o_val <= 16'b0111111100100111;
            14'h3b50 	:	o_val <= 16'b0111111100100111;
            14'h3b51 	:	o_val <= 16'b0111111100100111;
            14'h3b52 	:	o_val <= 16'b0111111100101000;
            14'h3b53 	:	o_val <= 16'b0111111100101000;
            14'h3b54 	:	o_val <= 16'b0111111100101000;
            14'h3b55 	:	o_val <= 16'b0111111100101001;
            14'h3b56 	:	o_val <= 16'b0111111100101001;
            14'h3b57 	:	o_val <= 16'b0111111100101010;
            14'h3b58 	:	o_val <= 16'b0111111100101010;
            14'h3b59 	:	o_val <= 16'b0111111100101010;
            14'h3b5a 	:	o_val <= 16'b0111111100101011;
            14'h3b5b 	:	o_val <= 16'b0111111100101011;
            14'h3b5c 	:	o_val <= 16'b0111111100101011;
            14'h3b5d 	:	o_val <= 16'b0111111100101100;
            14'h3b5e 	:	o_val <= 16'b0111111100101100;
            14'h3b5f 	:	o_val <= 16'b0111111100101100;
            14'h3b60 	:	o_val <= 16'b0111111100101101;
            14'h3b61 	:	o_val <= 16'b0111111100101101;
            14'h3b62 	:	o_val <= 16'b0111111100101101;
            14'h3b63 	:	o_val <= 16'b0111111100101110;
            14'h3b64 	:	o_val <= 16'b0111111100101110;
            14'h3b65 	:	o_val <= 16'b0111111100101111;
            14'h3b66 	:	o_val <= 16'b0111111100101111;
            14'h3b67 	:	o_val <= 16'b0111111100101111;
            14'h3b68 	:	o_val <= 16'b0111111100110000;
            14'h3b69 	:	o_val <= 16'b0111111100110000;
            14'h3b6a 	:	o_val <= 16'b0111111100110000;
            14'h3b6b 	:	o_val <= 16'b0111111100110001;
            14'h3b6c 	:	o_val <= 16'b0111111100110001;
            14'h3b6d 	:	o_val <= 16'b0111111100110001;
            14'h3b6e 	:	o_val <= 16'b0111111100110010;
            14'h3b6f 	:	o_val <= 16'b0111111100110010;
            14'h3b70 	:	o_val <= 16'b0111111100110010;
            14'h3b71 	:	o_val <= 16'b0111111100110011;
            14'h3b72 	:	o_val <= 16'b0111111100110011;
            14'h3b73 	:	o_val <= 16'b0111111100110011;
            14'h3b74 	:	o_val <= 16'b0111111100110100;
            14'h3b75 	:	o_val <= 16'b0111111100110100;
            14'h3b76 	:	o_val <= 16'b0111111100110101;
            14'h3b77 	:	o_val <= 16'b0111111100110101;
            14'h3b78 	:	o_val <= 16'b0111111100110101;
            14'h3b79 	:	o_val <= 16'b0111111100110110;
            14'h3b7a 	:	o_val <= 16'b0111111100110110;
            14'h3b7b 	:	o_val <= 16'b0111111100110110;
            14'h3b7c 	:	o_val <= 16'b0111111100110111;
            14'h3b7d 	:	o_val <= 16'b0111111100110111;
            14'h3b7e 	:	o_val <= 16'b0111111100110111;
            14'h3b7f 	:	o_val <= 16'b0111111100111000;
            14'h3b80 	:	o_val <= 16'b0111111100111000;
            14'h3b81 	:	o_val <= 16'b0111111100111000;
            14'h3b82 	:	o_val <= 16'b0111111100111001;
            14'h3b83 	:	o_val <= 16'b0111111100111001;
            14'h3b84 	:	o_val <= 16'b0111111100111001;
            14'h3b85 	:	o_val <= 16'b0111111100111010;
            14'h3b86 	:	o_val <= 16'b0111111100111010;
            14'h3b87 	:	o_val <= 16'b0111111100111010;
            14'h3b88 	:	o_val <= 16'b0111111100111011;
            14'h3b89 	:	o_val <= 16'b0111111100111011;
            14'h3b8a 	:	o_val <= 16'b0111111100111011;
            14'h3b8b 	:	o_val <= 16'b0111111100111100;
            14'h3b8c 	:	o_val <= 16'b0111111100111100;
            14'h3b8d 	:	o_val <= 16'b0111111100111100;
            14'h3b8e 	:	o_val <= 16'b0111111100111101;
            14'h3b8f 	:	o_val <= 16'b0111111100111101;
            14'h3b90 	:	o_val <= 16'b0111111100111110;
            14'h3b91 	:	o_val <= 16'b0111111100111110;
            14'h3b92 	:	o_val <= 16'b0111111100111110;
            14'h3b93 	:	o_val <= 16'b0111111100111111;
            14'h3b94 	:	o_val <= 16'b0111111100111111;
            14'h3b95 	:	o_val <= 16'b0111111100111111;
            14'h3b96 	:	o_val <= 16'b0111111101000000;
            14'h3b97 	:	o_val <= 16'b0111111101000000;
            14'h3b98 	:	o_val <= 16'b0111111101000000;
            14'h3b99 	:	o_val <= 16'b0111111101000001;
            14'h3b9a 	:	o_val <= 16'b0111111101000001;
            14'h3b9b 	:	o_val <= 16'b0111111101000001;
            14'h3b9c 	:	o_val <= 16'b0111111101000010;
            14'h3b9d 	:	o_val <= 16'b0111111101000010;
            14'h3b9e 	:	o_val <= 16'b0111111101000010;
            14'h3b9f 	:	o_val <= 16'b0111111101000011;
            14'h3ba0 	:	o_val <= 16'b0111111101000011;
            14'h3ba1 	:	o_val <= 16'b0111111101000011;
            14'h3ba2 	:	o_val <= 16'b0111111101000100;
            14'h3ba3 	:	o_val <= 16'b0111111101000100;
            14'h3ba4 	:	o_val <= 16'b0111111101000100;
            14'h3ba5 	:	o_val <= 16'b0111111101000101;
            14'h3ba6 	:	o_val <= 16'b0111111101000101;
            14'h3ba7 	:	o_val <= 16'b0111111101000101;
            14'h3ba8 	:	o_val <= 16'b0111111101000110;
            14'h3ba9 	:	o_val <= 16'b0111111101000110;
            14'h3baa 	:	o_val <= 16'b0111111101000110;
            14'h3bab 	:	o_val <= 16'b0111111101000111;
            14'h3bac 	:	o_val <= 16'b0111111101000111;
            14'h3bad 	:	o_val <= 16'b0111111101000111;
            14'h3bae 	:	o_val <= 16'b0111111101001000;
            14'h3baf 	:	o_val <= 16'b0111111101001000;
            14'h3bb0 	:	o_val <= 16'b0111111101001000;
            14'h3bb1 	:	o_val <= 16'b0111111101001001;
            14'h3bb2 	:	o_val <= 16'b0111111101001001;
            14'h3bb3 	:	o_val <= 16'b0111111101001001;
            14'h3bb4 	:	o_val <= 16'b0111111101001010;
            14'h3bb5 	:	o_val <= 16'b0111111101001010;
            14'h3bb6 	:	o_val <= 16'b0111111101001010;
            14'h3bb7 	:	o_val <= 16'b0111111101001011;
            14'h3bb8 	:	o_val <= 16'b0111111101001011;
            14'h3bb9 	:	o_val <= 16'b0111111101001011;
            14'h3bba 	:	o_val <= 16'b0111111101001100;
            14'h3bbb 	:	o_val <= 16'b0111111101001100;
            14'h3bbc 	:	o_val <= 16'b0111111101001100;
            14'h3bbd 	:	o_val <= 16'b0111111101001101;
            14'h3bbe 	:	o_val <= 16'b0111111101001101;
            14'h3bbf 	:	o_val <= 16'b0111111101001101;
            14'h3bc0 	:	o_val <= 16'b0111111101001110;
            14'h3bc1 	:	o_val <= 16'b0111111101001110;
            14'h3bc2 	:	o_val <= 16'b0111111101001110;
            14'h3bc3 	:	o_val <= 16'b0111111101001111;
            14'h3bc4 	:	o_val <= 16'b0111111101001111;
            14'h3bc5 	:	o_val <= 16'b0111111101001111;
            14'h3bc6 	:	o_val <= 16'b0111111101010000;
            14'h3bc7 	:	o_val <= 16'b0111111101010000;
            14'h3bc8 	:	o_val <= 16'b0111111101010000;
            14'h3bc9 	:	o_val <= 16'b0111111101010000;
            14'h3bca 	:	o_val <= 16'b0111111101010001;
            14'h3bcb 	:	o_val <= 16'b0111111101010001;
            14'h3bcc 	:	o_val <= 16'b0111111101010001;
            14'h3bcd 	:	o_val <= 16'b0111111101010010;
            14'h3bce 	:	o_val <= 16'b0111111101010010;
            14'h3bcf 	:	o_val <= 16'b0111111101010010;
            14'h3bd0 	:	o_val <= 16'b0111111101010011;
            14'h3bd1 	:	o_val <= 16'b0111111101010011;
            14'h3bd2 	:	o_val <= 16'b0111111101010011;
            14'h3bd3 	:	o_val <= 16'b0111111101010100;
            14'h3bd4 	:	o_val <= 16'b0111111101010100;
            14'h3bd5 	:	o_val <= 16'b0111111101010100;
            14'h3bd6 	:	o_val <= 16'b0111111101010101;
            14'h3bd7 	:	o_val <= 16'b0111111101010101;
            14'h3bd8 	:	o_val <= 16'b0111111101010101;
            14'h3bd9 	:	o_val <= 16'b0111111101010110;
            14'h3bda 	:	o_val <= 16'b0111111101010110;
            14'h3bdb 	:	o_val <= 16'b0111111101010110;
            14'h3bdc 	:	o_val <= 16'b0111111101010111;
            14'h3bdd 	:	o_val <= 16'b0111111101010111;
            14'h3bde 	:	o_val <= 16'b0111111101010111;
            14'h3bdf 	:	o_val <= 16'b0111111101011000;
            14'h3be0 	:	o_val <= 16'b0111111101011000;
            14'h3be1 	:	o_val <= 16'b0111111101011000;
            14'h3be2 	:	o_val <= 16'b0111111101011000;
            14'h3be3 	:	o_val <= 16'b0111111101011001;
            14'h3be4 	:	o_val <= 16'b0111111101011001;
            14'h3be5 	:	o_val <= 16'b0111111101011001;
            14'h3be6 	:	o_val <= 16'b0111111101011010;
            14'h3be7 	:	o_val <= 16'b0111111101011010;
            14'h3be8 	:	o_val <= 16'b0111111101011010;
            14'h3be9 	:	o_val <= 16'b0111111101011011;
            14'h3bea 	:	o_val <= 16'b0111111101011011;
            14'h3beb 	:	o_val <= 16'b0111111101011011;
            14'h3bec 	:	o_val <= 16'b0111111101011100;
            14'h3bed 	:	o_val <= 16'b0111111101011100;
            14'h3bee 	:	o_val <= 16'b0111111101011100;
            14'h3bef 	:	o_val <= 16'b0111111101011101;
            14'h3bf0 	:	o_val <= 16'b0111111101011101;
            14'h3bf1 	:	o_val <= 16'b0111111101011101;
            14'h3bf2 	:	o_val <= 16'b0111111101011110;
            14'h3bf3 	:	o_val <= 16'b0111111101011110;
            14'h3bf4 	:	o_val <= 16'b0111111101011110;
            14'h3bf5 	:	o_val <= 16'b0111111101011110;
            14'h3bf6 	:	o_val <= 16'b0111111101011111;
            14'h3bf7 	:	o_val <= 16'b0111111101011111;
            14'h3bf8 	:	o_val <= 16'b0111111101011111;
            14'h3bf9 	:	o_val <= 16'b0111111101100000;
            14'h3bfa 	:	o_val <= 16'b0111111101100000;
            14'h3bfb 	:	o_val <= 16'b0111111101100000;
            14'h3bfc 	:	o_val <= 16'b0111111101100001;
            14'h3bfd 	:	o_val <= 16'b0111111101100001;
            14'h3bfe 	:	o_val <= 16'b0111111101100001;
            14'h3bff 	:	o_val <= 16'b0111111101100010;
            14'h3c00 	:	o_val <= 16'b0111111101100010;
            14'h3c01 	:	o_val <= 16'b0111111101100010;
            14'h3c02 	:	o_val <= 16'b0111111101100010;
            14'h3c03 	:	o_val <= 16'b0111111101100011;
            14'h3c04 	:	o_val <= 16'b0111111101100011;
            14'h3c05 	:	o_val <= 16'b0111111101100011;
            14'h3c06 	:	o_val <= 16'b0111111101100100;
            14'h3c07 	:	o_val <= 16'b0111111101100100;
            14'h3c08 	:	o_val <= 16'b0111111101100100;
            14'h3c09 	:	o_val <= 16'b0111111101100101;
            14'h3c0a 	:	o_val <= 16'b0111111101100101;
            14'h3c0b 	:	o_val <= 16'b0111111101100101;
            14'h3c0c 	:	o_val <= 16'b0111111101100110;
            14'h3c0d 	:	o_val <= 16'b0111111101100110;
            14'h3c0e 	:	o_val <= 16'b0111111101100110;
            14'h3c0f 	:	o_val <= 16'b0111111101100110;
            14'h3c10 	:	o_val <= 16'b0111111101100111;
            14'h3c11 	:	o_val <= 16'b0111111101100111;
            14'h3c12 	:	o_val <= 16'b0111111101100111;
            14'h3c13 	:	o_val <= 16'b0111111101101000;
            14'h3c14 	:	o_val <= 16'b0111111101101000;
            14'h3c15 	:	o_val <= 16'b0111111101101000;
            14'h3c16 	:	o_val <= 16'b0111111101101001;
            14'h3c17 	:	o_val <= 16'b0111111101101001;
            14'h3c18 	:	o_val <= 16'b0111111101101001;
            14'h3c19 	:	o_val <= 16'b0111111101101001;
            14'h3c1a 	:	o_val <= 16'b0111111101101010;
            14'h3c1b 	:	o_val <= 16'b0111111101101010;
            14'h3c1c 	:	o_val <= 16'b0111111101101010;
            14'h3c1d 	:	o_val <= 16'b0111111101101011;
            14'h3c1e 	:	o_val <= 16'b0111111101101011;
            14'h3c1f 	:	o_val <= 16'b0111111101101011;
            14'h3c20 	:	o_val <= 16'b0111111101101100;
            14'h3c21 	:	o_val <= 16'b0111111101101100;
            14'h3c22 	:	o_val <= 16'b0111111101101100;
            14'h3c23 	:	o_val <= 16'b0111111101101100;
            14'h3c24 	:	o_val <= 16'b0111111101101101;
            14'h3c25 	:	o_val <= 16'b0111111101101101;
            14'h3c26 	:	o_val <= 16'b0111111101101101;
            14'h3c27 	:	o_val <= 16'b0111111101101110;
            14'h3c28 	:	o_val <= 16'b0111111101101110;
            14'h3c29 	:	o_val <= 16'b0111111101101110;
            14'h3c2a 	:	o_val <= 16'b0111111101101111;
            14'h3c2b 	:	o_val <= 16'b0111111101101111;
            14'h3c2c 	:	o_val <= 16'b0111111101101111;
            14'h3c2d 	:	o_val <= 16'b0111111101101111;
            14'h3c2e 	:	o_val <= 16'b0111111101110000;
            14'h3c2f 	:	o_val <= 16'b0111111101110000;
            14'h3c30 	:	o_val <= 16'b0111111101110000;
            14'h3c31 	:	o_val <= 16'b0111111101110001;
            14'h3c32 	:	o_val <= 16'b0111111101110001;
            14'h3c33 	:	o_val <= 16'b0111111101110001;
            14'h3c34 	:	o_val <= 16'b0111111101110001;
            14'h3c35 	:	o_val <= 16'b0111111101110010;
            14'h3c36 	:	o_val <= 16'b0111111101110010;
            14'h3c37 	:	o_val <= 16'b0111111101110010;
            14'h3c38 	:	o_val <= 16'b0111111101110011;
            14'h3c39 	:	o_val <= 16'b0111111101110011;
            14'h3c3a 	:	o_val <= 16'b0111111101110011;
            14'h3c3b 	:	o_val <= 16'b0111111101110100;
            14'h3c3c 	:	o_val <= 16'b0111111101110100;
            14'h3c3d 	:	o_val <= 16'b0111111101110100;
            14'h3c3e 	:	o_val <= 16'b0111111101110100;
            14'h3c3f 	:	o_val <= 16'b0111111101110101;
            14'h3c40 	:	o_val <= 16'b0111111101110101;
            14'h3c41 	:	o_val <= 16'b0111111101110101;
            14'h3c42 	:	o_val <= 16'b0111111101110110;
            14'h3c43 	:	o_val <= 16'b0111111101110110;
            14'h3c44 	:	o_val <= 16'b0111111101110110;
            14'h3c45 	:	o_val <= 16'b0111111101110110;
            14'h3c46 	:	o_val <= 16'b0111111101110111;
            14'h3c47 	:	o_val <= 16'b0111111101110111;
            14'h3c48 	:	o_val <= 16'b0111111101110111;
            14'h3c49 	:	o_val <= 16'b0111111101111000;
            14'h3c4a 	:	o_val <= 16'b0111111101111000;
            14'h3c4b 	:	o_val <= 16'b0111111101111000;
            14'h3c4c 	:	o_val <= 16'b0111111101111000;
            14'h3c4d 	:	o_val <= 16'b0111111101111001;
            14'h3c4e 	:	o_val <= 16'b0111111101111001;
            14'h3c4f 	:	o_val <= 16'b0111111101111001;
            14'h3c50 	:	o_val <= 16'b0111111101111010;
            14'h3c51 	:	o_val <= 16'b0111111101111010;
            14'h3c52 	:	o_val <= 16'b0111111101111010;
            14'h3c53 	:	o_val <= 16'b0111111101111010;
            14'h3c54 	:	o_val <= 16'b0111111101111011;
            14'h3c55 	:	o_val <= 16'b0111111101111011;
            14'h3c56 	:	o_val <= 16'b0111111101111011;
            14'h3c57 	:	o_val <= 16'b0111111101111100;
            14'h3c58 	:	o_val <= 16'b0111111101111100;
            14'h3c59 	:	o_val <= 16'b0111111101111100;
            14'h3c5a 	:	o_val <= 16'b0111111101111100;
            14'h3c5b 	:	o_val <= 16'b0111111101111101;
            14'h3c5c 	:	o_val <= 16'b0111111101111101;
            14'h3c5d 	:	o_val <= 16'b0111111101111101;
            14'h3c5e 	:	o_val <= 16'b0111111101111101;
            14'h3c5f 	:	o_val <= 16'b0111111101111110;
            14'h3c60 	:	o_val <= 16'b0111111101111110;
            14'h3c61 	:	o_val <= 16'b0111111101111110;
            14'h3c62 	:	o_val <= 16'b0111111101111111;
            14'h3c63 	:	o_val <= 16'b0111111101111111;
            14'h3c64 	:	o_val <= 16'b0111111101111111;
            14'h3c65 	:	o_val <= 16'b0111111101111111;
            14'h3c66 	:	o_val <= 16'b0111111110000000;
            14'h3c67 	:	o_val <= 16'b0111111110000000;
            14'h3c68 	:	o_val <= 16'b0111111110000000;
            14'h3c69 	:	o_val <= 16'b0111111110000001;
            14'h3c6a 	:	o_val <= 16'b0111111110000001;
            14'h3c6b 	:	o_val <= 16'b0111111110000001;
            14'h3c6c 	:	o_val <= 16'b0111111110000001;
            14'h3c6d 	:	o_val <= 16'b0111111110000010;
            14'h3c6e 	:	o_val <= 16'b0111111110000010;
            14'h3c6f 	:	o_val <= 16'b0111111110000010;
            14'h3c70 	:	o_val <= 16'b0111111110000010;
            14'h3c71 	:	o_val <= 16'b0111111110000011;
            14'h3c72 	:	o_val <= 16'b0111111110000011;
            14'h3c73 	:	o_val <= 16'b0111111110000011;
            14'h3c74 	:	o_val <= 16'b0111111110000100;
            14'h3c75 	:	o_val <= 16'b0111111110000100;
            14'h3c76 	:	o_val <= 16'b0111111110000100;
            14'h3c77 	:	o_val <= 16'b0111111110000100;
            14'h3c78 	:	o_val <= 16'b0111111110000101;
            14'h3c79 	:	o_val <= 16'b0111111110000101;
            14'h3c7a 	:	o_val <= 16'b0111111110000101;
            14'h3c7b 	:	o_val <= 16'b0111111110000101;
            14'h3c7c 	:	o_val <= 16'b0111111110000110;
            14'h3c7d 	:	o_val <= 16'b0111111110000110;
            14'h3c7e 	:	o_val <= 16'b0111111110000110;
            14'h3c7f 	:	o_val <= 16'b0111111110000111;
            14'h3c80 	:	o_val <= 16'b0111111110000111;
            14'h3c81 	:	o_val <= 16'b0111111110000111;
            14'h3c82 	:	o_val <= 16'b0111111110000111;
            14'h3c83 	:	o_val <= 16'b0111111110001000;
            14'h3c84 	:	o_val <= 16'b0111111110001000;
            14'h3c85 	:	o_val <= 16'b0111111110001000;
            14'h3c86 	:	o_val <= 16'b0111111110001000;
            14'h3c87 	:	o_val <= 16'b0111111110001001;
            14'h3c88 	:	o_val <= 16'b0111111110001001;
            14'h3c89 	:	o_val <= 16'b0111111110001001;
            14'h3c8a 	:	o_val <= 16'b0111111110001001;
            14'h3c8b 	:	o_val <= 16'b0111111110001010;
            14'h3c8c 	:	o_val <= 16'b0111111110001010;
            14'h3c8d 	:	o_val <= 16'b0111111110001010;
            14'h3c8e 	:	o_val <= 16'b0111111110001011;
            14'h3c8f 	:	o_val <= 16'b0111111110001011;
            14'h3c90 	:	o_val <= 16'b0111111110001011;
            14'h3c91 	:	o_val <= 16'b0111111110001011;
            14'h3c92 	:	o_val <= 16'b0111111110001100;
            14'h3c93 	:	o_val <= 16'b0111111110001100;
            14'h3c94 	:	o_val <= 16'b0111111110001100;
            14'h3c95 	:	o_val <= 16'b0111111110001100;
            14'h3c96 	:	o_val <= 16'b0111111110001101;
            14'h3c97 	:	o_val <= 16'b0111111110001101;
            14'h3c98 	:	o_val <= 16'b0111111110001101;
            14'h3c99 	:	o_val <= 16'b0111111110001101;
            14'h3c9a 	:	o_val <= 16'b0111111110001110;
            14'h3c9b 	:	o_val <= 16'b0111111110001110;
            14'h3c9c 	:	o_val <= 16'b0111111110001110;
            14'h3c9d 	:	o_val <= 16'b0111111110001110;
            14'h3c9e 	:	o_val <= 16'b0111111110001111;
            14'h3c9f 	:	o_val <= 16'b0111111110001111;
            14'h3ca0 	:	o_val <= 16'b0111111110001111;
            14'h3ca1 	:	o_val <= 16'b0111111110010000;
            14'h3ca2 	:	o_val <= 16'b0111111110010000;
            14'h3ca3 	:	o_val <= 16'b0111111110010000;
            14'h3ca4 	:	o_val <= 16'b0111111110010000;
            14'h3ca5 	:	o_val <= 16'b0111111110010001;
            14'h3ca6 	:	o_val <= 16'b0111111110010001;
            14'h3ca7 	:	o_val <= 16'b0111111110010001;
            14'h3ca8 	:	o_val <= 16'b0111111110010001;
            14'h3ca9 	:	o_val <= 16'b0111111110010010;
            14'h3caa 	:	o_val <= 16'b0111111110010010;
            14'h3cab 	:	o_val <= 16'b0111111110010010;
            14'h3cac 	:	o_val <= 16'b0111111110010010;
            14'h3cad 	:	o_val <= 16'b0111111110010011;
            14'h3cae 	:	o_val <= 16'b0111111110010011;
            14'h3caf 	:	o_val <= 16'b0111111110010011;
            14'h3cb0 	:	o_val <= 16'b0111111110010011;
            14'h3cb1 	:	o_val <= 16'b0111111110010100;
            14'h3cb2 	:	o_val <= 16'b0111111110010100;
            14'h3cb3 	:	o_val <= 16'b0111111110010100;
            14'h3cb4 	:	o_val <= 16'b0111111110010100;
            14'h3cb5 	:	o_val <= 16'b0111111110010101;
            14'h3cb6 	:	o_val <= 16'b0111111110010101;
            14'h3cb7 	:	o_val <= 16'b0111111110010101;
            14'h3cb8 	:	o_val <= 16'b0111111110010101;
            14'h3cb9 	:	o_val <= 16'b0111111110010110;
            14'h3cba 	:	o_val <= 16'b0111111110010110;
            14'h3cbb 	:	o_val <= 16'b0111111110010110;
            14'h3cbc 	:	o_val <= 16'b0111111110010110;
            14'h3cbd 	:	o_val <= 16'b0111111110010111;
            14'h3cbe 	:	o_val <= 16'b0111111110010111;
            14'h3cbf 	:	o_val <= 16'b0111111110010111;
            14'h3cc0 	:	o_val <= 16'b0111111110010111;
            14'h3cc1 	:	o_val <= 16'b0111111110011000;
            14'h3cc2 	:	o_val <= 16'b0111111110011000;
            14'h3cc3 	:	o_val <= 16'b0111111110011000;
            14'h3cc4 	:	o_val <= 16'b0111111110011000;
            14'h3cc5 	:	o_val <= 16'b0111111110011001;
            14'h3cc6 	:	o_val <= 16'b0111111110011001;
            14'h3cc7 	:	o_val <= 16'b0111111110011001;
            14'h3cc8 	:	o_val <= 16'b0111111110011001;
            14'h3cc9 	:	o_val <= 16'b0111111110011010;
            14'h3cca 	:	o_val <= 16'b0111111110011010;
            14'h3ccb 	:	o_val <= 16'b0111111110011010;
            14'h3ccc 	:	o_val <= 16'b0111111110011010;
            14'h3ccd 	:	o_val <= 16'b0111111110011011;
            14'h3cce 	:	o_val <= 16'b0111111110011011;
            14'h3ccf 	:	o_val <= 16'b0111111110011011;
            14'h3cd0 	:	o_val <= 16'b0111111110011011;
            14'h3cd1 	:	o_val <= 16'b0111111110011100;
            14'h3cd2 	:	o_val <= 16'b0111111110011100;
            14'h3cd3 	:	o_val <= 16'b0111111110011100;
            14'h3cd4 	:	o_val <= 16'b0111111110011100;
            14'h3cd5 	:	o_val <= 16'b0111111110011101;
            14'h3cd6 	:	o_val <= 16'b0111111110011101;
            14'h3cd7 	:	o_val <= 16'b0111111110011101;
            14'h3cd8 	:	o_val <= 16'b0111111110011101;
            14'h3cd9 	:	o_val <= 16'b0111111110011110;
            14'h3cda 	:	o_val <= 16'b0111111110011110;
            14'h3cdb 	:	o_val <= 16'b0111111110011110;
            14'h3cdc 	:	o_val <= 16'b0111111110011110;
            14'h3cdd 	:	o_val <= 16'b0111111110011111;
            14'h3cde 	:	o_val <= 16'b0111111110011111;
            14'h3cdf 	:	o_val <= 16'b0111111110011111;
            14'h3ce0 	:	o_val <= 16'b0111111110011111;
            14'h3ce1 	:	o_val <= 16'b0111111110100000;
            14'h3ce2 	:	o_val <= 16'b0111111110100000;
            14'h3ce3 	:	o_val <= 16'b0111111110100000;
            14'h3ce4 	:	o_val <= 16'b0111111110100000;
            14'h3ce5 	:	o_val <= 16'b0111111110100000;
            14'h3ce6 	:	o_val <= 16'b0111111110100001;
            14'h3ce7 	:	o_val <= 16'b0111111110100001;
            14'h3ce8 	:	o_val <= 16'b0111111110100001;
            14'h3ce9 	:	o_val <= 16'b0111111110100001;
            14'h3cea 	:	o_val <= 16'b0111111110100010;
            14'h3ceb 	:	o_val <= 16'b0111111110100010;
            14'h3cec 	:	o_val <= 16'b0111111110100010;
            14'h3ced 	:	o_val <= 16'b0111111110100010;
            14'h3cee 	:	o_val <= 16'b0111111110100011;
            14'h3cef 	:	o_val <= 16'b0111111110100011;
            14'h3cf0 	:	o_val <= 16'b0111111110100011;
            14'h3cf1 	:	o_val <= 16'b0111111110100011;
            14'h3cf2 	:	o_val <= 16'b0111111110100100;
            14'h3cf3 	:	o_val <= 16'b0111111110100100;
            14'h3cf4 	:	o_val <= 16'b0111111110100100;
            14'h3cf5 	:	o_val <= 16'b0111111110100100;
            14'h3cf6 	:	o_val <= 16'b0111111110100101;
            14'h3cf7 	:	o_val <= 16'b0111111110100101;
            14'h3cf8 	:	o_val <= 16'b0111111110100101;
            14'h3cf9 	:	o_val <= 16'b0111111110100101;
            14'h3cfa 	:	o_val <= 16'b0111111110100101;
            14'h3cfb 	:	o_val <= 16'b0111111110100110;
            14'h3cfc 	:	o_val <= 16'b0111111110100110;
            14'h3cfd 	:	o_val <= 16'b0111111110100110;
            14'h3cfe 	:	o_val <= 16'b0111111110100110;
            14'h3cff 	:	o_val <= 16'b0111111110100111;
            14'h3d00 	:	o_val <= 16'b0111111110100111;
            14'h3d01 	:	o_val <= 16'b0111111110100111;
            14'h3d02 	:	o_val <= 16'b0111111110100111;
            14'h3d03 	:	o_val <= 16'b0111111110101000;
            14'h3d04 	:	o_val <= 16'b0111111110101000;
            14'h3d05 	:	o_val <= 16'b0111111110101000;
            14'h3d06 	:	o_val <= 16'b0111111110101000;
            14'h3d07 	:	o_val <= 16'b0111111110101000;
            14'h3d08 	:	o_val <= 16'b0111111110101001;
            14'h3d09 	:	o_val <= 16'b0111111110101001;
            14'h3d0a 	:	o_val <= 16'b0111111110101001;
            14'h3d0b 	:	o_val <= 16'b0111111110101001;
            14'h3d0c 	:	o_val <= 16'b0111111110101010;
            14'h3d0d 	:	o_val <= 16'b0111111110101010;
            14'h3d0e 	:	o_val <= 16'b0111111110101010;
            14'h3d0f 	:	o_val <= 16'b0111111110101010;
            14'h3d10 	:	o_val <= 16'b0111111110101010;
            14'h3d11 	:	o_val <= 16'b0111111110101011;
            14'h3d12 	:	o_val <= 16'b0111111110101011;
            14'h3d13 	:	o_val <= 16'b0111111110101011;
            14'h3d14 	:	o_val <= 16'b0111111110101011;
            14'h3d15 	:	o_val <= 16'b0111111110101100;
            14'h3d16 	:	o_val <= 16'b0111111110101100;
            14'h3d17 	:	o_val <= 16'b0111111110101100;
            14'h3d18 	:	o_val <= 16'b0111111110101100;
            14'h3d19 	:	o_val <= 16'b0111111110101101;
            14'h3d1a 	:	o_val <= 16'b0111111110101101;
            14'h3d1b 	:	o_val <= 16'b0111111110101101;
            14'h3d1c 	:	o_val <= 16'b0111111110101101;
            14'h3d1d 	:	o_val <= 16'b0111111110101101;
            14'h3d1e 	:	o_val <= 16'b0111111110101110;
            14'h3d1f 	:	o_val <= 16'b0111111110101110;
            14'h3d20 	:	o_val <= 16'b0111111110101110;
            14'h3d21 	:	o_val <= 16'b0111111110101110;
            14'h3d22 	:	o_val <= 16'b0111111110101111;
            14'h3d23 	:	o_val <= 16'b0111111110101111;
            14'h3d24 	:	o_val <= 16'b0111111110101111;
            14'h3d25 	:	o_val <= 16'b0111111110101111;
            14'h3d26 	:	o_val <= 16'b0111111110101111;
            14'h3d27 	:	o_val <= 16'b0111111110110000;
            14'h3d28 	:	o_val <= 16'b0111111110110000;
            14'h3d29 	:	o_val <= 16'b0111111110110000;
            14'h3d2a 	:	o_val <= 16'b0111111110110000;
            14'h3d2b 	:	o_val <= 16'b0111111110110000;
            14'h3d2c 	:	o_val <= 16'b0111111110110001;
            14'h3d2d 	:	o_val <= 16'b0111111110110001;
            14'h3d2e 	:	o_val <= 16'b0111111110110001;
            14'h3d2f 	:	o_val <= 16'b0111111110110001;
            14'h3d30 	:	o_val <= 16'b0111111110110010;
            14'h3d31 	:	o_val <= 16'b0111111110110010;
            14'h3d32 	:	o_val <= 16'b0111111110110010;
            14'h3d33 	:	o_val <= 16'b0111111110110010;
            14'h3d34 	:	o_val <= 16'b0111111110110010;
            14'h3d35 	:	o_val <= 16'b0111111110110011;
            14'h3d36 	:	o_val <= 16'b0111111110110011;
            14'h3d37 	:	o_val <= 16'b0111111110110011;
            14'h3d38 	:	o_val <= 16'b0111111110110011;
            14'h3d39 	:	o_val <= 16'b0111111110110100;
            14'h3d3a 	:	o_val <= 16'b0111111110110100;
            14'h3d3b 	:	o_val <= 16'b0111111110110100;
            14'h3d3c 	:	o_val <= 16'b0111111110110100;
            14'h3d3d 	:	o_val <= 16'b0111111110110100;
            14'h3d3e 	:	o_val <= 16'b0111111110110101;
            14'h3d3f 	:	o_val <= 16'b0111111110110101;
            14'h3d40 	:	o_val <= 16'b0111111110110101;
            14'h3d41 	:	o_val <= 16'b0111111110110101;
            14'h3d42 	:	o_val <= 16'b0111111110110101;
            14'h3d43 	:	o_val <= 16'b0111111110110110;
            14'h3d44 	:	o_val <= 16'b0111111110110110;
            14'h3d45 	:	o_val <= 16'b0111111110110110;
            14'h3d46 	:	o_val <= 16'b0111111110110110;
            14'h3d47 	:	o_val <= 16'b0111111110110110;
            14'h3d48 	:	o_val <= 16'b0111111110110111;
            14'h3d49 	:	o_val <= 16'b0111111110110111;
            14'h3d4a 	:	o_val <= 16'b0111111110110111;
            14'h3d4b 	:	o_val <= 16'b0111111110110111;
            14'h3d4c 	:	o_val <= 16'b0111111110111000;
            14'h3d4d 	:	o_val <= 16'b0111111110111000;
            14'h3d4e 	:	o_val <= 16'b0111111110111000;
            14'h3d4f 	:	o_val <= 16'b0111111110111000;
            14'h3d50 	:	o_val <= 16'b0111111110111000;
            14'h3d51 	:	o_val <= 16'b0111111110111001;
            14'h3d52 	:	o_val <= 16'b0111111110111001;
            14'h3d53 	:	o_val <= 16'b0111111110111001;
            14'h3d54 	:	o_val <= 16'b0111111110111001;
            14'h3d55 	:	o_val <= 16'b0111111110111001;
            14'h3d56 	:	o_val <= 16'b0111111110111010;
            14'h3d57 	:	o_val <= 16'b0111111110111010;
            14'h3d58 	:	o_val <= 16'b0111111110111010;
            14'h3d59 	:	o_val <= 16'b0111111110111010;
            14'h3d5a 	:	o_val <= 16'b0111111110111010;
            14'h3d5b 	:	o_val <= 16'b0111111110111011;
            14'h3d5c 	:	o_val <= 16'b0111111110111011;
            14'h3d5d 	:	o_val <= 16'b0111111110111011;
            14'h3d5e 	:	o_val <= 16'b0111111110111011;
            14'h3d5f 	:	o_val <= 16'b0111111110111011;
            14'h3d60 	:	o_val <= 16'b0111111110111100;
            14'h3d61 	:	o_val <= 16'b0111111110111100;
            14'h3d62 	:	o_val <= 16'b0111111110111100;
            14'h3d63 	:	o_val <= 16'b0111111110111100;
            14'h3d64 	:	o_val <= 16'b0111111110111100;
            14'h3d65 	:	o_val <= 16'b0111111110111101;
            14'h3d66 	:	o_val <= 16'b0111111110111101;
            14'h3d67 	:	o_val <= 16'b0111111110111101;
            14'h3d68 	:	o_val <= 16'b0111111110111101;
            14'h3d69 	:	o_val <= 16'b0111111110111101;
            14'h3d6a 	:	o_val <= 16'b0111111110111110;
            14'h3d6b 	:	o_val <= 16'b0111111110111110;
            14'h3d6c 	:	o_val <= 16'b0111111110111110;
            14'h3d6d 	:	o_val <= 16'b0111111110111110;
            14'h3d6e 	:	o_val <= 16'b0111111110111110;
            14'h3d6f 	:	o_val <= 16'b0111111110111111;
            14'h3d70 	:	o_val <= 16'b0111111110111111;
            14'h3d71 	:	o_val <= 16'b0111111110111111;
            14'h3d72 	:	o_val <= 16'b0111111110111111;
            14'h3d73 	:	o_val <= 16'b0111111110111111;
            14'h3d74 	:	o_val <= 16'b0111111111000000;
            14'h3d75 	:	o_val <= 16'b0111111111000000;
            14'h3d76 	:	o_val <= 16'b0111111111000000;
            14'h3d77 	:	o_val <= 16'b0111111111000000;
            14'h3d78 	:	o_val <= 16'b0111111111000000;
            14'h3d79 	:	o_val <= 16'b0111111111000001;
            14'h3d7a 	:	o_val <= 16'b0111111111000001;
            14'h3d7b 	:	o_val <= 16'b0111111111000001;
            14'h3d7c 	:	o_val <= 16'b0111111111000001;
            14'h3d7d 	:	o_val <= 16'b0111111111000001;
            14'h3d7e 	:	o_val <= 16'b0111111111000010;
            14'h3d7f 	:	o_val <= 16'b0111111111000010;
            14'h3d80 	:	o_val <= 16'b0111111111000010;
            14'h3d81 	:	o_val <= 16'b0111111111000010;
            14'h3d82 	:	o_val <= 16'b0111111111000010;
            14'h3d83 	:	o_val <= 16'b0111111111000011;
            14'h3d84 	:	o_val <= 16'b0111111111000011;
            14'h3d85 	:	o_val <= 16'b0111111111000011;
            14'h3d86 	:	o_val <= 16'b0111111111000011;
            14'h3d87 	:	o_val <= 16'b0111111111000011;
            14'h3d88 	:	o_val <= 16'b0111111111000011;
            14'h3d89 	:	o_val <= 16'b0111111111000100;
            14'h3d8a 	:	o_val <= 16'b0111111111000100;
            14'h3d8b 	:	o_val <= 16'b0111111111000100;
            14'h3d8c 	:	o_val <= 16'b0111111111000100;
            14'h3d8d 	:	o_val <= 16'b0111111111000100;
            14'h3d8e 	:	o_val <= 16'b0111111111000101;
            14'h3d8f 	:	o_val <= 16'b0111111111000101;
            14'h3d90 	:	o_val <= 16'b0111111111000101;
            14'h3d91 	:	o_val <= 16'b0111111111000101;
            14'h3d92 	:	o_val <= 16'b0111111111000101;
            14'h3d93 	:	o_val <= 16'b0111111111000110;
            14'h3d94 	:	o_val <= 16'b0111111111000110;
            14'h3d95 	:	o_val <= 16'b0111111111000110;
            14'h3d96 	:	o_val <= 16'b0111111111000110;
            14'h3d97 	:	o_val <= 16'b0111111111000110;
            14'h3d98 	:	o_val <= 16'b0111111111000110;
            14'h3d99 	:	o_val <= 16'b0111111111000111;
            14'h3d9a 	:	o_val <= 16'b0111111111000111;
            14'h3d9b 	:	o_val <= 16'b0111111111000111;
            14'h3d9c 	:	o_val <= 16'b0111111111000111;
            14'h3d9d 	:	o_val <= 16'b0111111111000111;
            14'h3d9e 	:	o_val <= 16'b0111111111001000;
            14'h3d9f 	:	o_val <= 16'b0111111111001000;
            14'h3da0 	:	o_val <= 16'b0111111111001000;
            14'h3da1 	:	o_val <= 16'b0111111111001000;
            14'h3da2 	:	o_val <= 16'b0111111111001000;
            14'h3da3 	:	o_val <= 16'b0111111111001000;
            14'h3da4 	:	o_val <= 16'b0111111111001001;
            14'h3da5 	:	o_val <= 16'b0111111111001001;
            14'h3da6 	:	o_val <= 16'b0111111111001001;
            14'h3da7 	:	o_val <= 16'b0111111111001001;
            14'h3da8 	:	o_val <= 16'b0111111111001001;
            14'h3da9 	:	o_val <= 16'b0111111111001010;
            14'h3daa 	:	o_val <= 16'b0111111111001010;
            14'h3dab 	:	o_val <= 16'b0111111111001010;
            14'h3dac 	:	o_val <= 16'b0111111111001010;
            14'h3dad 	:	o_val <= 16'b0111111111001010;
            14'h3dae 	:	o_val <= 16'b0111111111001010;
            14'h3daf 	:	o_val <= 16'b0111111111001011;
            14'h3db0 	:	o_val <= 16'b0111111111001011;
            14'h3db1 	:	o_val <= 16'b0111111111001011;
            14'h3db2 	:	o_val <= 16'b0111111111001011;
            14'h3db3 	:	o_val <= 16'b0111111111001011;
            14'h3db4 	:	o_val <= 16'b0111111111001100;
            14'h3db5 	:	o_val <= 16'b0111111111001100;
            14'h3db6 	:	o_val <= 16'b0111111111001100;
            14'h3db7 	:	o_val <= 16'b0111111111001100;
            14'h3db8 	:	o_val <= 16'b0111111111001100;
            14'h3db9 	:	o_val <= 16'b0111111111001100;
            14'h3dba 	:	o_val <= 16'b0111111111001101;
            14'h3dbb 	:	o_val <= 16'b0111111111001101;
            14'h3dbc 	:	o_val <= 16'b0111111111001101;
            14'h3dbd 	:	o_val <= 16'b0111111111001101;
            14'h3dbe 	:	o_val <= 16'b0111111111001101;
            14'h3dbf 	:	o_val <= 16'b0111111111001101;
            14'h3dc0 	:	o_val <= 16'b0111111111001110;
            14'h3dc1 	:	o_val <= 16'b0111111111001110;
            14'h3dc2 	:	o_val <= 16'b0111111111001110;
            14'h3dc3 	:	o_val <= 16'b0111111111001110;
            14'h3dc4 	:	o_val <= 16'b0111111111001110;
            14'h3dc5 	:	o_val <= 16'b0111111111001110;
            14'h3dc6 	:	o_val <= 16'b0111111111001111;
            14'h3dc7 	:	o_val <= 16'b0111111111001111;
            14'h3dc8 	:	o_val <= 16'b0111111111001111;
            14'h3dc9 	:	o_val <= 16'b0111111111001111;
            14'h3dca 	:	o_val <= 16'b0111111111001111;
            14'h3dcb 	:	o_val <= 16'b0111111111010000;
            14'h3dcc 	:	o_val <= 16'b0111111111010000;
            14'h3dcd 	:	o_val <= 16'b0111111111010000;
            14'h3dce 	:	o_val <= 16'b0111111111010000;
            14'h3dcf 	:	o_val <= 16'b0111111111010000;
            14'h3dd0 	:	o_val <= 16'b0111111111010000;
            14'h3dd1 	:	o_val <= 16'b0111111111010001;
            14'h3dd2 	:	o_val <= 16'b0111111111010001;
            14'h3dd3 	:	o_val <= 16'b0111111111010001;
            14'h3dd4 	:	o_val <= 16'b0111111111010001;
            14'h3dd5 	:	o_val <= 16'b0111111111010001;
            14'h3dd6 	:	o_val <= 16'b0111111111010001;
            14'h3dd7 	:	o_val <= 16'b0111111111010010;
            14'h3dd8 	:	o_val <= 16'b0111111111010010;
            14'h3dd9 	:	o_val <= 16'b0111111111010010;
            14'h3dda 	:	o_val <= 16'b0111111111010010;
            14'h3ddb 	:	o_val <= 16'b0111111111010010;
            14'h3ddc 	:	o_val <= 16'b0111111111010010;
            14'h3ddd 	:	o_val <= 16'b0111111111010011;
            14'h3dde 	:	o_val <= 16'b0111111111010011;
            14'h3ddf 	:	o_val <= 16'b0111111111010011;
            14'h3de0 	:	o_val <= 16'b0111111111010011;
            14'h3de1 	:	o_val <= 16'b0111111111010011;
            14'h3de2 	:	o_val <= 16'b0111111111010011;
            14'h3de3 	:	o_val <= 16'b0111111111010100;
            14'h3de4 	:	o_val <= 16'b0111111111010100;
            14'h3de5 	:	o_val <= 16'b0111111111010100;
            14'h3de6 	:	o_val <= 16'b0111111111010100;
            14'h3de7 	:	o_val <= 16'b0111111111010100;
            14'h3de8 	:	o_val <= 16'b0111111111010100;
            14'h3de9 	:	o_val <= 16'b0111111111010100;
            14'h3dea 	:	o_val <= 16'b0111111111010101;
            14'h3deb 	:	o_val <= 16'b0111111111010101;
            14'h3dec 	:	o_val <= 16'b0111111111010101;
            14'h3ded 	:	o_val <= 16'b0111111111010101;
            14'h3dee 	:	o_val <= 16'b0111111111010101;
            14'h3def 	:	o_val <= 16'b0111111111010101;
            14'h3df0 	:	o_val <= 16'b0111111111010110;
            14'h3df1 	:	o_val <= 16'b0111111111010110;
            14'h3df2 	:	o_val <= 16'b0111111111010110;
            14'h3df3 	:	o_val <= 16'b0111111111010110;
            14'h3df4 	:	o_val <= 16'b0111111111010110;
            14'h3df5 	:	o_val <= 16'b0111111111010110;
            14'h3df6 	:	o_val <= 16'b0111111111010111;
            14'h3df7 	:	o_val <= 16'b0111111111010111;
            14'h3df8 	:	o_val <= 16'b0111111111010111;
            14'h3df9 	:	o_val <= 16'b0111111111010111;
            14'h3dfa 	:	o_val <= 16'b0111111111010111;
            14'h3dfb 	:	o_val <= 16'b0111111111010111;
            14'h3dfc 	:	o_val <= 16'b0111111111010111;
            14'h3dfd 	:	o_val <= 16'b0111111111011000;
            14'h3dfe 	:	o_val <= 16'b0111111111011000;
            14'h3dff 	:	o_val <= 16'b0111111111011000;
            14'h3e00 	:	o_val <= 16'b0111111111011000;
            14'h3e01 	:	o_val <= 16'b0111111111011000;
            14'h3e02 	:	o_val <= 16'b0111111111011000;
            14'h3e03 	:	o_val <= 16'b0111111111011001;
            14'h3e04 	:	o_val <= 16'b0111111111011001;
            14'h3e05 	:	o_val <= 16'b0111111111011001;
            14'h3e06 	:	o_val <= 16'b0111111111011001;
            14'h3e07 	:	o_val <= 16'b0111111111011001;
            14'h3e08 	:	o_val <= 16'b0111111111011001;
            14'h3e09 	:	o_val <= 16'b0111111111011001;
            14'h3e0a 	:	o_val <= 16'b0111111111011010;
            14'h3e0b 	:	o_val <= 16'b0111111111011010;
            14'h3e0c 	:	o_val <= 16'b0111111111011010;
            14'h3e0d 	:	o_val <= 16'b0111111111011010;
            14'h3e0e 	:	o_val <= 16'b0111111111011010;
            14'h3e0f 	:	o_val <= 16'b0111111111011010;
            14'h3e10 	:	o_val <= 16'b0111111111011011;
            14'h3e11 	:	o_val <= 16'b0111111111011011;
            14'h3e12 	:	o_val <= 16'b0111111111011011;
            14'h3e13 	:	o_val <= 16'b0111111111011011;
            14'h3e14 	:	o_val <= 16'b0111111111011011;
            14'h3e15 	:	o_val <= 16'b0111111111011011;
            14'h3e16 	:	o_val <= 16'b0111111111011011;
            14'h3e17 	:	o_val <= 16'b0111111111011100;
            14'h3e18 	:	o_val <= 16'b0111111111011100;
            14'h3e19 	:	o_val <= 16'b0111111111011100;
            14'h3e1a 	:	o_val <= 16'b0111111111011100;
            14'h3e1b 	:	o_val <= 16'b0111111111011100;
            14'h3e1c 	:	o_val <= 16'b0111111111011100;
            14'h3e1d 	:	o_val <= 16'b0111111111011100;
            14'h3e1e 	:	o_val <= 16'b0111111111011101;
            14'h3e1f 	:	o_val <= 16'b0111111111011101;
            14'h3e20 	:	o_val <= 16'b0111111111011101;
            14'h3e21 	:	o_val <= 16'b0111111111011101;
            14'h3e22 	:	o_val <= 16'b0111111111011101;
            14'h3e23 	:	o_val <= 16'b0111111111011101;
            14'h3e24 	:	o_val <= 16'b0111111111011101;
            14'h3e25 	:	o_val <= 16'b0111111111011110;
            14'h3e26 	:	o_val <= 16'b0111111111011110;
            14'h3e27 	:	o_val <= 16'b0111111111011110;
            14'h3e28 	:	o_val <= 16'b0111111111011110;
            14'h3e29 	:	o_val <= 16'b0111111111011110;
            14'h3e2a 	:	o_val <= 16'b0111111111011110;
            14'h3e2b 	:	o_val <= 16'b0111111111011110;
            14'h3e2c 	:	o_val <= 16'b0111111111011111;
            14'h3e2d 	:	o_val <= 16'b0111111111011111;
            14'h3e2e 	:	o_val <= 16'b0111111111011111;
            14'h3e2f 	:	o_val <= 16'b0111111111011111;
            14'h3e30 	:	o_val <= 16'b0111111111011111;
            14'h3e31 	:	o_val <= 16'b0111111111011111;
            14'h3e32 	:	o_val <= 16'b0111111111011111;
            14'h3e33 	:	o_val <= 16'b0111111111100000;
            14'h3e34 	:	o_val <= 16'b0111111111100000;
            14'h3e35 	:	o_val <= 16'b0111111111100000;
            14'h3e36 	:	o_val <= 16'b0111111111100000;
            14'h3e37 	:	o_val <= 16'b0111111111100000;
            14'h3e38 	:	o_val <= 16'b0111111111100000;
            14'h3e39 	:	o_val <= 16'b0111111111100000;
            14'h3e3a 	:	o_val <= 16'b0111111111100001;
            14'h3e3b 	:	o_val <= 16'b0111111111100001;
            14'h3e3c 	:	o_val <= 16'b0111111111100001;
            14'h3e3d 	:	o_val <= 16'b0111111111100001;
            14'h3e3e 	:	o_val <= 16'b0111111111100001;
            14'h3e3f 	:	o_val <= 16'b0111111111100001;
            14'h3e40 	:	o_val <= 16'b0111111111100001;
            14'h3e41 	:	o_val <= 16'b0111111111100001;
            14'h3e42 	:	o_val <= 16'b0111111111100010;
            14'h3e43 	:	o_val <= 16'b0111111111100010;
            14'h3e44 	:	o_val <= 16'b0111111111100010;
            14'h3e45 	:	o_val <= 16'b0111111111100010;
            14'h3e46 	:	o_val <= 16'b0111111111100010;
            14'h3e47 	:	o_val <= 16'b0111111111100010;
            14'h3e48 	:	o_val <= 16'b0111111111100010;
            14'h3e49 	:	o_val <= 16'b0111111111100011;
            14'h3e4a 	:	o_val <= 16'b0111111111100011;
            14'h3e4b 	:	o_val <= 16'b0111111111100011;
            14'h3e4c 	:	o_val <= 16'b0111111111100011;
            14'h3e4d 	:	o_val <= 16'b0111111111100011;
            14'h3e4e 	:	o_val <= 16'b0111111111100011;
            14'h3e4f 	:	o_val <= 16'b0111111111100011;
            14'h3e50 	:	o_val <= 16'b0111111111100011;
            14'h3e51 	:	o_val <= 16'b0111111111100100;
            14'h3e52 	:	o_val <= 16'b0111111111100100;
            14'h3e53 	:	o_val <= 16'b0111111111100100;
            14'h3e54 	:	o_val <= 16'b0111111111100100;
            14'h3e55 	:	o_val <= 16'b0111111111100100;
            14'h3e56 	:	o_val <= 16'b0111111111100100;
            14'h3e57 	:	o_val <= 16'b0111111111100100;
            14'h3e58 	:	o_val <= 16'b0111111111100100;
            14'h3e59 	:	o_val <= 16'b0111111111100101;
            14'h3e5a 	:	o_val <= 16'b0111111111100101;
            14'h3e5b 	:	o_val <= 16'b0111111111100101;
            14'h3e5c 	:	o_val <= 16'b0111111111100101;
            14'h3e5d 	:	o_val <= 16'b0111111111100101;
            14'h3e5e 	:	o_val <= 16'b0111111111100101;
            14'h3e5f 	:	o_val <= 16'b0111111111100101;
            14'h3e60 	:	o_val <= 16'b0111111111100110;
            14'h3e61 	:	o_val <= 16'b0111111111100110;
            14'h3e62 	:	o_val <= 16'b0111111111100110;
            14'h3e63 	:	o_val <= 16'b0111111111100110;
            14'h3e64 	:	o_val <= 16'b0111111111100110;
            14'h3e65 	:	o_val <= 16'b0111111111100110;
            14'h3e66 	:	o_val <= 16'b0111111111100110;
            14'h3e67 	:	o_val <= 16'b0111111111100110;
            14'h3e68 	:	o_val <= 16'b0111111111100110;
            14'h3e69 	:	o_val <= 16'b0111111111100111;
            14'h3e6a 	:	o_val <= 16'b0111111111100111;
            14'h3e6b 	:	o_val <= 16'b0111111111100111;
            14'h3e6c 	:	o_val <= 16'b0111111111100111;
            14'h3e6d 	:	o_val <= 16'b0111111111100111;
            14'h3e6e 	:	o_val <= 16'b0111111111100111;
            14'h3e6f 	:	o_val <= 16'b0111111111100111;
            14'h3e70 	:	o_val <= 16'b0111111111100111;
            14'h3e71 	:	o_val <= 16'b0111111111101000;
            14'h3e72 	:	o_val <= 16'b0111111111101000;
            14'h3e73 	:	o_val <= 16'b0111111111101000;
            14'h3e74 	:	o_val <= 16'b0111111111101000;
            14'h3e75 	:	o_val <= 16'b0111111111101000;
            14'h3e76 	:	o_val <= 16'b0111111111101000;
            14'h3e77 	:	o_val <= 16'b0111111111101000;
            14'h3e78 	:	o_val <= 16'b0111111111101000;
            14'h3e79 	:	o_val <= 16'b0111111111101001;
            14'h3e7a 	:	o_val <= 16'b0111111111101001;
            14'h3e7b 	:	o_val <= 16'b0111111111101001;
            14'h3e7c 	:	o_val <= 16'b0111111111101001;
            14'h3e7d 	:	o_val <= 16'b0111111111101001;
            14'h3e7e 	:	o_val <= 16'b0111111111101001;
            14'h3e7f 	:	o_val <= 16'b0111111111101001;
            14'h3e80 	:	o_val <= 16'b0111111111101001;
            14'h3e81 	:	o_val <= 16'b0111111111101001;
            14'h3e82 	:	o_val <= 16'b0111111111101010;
            14'h3e83 	:	o_val <= 16'b0111111111101010;
            14'h3e84 	:	o_val <= 16'b0111111111101010;
            14'h3e85 	:	o_val <= 16'b0111111111101010;
            14'h3e86 	:	o_val <= 16'b0111111111101010;
            14'h3e87 	:	o_val <= 16'b0111111111101010;
            14'h3e88 	:	o_val <= 16'b0111111111101010;
            14'h3e89 	:	o_val <= 16'b0111111111101010;
            14'h3e8a 	:	o_val <= 16'b0111111111101010;
            14'h3e8b 	:	o_val <= 16'b0111111111101011;
            14'h3e8c 	:	o_val <= 16'b0111111111101011;
            14'h3e8d 	:	o_val <= 16'b0111111111101011;
            14'h3e8e 	:	o_val <= 16'b0111111111101011;
            14'h3e8f 	:	o_val <= 16'b0111111111101011;
            14'h3e90 	:	o_val <= 16'b0111111111101011;
            14'h3e91 	:	o_val <= 16'b0111111111101011;
            14'h3e92 	:	o_val <= 16'b0111111111101011;
            14'h3e93 	:	o_val <= 16'b0111111111101011;
            14'h3e94 	:	o_val <= 16'b0111111111101100;
            14'h3e95 	:	o_val <= 16'b0111111111101100;
            14'h3e96 	:	o_val <= 16'b0111111111101100;
            14'h3e97 	:	o_val <= 16'b0111111111101100;
            14'h3e98 	:	o_val <= 16'b0111111111101100;
            14'h3e99 	:	o_val <= 16'b0111111111101100;
            14'h3e9a 	:	o_val <= 16'b0111111111101100;
            14'h3e9b 	:	o_val <= 16'b0111111111101100;
            14'h3e9c 	:	o_val <= 16'b0111111111101100;
            14'h3e9d 	:	o_val <= 16'b0111111111101101;
            14'h3e9e 	:	o_val <= 16'b0111111111101101;
            14'h3e9f 	:	o_val <= 16'b0111111111101101;
            14'h3ea0 	:	o_val <= 16'b0111111111101101;
            14'h3ea1 	:	o_val <= 16'b0111111111101101;
            14'h3ea2 	:	o_val <= 16'b0111111111101101;
            14'h3ea3 	:	o_val <= 16'b0111111111101101;
            14'h3ea4 	:	o_val <= 16'b0111111111101101;
            14'h3ea5 	:	o_val <= 16'b0111111111101101;
            14'h3ea6 	:	o_val <= 16'b0111111111101110;
            14'h3ea7 	:	o_val <= 16'b0111111111101110;
            14'h3ea8 	:	o_val <= 16'b0111111111101110;
            14'h3ea9 	:	o_val <= 16'b0111111111101110;
            14'h3eaa 	:	o_val <= 16'b0111111111101110;
            14'h3eab 	:	o_val <= 16'b0111111111101110;
            14'h3eac 	:	o_val <= 16'b0111111111101110;
            14'h3ead 	:	o_val <= 16'b0111111111101110;
            14'h3eae 	:	o_val <= 16'b0111111111101110;
            14'h3eaf 	:	o_val <= 16'b0111111111101110;
            14'h3eb0 	:	o_val <= 16'b0111111111101111;
            14'h3eb1 	:	o_val <= 16'b0111111111101111;
            14'h3eb2 	:	o_val <= 16'b0111111111101111;
            14'h3eb3 	:	o_val <= 16'b0111111111101111;
            14'h3eb4 	:	o_val <= 16'b0111111111101111;
            14'h3eb5 	:	o_val <= 16'b0111111111101111;
            14'h3eb6 	:	o_val <= 16'b0111111111101111;
            14'h3eb7 	:	o_val <= 16'b0111111111101111;
            14'h3eb8 	:	o_val <= 16'b0111111111101111;
            14'h3eb9 	:	o_val <= 16'b0111111111101111;
            14'h3eba 	:	o_val <= 16'b0111111111110000;
            14'h3ebb 	:	o_val <= 16'b0111111111110000;
            14'h3ebc 	:	o_val <= 16'b0111111111110000;
            14'h3ebd 	:	o_val <= 16'b0111111111110000;
            14'h3ebe 	:	o_val <= 16'b0111111111110000;
            14'h3ebf 	:	o_val <= 16'b0111111111110000;
            14'h3ec0 	:	o_val <= 16'b0111111111110000;
            14'h3ec1 	:	o_val <= 16'b0111111111110000;
            14'h3ec2 	:	o_val <= 16'b0111111111110000;
            14'h3ec3 	:	o_val <= 16'b0111111111110000;
            14'h3ec4 	:	o_val <= 16'b0111111111110001;
            14'h3ec5 	:	o_val <= 16'b0111111111110001;
            14'h3ec6 	:	o_val <= 16'b0111111111110001;
            14'h3ec7 	:	o_val <= 16'b0111111111110001;
            14'h3ec8 	:	o_val <= 16'b0111111111110001;
            14'h3ec9 	:	o_val <= 16'b0111111111110001;
            14'h3eca 	:	o_val <= 16'b0111111111110001;
            14'h3ecb 	:	o_val <= 16'b0111111111110001;
            14'h3ecc 	:	o_val <= 16'b0111111111110001;
            14'h3ecd 	:	o_val <= 16'b0111111111110001;
            14'h3ece 	:	o_val <= 16'b0111111111110001;
            14'h3ecf 	:	o_val <= 16'b0111111111110010;
            14'h3ed0 	:	o_val <= 16'b0111111111110010;
            14'h3ed1 	:	o_val <= 16'b0111111111110010;
            14'h3ed2 	:	o_val <= 16'b0111111111110010;
            14'h3ed3 	:	o_val <= 16'b0111111111110010;
            14'h3ed4 	:	o_val <= 16'b0111111111110010;
            14'h3ed5 	:	o_val <= 16'b0111111111110010;
            14'h3ed6 	:	o_val <= 16'b0111111111110010;
            14'h3ed7 	:	o_val <= 16'b0111111111110010;
            14'h3ed8 	:	o_val <= 16'b0111111111110010;
            14'h3ed9 	:	o_val <= 16'b0111111111110010;
            14'h3eda 	:	o_val <= 16'b0111111111110011;
            14'h3edb 	:	o_val <= 16'b0111111111110011;
            14'h3edc 	:	o_val <= 16'b0111111111110011;
            14'h3edd 	:	o_val <= 16'b0111111111110011;
            14'h3ede 	:	o_val <= 16'b0111111111110011;
            14'h3edf 	:	o_val <= 16'b0111111111110011;
            14'h3ee0 	:	o_val <= 16'b0111111111110011;
            14'h3ee1 	:	o_val <= 16'b0111111111110011;
            14'h3ee2 	:	o_val <= 16'b0111111111110011;
            14'h3ee3 	:	o_val <= 16'b0111111111110011;
            14'h3ee4 	:	o_val <= 16'b0111111111110011;
            14'h3ee5 	:	o_val <= 16'b0111111111110011;
            14'h3ee6 	:	o_val <= 16'b0111111111110100;
            14'h3ee7 	:	o_val <= 16'b0111111111110100;
            14'h3ee8 	:	o_val <= 16'b0111111111110100;
            14'h3ee9 	:	o_val <= 16'b0111111111110100;
            14'h3eea 	:	o_val <= 16'b0111111111110100;
            14'h3eeb 	:	o_val <= 16'b0111111111110100;
            14'h3eec 	:	o_val <= 16'b0111111111110100;
            14'h3eed 	:	o_val <= 16'b0111111111110100;
            14'h3eee 	:	o_val <= 16'b0111111111110100;
            14'h3eef 	:	o_val <= 16'b0111111111110100;
            14'h3ef0 	:	o_val <= 16'b0111111111110100;
            14'h3ef1 	:	o_val <= 16'b0111111111110100;
            14'h3ef2 	:	o_val <= 16'b0111111111110101;
            14'h3ef3 	:	o_val <= 16'b0111111111110101;
            14'h3ef4 	:	o_val <= 16'b0111111111110101;
            14'h3ef5 	:	o_val <= 16'b0111111111110101;
            14'h3ef6 	:	o_val <= 16'b0111111111110101;
            14'h3ef7 	:	o_val <= 16'b0111111111110101;
            14'h3ef8 	:	o_val <= 16'b0111111111110101;
            14'h3ef9 	:	o_val <= 16'b0111111111110101;
            14'h3efa 	:	o_val <= 16'b0111111111110101;
            14'h3efb 	:	o_val <= 16'b0111111111110101;
            14'h3efc 	:	o_val <= 16'b0111111111110101;
            14'h3efd 	:	o_val <= 16'b0111111111110101;
            14'h3efe 	:	o_val <= 16'b0111111111110110;
            14'h3eff 	:	o_val <= 16'b0111111111110110;
            14'h3f00 	:	o_val <= 16'b0111111111110110;
            14'h3f01 	:	o_val <= 16'b0111111111110110;
            14'h3f02 	:	o_val <= 16'b0111111111110110;
            14'h3f03 	:	o_val <= 16'b0111111111110110;
            14'h3f04 	:	o_val <= 16'b0111111111110110;
            14'h3f05 	:	o_val <= 16'b0111111111110110;
            14'h3f06 	:	o_val <= 16'b0111111111110110;
            14'h3f07 	:	o_val <= 16'b0111111111110110;
            14'h3f08 	:	o_val <= 16'b0111111111110110;
            14'h3f09 	:	o_val <= 16'b0111111111110110;
            14'h3f0a 	:	o_val <= 16'b0111111111110110;
            14'h3f0b 	:	o_val <= 16'b0111111111110110;
            14'h3f0c 	:	o_val <= 16'b0111111111110111;
            14'h3f0d 	:	o_val <= 16'b0111111111110111;
            14'h3f0e 	:	o_val <= 16'b0111111111110111;
            14'h3f0f 	:	o_val <= 16'b0111111111110111;
            14'h3f10 	:	o_val <= 16'b0111111111110111;
            14'h3f11 	:	o_val <= 16'b0111111111110111;
            14'h3f12 	:	o_val <= 16'b0111111111110111;
            14'h3f13 	:	o_val <= 16'b0111111111110111;
            14'h3f14 	:	o_val <= 16'b0111111111110111;
            14'h3f15 	:	o_val <= 16'b0111111111110111;
            14'h3f16 	:	o_val <= 16'b0111111111110111;
            14'h3f17 	:	o_val <= 16'b0111111111110111;
            14'h3f18 	:	o_val <= 16'b0111111111110111;
            14'h3f19 	:	o_val <= 16'b0111111111110111;
            14'h3f1a 	:	o_val <= 16'b0111111111111000;
            14'h3f1b 	:	o_val <= 16'b0111111111111000;
            14'h3f1c 	:	o_val <= 16'b0111111111111000;
            14'h3f1d 	:	o_val <= 16'b0111111111111000;
            14'h3f1e 	:	o_val <= 16'b0111111111111000;
            14'h3f1f 	:	o_val <= 16'b0111111111111000;
            14'h3f20 	:	o_val <= 16'b0111111111111000;
            14'h3f21 	:	o_val <= 16'b0111111111111000;
            14'h3f22 	:	o_val <= 16'b0111111111111000;
            14'h3f23 	:	o_val <= 16'b0111111111111000;
            14'h3f24 	:	o_val <= 16'b0111111111111000;
            14'h3f25 	:	o_val <= 16'b0111111111111000;
            14'h3f26 	:	o_val <= 16'b0111111111111000;
            14'h3f27 	:	o_val <= 16'b0111111111111000;
            14'h3f28 	:	o_val <= 16'b0111111111111001;
            14'h3f29 	:	o_val <= 16'b0111111111111001;
            14'h3f2a 	:	o_val <= 16'b0111111111111001;
            14'h3f2b 	:	o_val <= 16'b0111111111111001;
            14'h3f2c 	:	o_val <= 16'b0111111111111001;
            14'h3f2d 	:	o_val <= 16'b0111111111111001;
            14'h3f2e 	:	o_val <= 16'b0111111111111001;
            14'h3f2f 	:	o_val <= 16'b0111111111111001;
            14'h3f30 	:	o_val <= 16'b0111111111111001;
            14'h3f31 	:	o_val <= 16'b0111111111111001;
            14'h3f32 	:	o_val <= 16'b0111111111111001;
            14'h3f33 	:	o_val <= 16'b0111111111111001;
            14'h3f34 	:	o_val <= 16'b0111111111111001;
            14'h3f35 	:	o_val <= 16'b0111111111111001;
            14'h3f36 	:	o_val <= 16'b0111111111111001;
            14'h3f37 	:	o_val <= 16'b0111111111111001;
            14'h3f38 	:	o_val <= 16'b0111111111111010;
            14'h3f39 	:	o_val <= 16'b0111111111111010;
            14'h3f3a 	:	o_val <= 16'b0111111111111010;
            14'h3f3b 	:	o_val <= 16'b0111111111111010;
            14'h3f3c 	:	o_val <= 16'b0111111111111010;
            14'h3f3d 	:	o_val <= 16'b0111111111111010;
            14'h3f3e 	:	o_val <= 16'b0111111111111010;
            14'h3f3f 	:	o_val <= 16'b0111111111111010;
            14'h3f40 	:	o_val <= 16'b0111111111111010;
            14'h3f41 	:	o_val <= 16'b0111111111111010;
            14'h3f42 	:	o_val <= 16'b0111111111111010;
            14'h3f43 	:	o_val <= 16'b0111111111111010;
            14'h3f44 	:	o_val <= 16'b0111111111111010;
            14'h3f45 	:	o_val <= 16'b0111111111111010;
            14'h3f46 	:	o_val <= 16'b0111111111111010;
            14'h3f47 	:	o_val <= 16'b0111111111111010;
            14'h3f48 	:	o_val <= 16'b0111111111111010;
            14'h3f49 	:	o_val <= 16'b0111111111111010;
            14'h3f4a 	:	o_val <= 16'b0111111111111011;
            14'h3f4b 	:	o_val <= 16'b0111111111111011;
            14'h3f4c 	:	o_val <= 16'b0111111111111011;
            14'h3f4d 	:	o_val <= 16'b0111111111111011;
            14'h3f4e 	:	o_val <= 16'b0111111111111011;
            14'h3f4f 	:	o_val <= 16'b0111111111111011;
            14'h3f50 	:	o_val <= 16'b0111111111111011;
            14'h3f51 	:	o_val <= 16'b0111111111111011;
            14'h3f52 	:	o_val <= 16'b0111111111111011;
            14'h3f53 	:	o_val <= 16'b0111111111111011;
            14'h3f54 	:	o_val <= 16'b0111111111111011;
            14'h3f55 	:	o_val <= 16'b0111111111111011;
            14'h3f56 	:	o_val <= 16'b0111111111111011;
            14'h3f57 	:	o_val <= 16'b0111111111111011;
            14'h3f58 	:	o_val <= 16'b0111111111111011;
            14'h3f59 	:	o_val <= 16'b0111111111111011;
            14'h3f5a 	:	o_val <= 16'b0111111111111011;
            14'h3f5b 	:	o_val <= 16'b0111111111111011;
            14'h3f5c 	:	o_val <= 16'b0111111111111011;
            14'h3f5d 	:	o_val <= 16'b0111111111111100;
            14'h3f5e 	:	o_val <= 16'b0111111111111100;
            14'h3f5f 	:	o_val <= 16'b0111111111111100;
            14'h3f60 	:	o_val <= 16'b0111111111111100;
            14'h3f61 	:	o_val <= 16'b0111111111111100;
            14'h3f62 	:	o_val <= 16'b0111111111111100;
            14'h3f63 	:	o_val <= 16'b0111111111111100;
            14'h3f64 	:	o_val <= 16'b0111111111111100;
            14'h3f65 	:	o_val <= 16'b0111111111111100;
            14'h3f66 	:	o_val <= 16'b0111111111111100;
            14'h3f67 	:	o_val <= 16'b0111111111111100;
            14'h3f68 	:	o_val <= 16'b0111111111111100;
            14'h3f69 	:	o_val <= 16'b0111111111111100;
            14'h3f6a 	:	o_val <= 16'b0111111111111100;
            14'h3f6b 	:	o_val <= 16'b0111111111111100;
            14'h3f6c 	:	o_val <= 16'b0111111111111100;
            14'h3f6d 	:	o_val <= 16'b0111111111111100;
            14'h3f6e 	:	o_val <= 16'b0111111111111100;
            14'h3f6f 	:	o_val <= 16'b0111111111111100;
            14'h3f70 	:	o_val <= 16'b0111111111111100;
            14'h3f71 	:	o_val <= 16'b0111111111111100;
            14'h3f72 	:	o_val <= 16'b0111111111111100;
            14'h3f73 	:	o_val <= 16'b0111111111111101;
            14'h3f74 	:	o_val <= 16'b0111111111111101;
            14'h3f75 	:	o_val <= 16'b0111111111111101;
            14'h3f76 	:	o_val <= 16'b0111111111111101;
            14'h3f77 	:	o_val <= 16'b0111111111111101;
            14'h3f78 	:	o_val <= 16'b0111111111111101;
            14'h3f79 	:	o_val <= 16'b0111111111111101;
            14'h3f7a 	:	o_val <= 16'b0111111111111101;
            14'h3f7b 	:	o_val <= 16'b0111111111111101;
            14'h3f7c 	:	o_val <= 16'b0111111111111101;
            14'h3f7d 	:	o_val <= 16'b0111111111111101;
            14'h3f7e 	:	o_val <= 16'b0111111111111101;
            14'h3f7f 	:	o_val <= 16'b0111111111111101;
            14'h3f80 	:	o_val <= 16'b0111111111111101;
            14'h3f81 	:	o_val <= 16'b0111111111111101;
            14'h3f82 	:	o_val <= 16'b0111111111111101;
            14'h3f83 	:	o_val <= 16'b0111111111111101;
            14'h3f84 	:	o_val <= 16'b0111111111111101;
            14'h3f85 	:	o_val <= 16'b0111111111111101;
            14'h3f86 	:	o_val <= 16'b0111111111111101;
            14'h3f87 	:	o_val <= 16'b0111111111111101;
            14'h3f88 	:	o_val <= 16'b0111111111111101;
            14'h3f89 	:	o_val <= 16'b0111111111111101;
            14'h3f8a 	:	o_val <= 16'b0111111111111101;
            14'h3f8b 	:	o_val <= 16'b0111111111111101;
            14'h3f8c 	:	o_val <= 16'b0111111111111101;
            14'h3f8d 	:	o_val <= 16'b0111111111111110;
            14'h3f8e 	:	o_val <= 16'b0111111111111110;
            14'h3f8f 	:	o_val <= 16'b0111111111111110;
            14'h3f90 	:	o_val <= 16'b0111111111111110;
            14'h3f91 	:	o_val <= 16'b0111111111111110;
            14'h3f92 	:	o_val <= 16'b0111111111111110;
            14'h3f93 	:	o_val <= 16'b0111111111111110;
            14'h3f94 	:	o_val <= 16'b0111111111111110;
            14'h3f95 	:	o_val <= 16'b0111111111111110;
            14'h3f96 	:	o_val <= 16'b0111111111111110;
            14'h3f97 	:	o_val <= 16'b0111111111111110;
            14'h3f98 	:	o_val <= 16'b0111111111111110;
            14'h3f99 	:	o_val <= 16'b0111111111111110;
            14'h3f9a 	:	o_val <= 16'b0111111111111110;
            14'h3f9b 	:	o_val <= 16'b0111111111111110;
            14'h3f9c 	:	o_val <= 16'b0111111111111110;
            14'h3f9d 	:	o_val <= 16'b0111111111111110;
            14'h3f9e 	:	o_val <= 16'b0111111111111110;
            14'h3f9f 	:	o_val <= 16'b0111111111111110;
            14'h3fa0 	:	o_val <= 16'b0111111111111110;
            14'h3fa1 	:	o_val <= 16'b0111111111111110;
            14'h3fa2 	:	o_val <= 16'b0111111111111110;
            14'h3fa3 	:	o_val <= 16'b0111111111111110;
            14'h3fa4 	:	o_val <= 16'b0111111111111110;
            14'h3fa5 	:	o_val <= 16'b0111111111111110;
            14'h3fa6 	:	o_val <= 16'b0111111111111110;
            14'h3fa7 	:	o_val <= 16'b0111111111111110;
            14'h3fa8 	:	o_val <= 16'b0111111111111110;
            14'h3fa9 	:	o_val <= 16'b0111111111111110;
            14'h3faa 	:	o_val <= 16'b0111111111111110;
            14'h3fab 	:	o_val <= 16'b0111111111111110;
            14'h3fac 	:	o_val <= 16'b0111111111111110;
            14'h3fad 	:	o_val <= 16'b0111111111111110;
            14'h3fae 	:	o_val <= 16'b0111111111111110;
            14'h3faf 	:	o_val <= 16'b0111111111111111;
            14'h3fb0 	:	o_val <= 16'b0111111111111111;
            14'h3fb1 	:	o_val <= 16'b0111111111111111;
            14'h3fb2 	:	o_val <= 16'b0111111111111111;
            14'h3fb3 	:	o_val <= 16'b0111111111111111;
            14'h3fb4 	:	o_val <= 16'b0111111111111111;
            14'h3fb5 	:	o_val <= 16'b0111111111111111;
            14'h3fb6 	:	o_val <= 16'b0111111111111111;
            14'h3fb7 	:	o_val <= 16'b0111111111111111;
            14'h3fb8 	:	o_val <= 16'b0111111111111111;
            14'h3fb9 	:	o_val <= 16'b0111111111111111;
            14'h3fba 	:	o_val <= 16'b0111111111111111;
            14'h3fbb 	:	o_val <= 16'b0111111111111111;
            14'h3fbc 	:	o_val <= 16'b0111111111111111;
            14'h3fbd 	:	o_val <= 16'b0111111111111111;
            14'h3fbe 	:	o_val <= 16'b0111111111111111;
            14'h3fbf 	:	o_val <= 16'b0111111111111111;
            14'h3fc0 	:	o_val <= 16'b0111111111111111;
            14'h3fc1 	:	o_val <= 16'b0111111111111111;
            14'h3fc2 	:	o_val <= 16'b0111111111111111;
            14'h3fc3 	:	o_val <= 16'b0111111111111111;
            14'h3fc4 	:	o_val <= 16'b0111111111111111;
            14'h3fc5 	:	o_val <= 16'b0111111111111111;
            14'h3fc6 	:	o_val <= 16'b0111111111111111;
            14'h3fc7 	:	o_val <= 16'b0111111111111111;
            14'h3fc8 	:	o_val <= 16'b0111111111111111;
            14'h3fc9 	:	o_val <= 16'b0111111111111111;
            14'h3fca 	:	o_val <= 16'b0111111111111111;
            14'h3fcb 	:	o_val <= 16'b0111111111111111;
            14'h3fcc 	:	o_val <= 16'b0111111111111111;
            14'h3fcd 	:	o_val <= 16'b0111111111111111;
            14'h3fce 	:	o_val <= 16'b0111111111111111;
            14'h3fcf 	:	o_val <= 16'b0111111111111111;
            14'h3fd0 	:	o_val <= 16'b0111111111111111;
            14'h3fd1 	:	o_val <= 16'b0111111111111111;
            14'h3fd2 	:	o_val <= 16'b0111111111111111;
            14'h3fd3 	:	o_val <= 16'b0111111111111111;
            14'h3fd4 	:	o_val <= 16'b0111111111111111;
            14'h3fd5 	:	o_val <= 16'b0111111111111111;
            14'h3fd6 	:	o_val <= 16'b0111111111111111;
            14'h3fd7 	:	o_val <= 16'b0111111111111111;
            14'h3fd8 	:	o_val <= 16'b0111111111111111;
            14'h3fd9 	:	o_val <= 16'b0111111111111111;
            14'h3fda 	:	o_val <= 16'b0111111111111111;
            14'h3fdb 	:	o_val <= 16'b0111111111111111;
            14'h3fdc 	:	o_val <= 16'b0111111111111111;
            14'h3fdd 	:	o_val <= 16'b0111111111111111;
            14'h3fde 	:	o_val <= 16'b0111111111111111;
            14'h3fdf 	:	o_val <= 16'b0111111111111111;
            14'h3fe0 	:	o_val <= 16'b0111111111111111;
            14'h3fe1 	:	o_val <= 16'b0111111111111111;
            14'h3fe2 	:	o_val <= 16'b0111111111111111;
            14'h3fe3 	:	o_val <= 16'b0111111111111111;
            14'h3fe4 	:	o_val <= 16'b0111111111111111;
            14'h3fe5 	:	o_val <= 16'b0111111111111111;
            14'h3fe6 	:	o_val <= 16'b0111111111111111;
            14'h3fe7 	:	o_val <= 16'b0111111111111111;
            14'h3fe8 	:	o_val <= 16'b0111111111111111;
            14'h3fe9 	:	o_val <= 16'b0111111111111111;
            14'h3fea 	:	o_val <= 16'b0111111111111111;
            14'h3feb 	:	o_val <= 16'b0111111111111111;
            14'h3fec 	:	o_val <= 16'b0111111111111111;
            14'h3fed 	:	o_val <= 16'b0111111111111111;
            14'h3fee 	:	o_val <= 16'b0111111111111111;
            14'h3fef 	:	o_val <= 16'b0111111111111111;
            14'h3ff0 	:	o_val <= 16'b0111111111111111;
            14'h3ff1 	:	o_val <= 16'b0111111111111111;
            14'h3ff2 	:	o_val <= 16'b0111111111111111;
            14'h3ff3 	:	o_val <= 16'b0111111111111111;
            14'h3ff4 	:	o_val <= 16'b0111111111111111;
            14'h3ff5 	:	o_val <= 16'b0111111111111111;
            14'h3ff6 	:	o_val <= 16'b0111111111111111;
            14'h3ff7 	:	o_val <= 16'b0111111111111111;
            14'h3ff8 	:	o_val <= 16'b0111111111111111;
            14'h3ff9 	:	o_val <= 16'b0111111111111111;
            14'h3ffa 	:	o_val <= 16'b0111111111111111;
            14'h3ffb 	:	o_val <= 16'b0111111111111111;
            14'h3ffc 	:	o_val <= 16'b0111111111111111;
            14'h3ffd 	:	o_val <= 16'b0111111111111111;
            14'h3ffe 	:	o_val <= 16'b0111111111111111;
            14'h3fff 	:	o_val <= 16'b0111111111111111;
				 default		:	o_val <= 16'b0;
			endcase
		end
endmodule
                                        
