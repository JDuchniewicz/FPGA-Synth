

module quarter_sine_lut(input[13:0] phase,
								output reg[15:0] val_out); //is reg needed here? try removing
		always @(phase) begin
			case(phase)
             14'h000 	:	val_out <= 16'h0003;
             14'h001 	:	val_out <= 16'h0009;
             14'h002 	:	val_out <= 16'h000f;
             14'h003 	:	val_out <= 16'h0015;
             14'h004 	:	val_out <= 16'h001c;
             14'h005 	:	val_out <= 16'h0022;
             14'h006 	:	val_out <= 16'h0028;
             14'h007 	:	val_out <= 16'h002f;
             14'h008 	:	val_out <= 16'h0035;
             14'h009 	:	val_out <= 16'h003b;
             14'h00a 	:	val_out <= 16'h0041;
             14'h00b 	:	val_out <= 16'h0048;
             14'h00c 	:	val_out <= 16'h004e;
             14'h00d 	:	val_out <= 16'h0054;
             14'h00e 	:	val_out <= 16'h005b;
             14'h00f 	:	val_out <= 16'h0061;
             14'h010 	:	val_out <= 16'h0067;
             14'h011 	:	val_out <= 16'h006d;
             14'h012 	:	val_out <= 16'h0074;
             14'h013 	:	val_out <= 16'h007a;
             14'h014 	:	val_out <= 16'h0080;
             14'h015 	:	val_out <= 16'h0087;
             14'h016 	:	val_out <= 16'h008d;
             14'h017 	:	val_out <= 16'h0093;
             14'h018 	:	val_out <= 16'h0099;
             14'h019 	:	val_out <= 16'h00a0;
             14'h01a 	:	val_out <= 16'h00a6;
             14'h01b 	:	val_out <= 16'h00ac;
             14'h01c 	:	val_out <= 16'h00b3;
             14'h01d 	:	val_out <= 16'h00b9;
             14'h01e 	:	val_out <= 16'h00bf;
             14'h01f 	:	val_out <= 16'h00c5;
             14'h020 	:	val_out <= 16'h00cc;
             14'h021 	:	val_out <= 16'h00d2;
             14'h022 	:	val_out <= 16'h00d8;
             14'h023 	:	val_out <= 16'h00df;
             14'h024 	:	val_out <= 16'h00e5;
             14'h025 	:	val_out <= 16'h00eb;
             14'h026 	:	val_out <= 16'h00f1;
             14'h027 	:	val_out <= 16'h00f8;
             14'h028 	:	val_out <= 16'h00fe;
             14'h029 	:	val_out <= 16'h0104;
             14'h02a 	:	val_out <= 16'h010b;
             14'h02b 	:	val_out <= 16'h0111;
             14'h02c 	:	val_out <= 16'h0117;
             14'h02d 	:	val_out <= 16'h011d;
             14'h02e 	:	val_out <= 16'h0124;
             14'h02f 	:	val_out <= 16'h012a;
             14'h030 	:	val_out <= 16'h0130;
             14'h031 	:	val_out <= 16'h0137;
             14'h032 	:	val_out <= 16'h013d;
             14'h033 	:	val_out <= 16'h0143;
             14'h034 	:	val_out <= 16'h0149;
             14'h035 	:	val_out <= 16'h0150;
             14'h036 	:	val_out <= 16'h0156;
             14'h037 	:	val_out <= 16'h015c;
             14'h038 	:	val_out <= 16'h0162;
             14'h039 	:	val_out <= 16'h0169;
             14'h03a 	:	val_out <= 16'h016f;
             14'h03b 	:	val_out <= 16'h0175;
             14'h03c 	:	val_out <= 16'h017c;
             14'h03d 	:	val_out <= 16'h0182;
             14'h03e 	:	val_out <= 16'h0188;
             14'h03f 	:	val_out <= 16'h018e;
             14'h040 	:	val_out <= 16'h0195;
             14'h041 	:	val_out <= 16'h019b;
             14'h042 	:	val_out <= 16'h01a1;
             14'h043 	:	val_out <= 16'h01a8;
             14'h044 	:	val_out <= 16'h01ae;
             14'h045 	:	val_out <= 16'h01b4;
             14'h046 	:	val_out <= 16'h01ba;
             14'h047 	:	val_out <= 16'h01c1;
             14'h048 	:	val_out <= 16'h01c7;
             14'h049 	:	val_out <= 16'h01cd;
             14'h04a 	:	val_out <= 16'h01d4;
             14'h04b 	:	val_out <= 16'h01da;
             14'h04c 	:	val_out <= 16'h01e0;
             14'h04d 	:	val_out <= 16'h01e6;
             14'h04e 	:	val_out <= 16'h01ed;
             14'h04f 	:	val_out <= 16'h01f3;
             14'h050 	:	val_out <= 16'h01f9;
             14'h051 	:	val_out <= 16'h0200;
             14'h052 	:	val_out <= 16'h0206;
             14'h053 	:	val_out <= 16'h020c;
             14'h054 	:	val_out <= 16'h0212;
             14'h055 	:	val_out <= 16'h0219;
             14'h056 	:	val_out <= 16'h021f;
             14'h057 	:	val_out <= 16'h0225;
             14'h058 	:	val_out <= 16'h022c;
             14'h059 	:	val_out <= 16'h0232;
             14'h05a 	:	val_out <= 16'h0238;
             14'h05b 	:	val_out <= 16'h023e;
             14'h05c 	:	val_out <= 16'h0245;
             14'h05d 	:	val_out <= 16'h024b;
             14'h05e 	:	val_out <= 16'h0251;
             14'h05f 	:	val_out <= 16'h0258;
             14'h060 	:	val_out <= 16'h025e;
             14'h061 	:	val_out <= 16'h0264;
             14'h062 	:	val_out <= 16'h026a;
             14'h063 	:	val_out <= 16'h0271;
             14'h064 	:	val_out <= 16'h0277;
             14'h065 	:	val_out <= 16'h027d;
             14'h066 	:	val_out <= 16'h0284;
             14'h067 	:	val_out <= 16'h028a;
             14'h068 	:	val_out <= 16'h0290;
             14'h069 	:	val_out <= 16'h0296;
             14'h06a 	:	val_out <= 16'h029d;
             14'h06b 	:	val_out <= 16'h02a3;
             14'h06c 	:	val_out <= 16'h02a9;
             14'h06d 	:	val_out <= 16'h02af;
             14'h06e 	:	val_out <= 16'h02b6;
             14'h06f 	:	val_out <= 16'h02bc;
             14'h070 	:	val_out <= 16'h02c2;
             14'h071 	:	val_out <= 16'h02c9;
             14'h072 	:	val_out <= 16'h02cf;
             14'h073 	:	val_out <= 16'h02d5;
             14'h074 	:	val_out <= 16'h02db;
             14'h075 	:	val_out <= 16'h02e2;
             14'h076 	:	val_out <= 16'h02e8;
             14'h077 	:	val_out <= 16'h02ee;
             14'h078 	:	val_out <= 16'h02f5;
             14'h079 	:	val_out <= 16'h02fb;
             14'h07a 	:	val_out <= 16'h0301;
             14'h07b 	:	val_out <= 16'h0307;
             14'h07c 	:	val_out <= 16'h030e;
             14'h07d 	:	val_out <= 16'h0314;
             14'h07e 	:	val_out <= 16'h031a;
             14'h07f 	:	val_out <= 16'h0321;
             14'h080 	:	val_out <= 16'h0327;
             14'h081 	:	val_out <= 16'h032d;
             14'h082 	:	val_out <= 16'h0333;
             14'h083 	:	val_out <= 16'h033a;
             14'h084 	:	val_out <= 16'h0340;
             14'h085 	:	val_out <= 16'h0346;
             14'h086 	:	val_out <= 16'h034d;
             14'h087 	:	val_out <= 16'h0353;
             14'h088 	:	val_out <= 16'h0359;
             14'h089 	:	val_out <= 16'h035f;
             14'h08a 	:	val_out <= 16'h0366;
             14'h08b 	:	val_out <= 16'h036c;
             14'h08c 	:	val_out <= 16'h0372;
             14'h08d 	:	val_out <= 16'h0379;
             14'h08e 	:	val_out <= 16'h037f;
             14'h08f 	:	val_out <= 16'h0385;
             14'h090 	:	val_out <= 16'h038b;
             14'h091 	:	val_out <= 16'h0392;
             14'h092 	:	val_out <= 16'h0398;
             14'h093 	:	val_out <= 16'h039e;
             14'h094 	:	val_out <= 16'h03a5;
             14'h095 	:	val_out <= 16'h03ab;
             14'h096 	:	val_out <= 16'h03b1;
             14'h097 	:	val_out <= 16'h03b7;
             14'h098 	:	val_out <= 16'h03be;
             14'h099 	:	val_out <= 16'h03c4;
             14'h09a 	:	val_out <= 16'h03ca;
             14'h09b 	:	val_out <= 16'h03d0;
             14'h09c 	:	val_out <= 16'h03d7;
             14'h09d 	:	val_out <= 16'h03dd;
             14'h09e 	:	val_out <= 16'h03e3;
             14'h09f 	:	val_out <= 16'h03ea;
             14'h0a0 	:	val_out <= 16'h03f0;
             14'h0a1 	:	val_out <= 16'h03f6;
             14'h0a2 	:	val_out <= 16'h03fc;
             14'h0a3 	:	val_out <= 16'h0403;
             14'h0a4 	:	val_out <= 16'h0409;
             14'h0a5 	:	val_out <= 16'h040f;
             14'h0a6 	:	val_out <= 16'h0416;
             14'h0a7 	:	val_out <= 16'h041c;
             14'h0a8 	:	val_out <= 16'h0422;
             14'h0a9 	:	val_out <= 16'h0428;
             14'h0aa 	:	val_out <= 16'h042f;
             14'h0ab 	:	val_out <= 16'h0435;
             14'h0ac 	:	val_out <= 16'h043b;
             14'h0ad 	:	val_out <= 16'h0442;
             14'h0ae 	:	val_out <= 16'h0448;
             14'h0af 	:	val_out <= 16'h044e;
             14'h0b0 	:	val_out <= 16'h0454;
             14'h0b1 	:	val_out <= 16'h045b;
             14'h0b2 	:	val_out <= 16'h0461;
             14'h0b3 	:	val_out <= 16'h0467;
             14'h0b4 	:	val_out <= 16'h046e;
             14'h0b5 	:	val_out <= 16'h0474;
             14'h0b6 	:	val_out <= 16'h047a;
             14'h0b7 	:	val_out <= 16'h0480;
             14'h0b8 	:	val_out <= 16'h0487;
             14'h0b9 	:	val_out <= 16'h048d;
             14'h0ba 	:	val_out <= 16'h0493;
             14'h0bb 	:	val_out <= 16'h049a;
             14'h0bc 	:	val_out <= 16'h04a0;
             14'h0bd 	:	val_out <= 16'h04a6;
             14'h0be 	:	val_out <= 16'h04ac;
             14'h0bf 	:	val_out <= 16'h04b3;
             14'h0c0 	:	val_out <= 16'h04b9;
             14'h0c1 	:	val_out <= 16'h04bf;
             14'h0c2 	:	val_out <= 16'h04c6;
             14'h0c3 	:	val_out <= 16'h04cc;
             14'h0c4 	:	val_out <= 16'h04d2;
             14'h0c5 	:	val_out <= 16'h04d8;
             14'h0c6 	:	val_out <= 16'h04df;
             14'h0c7 	:	val_out <= 16'h04e5;
             14'h0c8 	:	val_out <= 16'h04eb;
             14'h0c9 	:	val_out <= 16'h04f1;
             14'h0ca 	:	val_out <= 16'h04f8;
             14'h0cb 	:	val_out <= 16'h04fe;
             14'h0cc 	:	val_out <= 16'h0504;
             14'h0cd 	:	val_out <= 16'h050b;
             14'h0ce 	:	val_out <= 16'h0511;
             14'h0cf 	:	val_out <= 16'h0517;
             14'h0d0 	:	val_out <= 16'h051d;
             14'h0d1 	:	val_out <= 16'h0524;
             14'h0d2 	:	val_out <= 16'h052a;
             14'h0d3 	:	val_out <= 16'h0530;
             14'h0d4 	:	val_out <= 16'h0537;
             14'h0d5 	:	val_out <= 16'h053d;
             14'h0d6 	:	val_out <= 16'h0543;
             14'h0d7 	:	val_out <= 16'h0549;
             14'h0d8 	:	val_out <= 16'h0550;
             14'h0d9 	:	val_out <= 16'h0556;
             14'h0da 	:	val_out <= 16'h055c;
             14'h0db 	:	val_out <= 16'h0563;
             14'h0dc 	:	val_out <= 16'h0569;
             14'h0dd 	:	val_out <= 16'h056f;
             14'h0de 	:	val_out <= 16'h0575;
             14'h0df 	:	val_out <= 16'h057c;
             14'h0e0 	:	val_out <= 16'h0582;
             14'h0e1 	:	val_out <= 16'h0588;
             14'h0e2 	:	val_out <= 16'h058f;
             14'h0e3 	:	val_out <= 16'h0595;
             14'h0e4 	:	val_out <= 16'h059b;
             14'h0e5 	:	val_out <= 16'h05a1;
             14'h0e6 	:	val_out <= 16'h05a8;
             14'h0e7 	:	val_out <= 16'h05ae;
             14'h0e8 	:	val_out <= 16'h05b4;
             14'h0e9 	:	val_out <= 16'h05bb;
             14'h0ea 	:	val_out <= 16'h05c1;
             14'h0eb 	:	val_out <= 16'h05c7;
             14'h0ec 	:	val_out <= 16'h05cd;
             14'h0ed 	:	val_out <= 16'h05d4;
             14'h0ee 	:	val_out <= 16'h05da;
             14'h0ef 	:	val_out <= 16'h05e0;
             14'h0f0 	:	val_out <= 16'h05e6;
             14'h0f1 	:	val_out <= 16'h05ed;
             14'h0f2 	:	val_out <= 16'h05f3;
             14'h0f3 	:	val_out <= 16'h05f9;
             14'h0f4 	:	val_out <= 16'h0600;
             14'h0f5 	:	val_out <= 16'h0606;
             14'h0f6 	:	val_out <= 16'h060c;
             14'h0f7 	:	val_out <= 16'h0612;
             14'h0f8 	:	val_out <= 16'h0619;
             14'h0f9 	:	val_out <= 16'h061f;
             14'h0fa 	:	val_out <= 16'h0625;
             14'h0fb 	:	val_out <= 16'h062c;
             14'h0fc 	:	val_out <= 16'h0632;
             14'h0fd 	:	val_out <= 16'h0638;
             14'h0fe 	:	val_out <= 16'h063e;
             14'h0ff 	:	val_out <= 16'h0645;
             14'h100 	:	val_out <= 16'h064b;
             14'h101 	:	val_out <= 16'h0651;
             14'h102 	:	val_out <= 16'h0658;
             14'h103 	:	val_out <= 16'h065e;
             14'h104 	:	val_out <= 16'h0664;
             14'h105 	:	val_out <= 16'h066a;
             14'h106 	:	val_out <= 16'h0671;
             14'h107 	:	val_out <= 16'h0677;
             14'h108 	:	val_out <= 16'h067d;
             14'h109 	:	val_out <= 16'h0684;
             14'h10a 	:	val_out <= 16'h068a;
             14'h10b 	:	val_out <= 16'h0690;
             14'h10c 	:	val_out <= 16'h0696;
             14'h10d 	:	val_out <= 16'h069d;
             14'h10e 	:	val_out <= 16'h06a3;
             14'h10f 	:	val_out <= 16'h06a9;
             14'h110 	:	val_out <= 16'h06af;
             14'h111 	:	val_out <= 16'h06b6;
             14'h112 	:	val_out <= 16'h06bc;
             14'h113 	:	val_out <= 16'h06c2;
             14'h114 	:	val_out <= 16'h06c9;
             14'h115 	:	val_out <= 16'h06cf;
             14'h116 	:	val_out <= 16'h06d5;
             14'h117 	:	val_out <= 16'h06db;
             14'h118 	:	val_out <= 16'h06e2;
             14'h119 	:	val_out <= 16'h06e8;
             14'h11a 	:	val_out <= 16'h06ee;
             14'h11b 	:	val_out <= 16'h06f5;
             14'h11c 	:	val_out <= 16'h06fb;
             14'h11d 	:	val_out <= 16'h0701;
             14'h11e 	:	val_out <= 16'h0707;
             14'h11f 	:	val_out <= 16'h070e;
             14'h120 	:	val_out <= 16'h0714;
             14'h121 	:	val_out <= 16'h071a;
             14'h122 	:	val_out <= 16'h0721;
             14'h123 	:	val_out <= 16'h0727;
             14'h124 	:	val_out <= 16'h072d;
             14'h125 	:	val_out <= 16'h0733;
             14'h126 	:	val_out <= 16'h073a;
             14'h127 	:	val_out <= 16'h0740;
             14'h128 	:	val_out <= 16'h0746;
             14'h129 	:	val_out <= 16'h074c;
             14'h12a 	:	val_out <= 16'h0753;
             14'h12b 	:	val_out <= 16'h0759;
             14'h12c 	:	val_out <= 16'h075f;
             14'h12d 	:	val_out <= 16'h0766;
             14'h12e 	:	val_out <= 16'h076c;
             14'h12f 	:	val_out <= 16'h0772;
             14'h130 	:	val_out <= 16'h0778;
             14'h131 	:	val_out <= 16'h077f;
             14'h132 	:	val_out <= 16'h0785;
             14'h133 	:	val_out <= 16'h078b;
             14'h134 	:	val_out <= 16'h0792;
             14'h135 	:	val_out <= 16'h0798;
             14'h136 	:	val_out <= 16'h079e;
             14'h137 	:	val_out <= 16'h07a4;
             14'h138 	:	val_out <= 16'h07ab;
             14'h139 	:	val_out <= 16'h07b1;
             14'h13a 	:	val_out <= 16'h07b7;
             14'h13b 	:	val_out <= 16'h07be;
             14'h13c 	:	val_out <= 16'h07c4;
             14'h13d 	:	val_out <= 16'h07ca;
             14'h13e 	:	val_out <= 16'h07d0;
             14'h13f 	:	val_out <= 16'h07d7;
             14'h140 	:	val_out <= 16'h07dd;
             14'h141 	:	val_out <= 16'h07e3;
             14'h142 	:	val_out <= 16'h07ea;
             14'h143 	:	val_out <= 16'h07f0;
             14'h144 	:	val_out <= 16'h07f6;
             14'h145 	:	val_out <= 16'h07fc;
             14'h146 	:	val_out <= 16'h0803;
             14'h147 	:	val_out <= 16'h0809;
             14'h148 	:	val_out <= 16'h080f;
             14'h149 	:	val_out <= 16'h0815;
             14'h14a 	:	val_out <= 16'h081c;
             14'h14b 	:	val_out <= 16'h0822;
             14'h14c 	:	val_out <= 16'h0828;
             14'h14d 	:	val_out <= 16'h082f;
             14'h14e 	:	val_out <= 16'h0835;
             14'h14f 	:	val_out <= 16'h083b;
             14'h150 	:	val_out <= 16'h0841;
             14'h151 	:	val_out <= 16'h0848;
             14'h152 	:	val_out <= 16'h084e;
             14'h153 	:	val_out <= 16'h0854;
             14'h154 	:	val_out <= 16'h085b;
             14'h155 	:	val_out <= 16'h0861;
             14'h156 	:	val_out <= 16'h0867;
             14'h157 	:	val_out <= 16'h086d;
             14'h158 	:	val_out <= 16'h0874;
             14'h159 	:	val_out <= 16'h087a;
             14'h15a 	:	val_out <= 16'h0880;
             14'h15b 	:	val_out <= 16'h0887;
             14'h15c 	:	val_out <= 16'h088d;
             14'h15d 	:	val_out <= 16'h0893;
             14'h15e 	:	val_out <= 16'h0899;
             14'h15f 	:	val_out <= 16'h08a0;
             14'h160 	:	val_out <= 16'h08a6;
             14'h161 	:	val_out <= 16'h08ac;
             14'h162 	:	val_out <= 16'h08b2;
             14'h163 	:	val_out <= 16'h08b9;
             14'h164 	:	val_out <= 16'h08bf;
             14'h165 	:	val_out <= 16'h08c5;
             14'h166 	:	val_out <= 16'h08cc;
             14'h167 	:	val_out <= 16'h08d2;
             14'h168 	:	val_out <= 16'h08d8;
             14'h169 	:	val_out <= 16'h08de;
             14'h16a 	:	val_out <= 16'h08e5;
             14'h16b 	:	val_out <= 16'h08eb;
             14'h16c 	:	val_out <= 16'h08f1;
             14'h16d 	:	val_out <= 16'h08f8;
             14'h16e 	:	val_out <= 16'h08fe;
             14'h16f 	:	val_out <= 16'h0904;
             14'h170 	:	val_out <= 16'h090a;
             14'h171 	:	val_out <= 16'h0911;
             14'h172 	:	val_out <= 16'h0917;
             14'h173 	:	val_out <= 16'h091d;
             14'h174 	:	val_out <= 16'h0923;
             14'h175 	:	val_out <= 16'h092a;
             14'h176 	:	val_out <= 16'h0930;
             14'h177 	:	val_out <= 16'h0936;
             14'h178 	:	val_out <= 16'h093d;
             14'h179 	:	val_out <= 16'h0943;
             14'h17a 	:	val_out <= 16'h0949;
             14'h17b 	:	val_out <= 16'h094f;
             14'h17c 	:	val_out <= 16'h0956;
             14'h17d 	:	val_out <= 16'h095c;
             14'h17e 	:	val_out <= 16'h0962;
             14'h17f 	:	val_out <= 16'h0969;
             14'h180 	:	val_out <= 16'h096f;
             14'h181 	:	val_out <= 16'h0975;
             14'h182 	:	val_out <= 16'h097b;
             14'h183 	:	val_out <= 16'h0982;
             14'h184 	:	val_out <= 16'h0988;
             14'h185 	:	val_out <= 16'h098e;
             14'h186 	:	val_out <= 16'h0995;
             14'h187 	:	val_out <= 16'h099b;
             14'h188 	:	val_out <= 16'h09a1;
             14'h189 	:	val_out <= 16'h09a7;
             14'h18a 	:	val_out <= 16'h09ae;
             14'h18b 	:	val_out <= 16'h09b4;
             14'h18c 	:	val_out <= 16'h09ba;
             14'h18d 	:	val_out <= 16'h09c0;
             14'h18e 	:	val_out <= 16'h09c7;
             14'h18f 	:	val_out <= 16'h09cd;
             14'h190 	:	val_out <= 16'h09d3;
             14'h191 	:	val_out <= 16'h09da;
             14'h192 	:	val_out <= 16'h09e0;
             14'h193 	:	val_out <= 16'h09e6;
             14'h194 	:	val_out <= 16'h09ec;
             14'h195 	:	val_out <= 16'h09f3;
             14'h196 	:	val_out <= 16'h09f9;
             14'h197 	:	val_out <= 16'h09ff;
             14'h198 	:	val_out <= 16'h0a06;
             14'h199 	:	val_out <= 16'h0a0c;
             14'h19a 	:	val_out <= 16'h0a12;
             14'h19b 	:	val_out <= 16'h0a18;
             14'h19c 	:	val_out <= 16'h0a1f;
             14'h19d 	:	val_out <= 16'h0a25;
             14'h19e 	:	val_out <= 16'h0a2b;
             14'h19f 	:	val_out <= 16'h0a31;
             14'h1a0 	:	val_out <= 16'h0a38;
             14'h1a1 	:	val_out <= 16'h0a3e;
             14'h1a2 	:	val_out <= 16'h0a44;
             14'h1a3 	:	val_out <= 16'h0a4b;
             14'h1a4 	:	val_out <= 16'h0a51;
             14'h1a5 	:	val_out <= 16'h0a57;
             14'h1a6 	:	val_out <= 16'h0a5d;
             14'h1a7 	:	val_out <= 16'h0a64;
             14'h1a8 	:	val_out <= 16'h0a6a;
             14'h1a9 	:	val_out <= 16'h0a70;
             14'h1aa 	:	val_out <= 16'h0a77;
             14'h1ab 	:	val_out <= 16'h0a7d;
             14'h1ac 	:	val_out <= 16'h0a83;
             14'h1ad 	:	val_out <= 16'h0a89;
             14'h1ae 	:	val_out <= 16'h0a90;
             14'h1af 	:	val_out <= 16'h0a96;
             14'h1b0 	:	val_out <= 16'h0a9c;
             14'h1b1 	:	val_out <= 16'h0aa2;
             14'h1b2 	:	val_out <= 16'h0aa9;
             14'h1b3 	:	val_out <= 16'h0aaf;
             14'h1b4 	:	val_out <= 16'h0ab5;
             14'h1b5 	:	val_out <= 16'h0abc;
             14'h1b6 	:	val_out <= 16'h0ac2;
             14'h1b7 	:	val_out <= 16'h0ac8;
             14'h1b8 	:	val_out <= 16'h0ace;
             14'h1b9 	:	val_out <= 16'h0ad5;
             14'h1ba 	:	val_out <= 16'h0adb;
             14'h1bb 	:	val_out <= 16'h0ae1;
             14'h1bc 	:	val_out <= 16'h0ae8;
             14'h1bd 	:	val_out <= 16'h0aee;
             14'h1be 	:	val_out <= 16'h0af4;
             14'h1bf 	:	val_out <= 16'h0afa;
             14'h1c0 	:	val_out <= 16'h0b01;
             14'h1c1 	:	val_out <= 16'h0b07;
             14'h1c2 	:	val_out <= 16'h0b0d;
             14'h1c3 	:	val_out <= 16'h0b13;
             14'h1c4 	:	val_out <= 16'h0b1a;
             14'h1c5 	:	val_out <= 16'h0b20;
             14'h1c6 	:	val_out <= 16'h0b26;
             14'h1c7 	:	val_out <= 16'h0b2d;
             14'h1c8 	:	val_out <= 16'h0b33;
             14'h1c9 	:	val_out <= 16'h0b39;
             14'h1ca 	:	val_out <= 16'h0b3f;
             14'h1cb 	:	val_out <= 16'h0b46;
             14'h1cc 	:	val_out <= 16'h0b4c;
             14'h1cd 	:	val_out <= 16'h0b52;
             14'h1ce 	:	val_out <= 16'h0b59;
             14'h1cf 	:	val_out <= 16'h0b5f;
             14'h1d0 	:	val_out <= 16'h0b65;
             14'h1d1 	:	val_out <= 16'h0b6b;
             14'h1d2 	:	val_out <= 16'h0b72;
             14'h1d3 	:	val_out <= 16'h0b78;
             14'h1d4 	:	val_out <= 16'h0b7e;
             14'h1d5 	:	val_out <= 16'h0b84;
             14'h1d6 	:	val_out <= 16'h0b8b;
             14'h1d7 	:	val_out <= 16'h0b91;
             14'h1d8 	:	val_out <= 16'h0b97;
             14'h1d9 	:	val_out <= 16'h0b9e;
             14'h1da 	:	val_out <= 16'h0ba4;
             14'h1db 	:	val_out <= 16'h0baa;
             14'h1dc 	:	val_out <= 16'h0bb0;
             14'h1dd 	:	val_out <= 16'h0bb7;
             14'h1de 	:	val_out <= 16'h0bbd;
             14'h1df 	:	val_out <= 16'h0bc3;
             14'h1e0 	:	val_out <= 16'h0bca;
             14'h1e1 	:	val_out <= 16'h0bd0;
             14'h1e2 	:	val_out <= 16'h0bd6;
             14'h1e3 	:	val_out <= 16'h0bdc;
             14'h1e4 	:	val_out <= 16'h0be3;
             14'h1e5 	:	val_out <= 16'h0be9;
             14'h1e6 	:	val_out <= 16'h0bef;
             14'h1e7 	:	val_out <= 16'h0bf5;
             14'h1e8 	:	val_out <= 16'h0bfc;
             14'h1e9 	:	val_out <= 16'h0c02;
             14'h1ea 	:	val_out <= 16'h0c08;
             14'h1eb 	:	val_out <= 16'h0c0f;
             14'h1ec 	:	val_out <= 16'h0c15;
             14'h1ed 	:	val_out <= 16'h0c1b;
             14'h1ee 	:	val_out <= 16'h0c21;
             14'h1ef 	:	val_out <= 16'h0c28;
             14'h1f0 	:	val_out <= 16'h0c2e;
             14'h1f1 	:	val_out <= 16'h0c34;
             14'h1f2 	:	val_out <= 16'h0c3a;
             14'h1f3 	:	val_out <= 16'h0c41;
             14'h1f4 	:	val_out <= 16'h0c47;
             14'h1f5 	:	val_out <= 16'h0c4d;
             14'h1f6 	:	val_out <= 16'h0c54;
             14'h1f7 	:	val_out <= 16'h0c5a;
             14'h1f8 	:	val_out <= 16'h0c60;
             14'h1f9 	:	val_out <= 16'h0c66;
             14'h1fa 	:	val_out <= 16'h0c6d;
             14'h1fb 	:	val_out <= 16'h0c73;
             14'h1fc 	:	val_out <= 16'h0c79;
             14'h1fd 	:	val_out <= 16'h0c80;
             14'h1fe 	:	val_out <= 16'h0c86;
             14'h1ff 	:	val_out <= 16'h0c8c;
             14'h200 	:	val_out <= 16'h0c92;
             14'h201 	:	val_out <= 16'h0c99;
             14'h202 	:	val_out <= 16'h0c9f;
             14'h203 	:	val_out <= 16'h0ca5;
             14'h204 	:	val_out <= 16'h0cab;
             14'h205 	:	val_out <= 16'h0cb2;
             14'h206 	:	val_out <= 16'h0cb8;
             14'h207 	:	val_out <= 16'h0cbe;
             14'h208 	:	val_out <= 16'h0cc5;
             14'h209 	:	val_out <= 16'h0ccb;
             14'h20a 	:	val_out <= 16'h0cd1;
             14'h20b 	:	val_out <= 16'h0cd7;
             14'h20c 	:	val_out <= 16'h0cde;
             14'h20d 	:	val_out <= 16'h0ce4;
             14'h20e 	:	val_out <= 16'h0cea;
             14'h20f 	:	val_out <= 16'h0cf0;
             14'h210 	:	val_out <= 16'h0cf7;
             14'h211 	:	val_out <= 16'h0cfd;
             14'h212 	:	val_out <= 16'h0d03;
             14'h213 	:	val_out <= 16'h0d0a;
             14'h214 	:	val_out <= 16'h0d10;
             14'h215 	:	val_out <= 16'h0d16;
             14'h216 	:	val_out <= 16'h0d1c;
             14'h217 	:	val_out <= 16'h0d23;
             14'h218 	:	val_out <= 16'h0d29;
             14'h219 	:	val_out <= 16'h0d2f;
             14'h21a 	:	val_out <= 16'h0d35;
             14'h21b 	:	val_out <= 16'h0d3c;
             14'h21c 	:	val_out <= 16'h0d42;
             14'h21d 	:	val_out <= 16'h0d48;
             14'h21e 	:	val_out <= 16'h0d4f;
             14'h21f 	:	val_out <= 16'h0d55;
             14'h220 	:	val_out <= 16'h0d5b;
             14'h221 	:	val_out <= 16'h0d61;
             14'h222 	:	val_out <= 16'h0d68;
             14'h223 	:	val_out <= 16'h0d6e;
             14'h224 	:	val_out <= 16'h0d74;
             14'h225 	:	val_out <= 16'h0d7b;
             14'h226 	:	val_out <= 16'h0d81;
             14'h227 	:	val_out <= 16'h0d87;
             14'h228 	:	val_out <= 16'h0d8d;
             14'h229 	:	val_out <= 16'h0d94;
             14'h22a 	:	val_out <= 16'h0d9a;
             14'h22b 	:	val_out <= 16'h0da0;
             14'h22c 	:	val_out <= 16'h0da6;
             14'h22d 	:	val_out <= 16'h0dad;
             14'h22e 	:	val_out <= 16'h0db3;
             14'h22f 	:	val_out <= 16'h0db9;
             14'h230 	:	val_out <= 16'h0dc0;
             14'h231 	:	val_out <= 16'h0dc6;
             14'h232 	:	val_out <= 16'h0dcc;
             14'h233 	:	val_out <= 16'h0dd2;
             14'h234 	:	val_out <= 16'h0dd9;
             14'h235 	:	val_out <= 16'h0ddf;
             14'h236 	:	val_out <= 16'h0de5;
             14'h237 	:	val_out <= 16'h0deb;
             14'h238 	:	val_out <= 16'h0df2;
             14'h239 	:	val_out <= 16'h0df8;
             14'h23a 	:	val_out <= 16'h0dfe;
             14'h23b 	:	val_out <= 16'h0e05;
             14'h23c 	:	val_out <= 16'h0e0b;
             14'h23d 	:	val_out <= 16'h0e11;
             14'h23e 	:	val_out <= 16'h0e17;
             14'h23f 	:	val_out <= 16'h0e1e;
             14'h240 	:	val_out <= 16'h0e24;
             14'h241 	:	val_out <= 16'h0e2a;
             14'h242 	:	val_out <= 16'h0e30;
             14'h243 	:	val_out <= 16'h0e37;
             14'h244 	:	val_out <= 16'h0e3d;
             14'h245 	:	val_out <= 16'h0e43;
             14'h246 	:	val_out <= 16'h0e4a;
             14'h247 	:	val_out <= 16'h0e50;
             14'h248 	:	val_out <= 16'h0e56;
             14'h249 	:	val_out <= 16'h0e5c;
             14'h24a 	:	val_out <= 16'h0e63;
             14'h24b 	:	val_out <= 16'h0e69;
             14'h24c 	:	val_out <= 16'h0e6f;
             14'h24d 	:	val_out <= 16'h0e75;
             14'h24e 	:	val_out <= 16'h0e7c;
             14'h24f 	:	val_out <= 16'h0e82;
             14'h250 	:	val_out <= 16'h0e88;
             14'h251 	:	val_out <= 16'h0e8f;
             14'h252 	:	val_out <= 16'h0e95;
             14'h253 	:	val_out <= 16'h0e9b;
             14'h254 	:	val_out <= 16'h0ea1;
             14'h255 	:	val_out <= 16'h0ea8;
             14'h256 	:	val_out <= 16'h0eae;
             14'h257 	:	val_out <= 16'h0eb4;
             14'h258 	:	val_out <= 16'h0eba;
             14'h259 	:	val_out <= 16'h0ec1;
             14'h25a 	:	val_out <= 16'h0ec7;
             14'h25b 	:	val_out <= 16'h0ecd;
             14'h25c 	:	val_out <= 16'h0ed4;
             14'h25d 	:	val_out <= 16'h0eda;
             14'h25e 	:	val_out <= 16'h0ee0;
             14'h25f 	:	val_out <= 16'h0ee6;
             14'h260 	:	val_out <= 16'h0eed;
             14'h261 	:	val_out <= 16'h0ef3;
             14'h262 	:	val_out <= 16'h0ef9;
             14'h263 	:	val_out <= 16'h0eff;
             14'h264 	:	val_out <= 16'h0f06;
             14'h265 	:	val_out <= 16'h0f0c;
             14'h266 	:	val_out <= 16'h0f12;
             14'h267 	:	val_out <= 16'h0f19;
             14'h268 	:	val_out <= 16'h0f1f;
             14'h269 	:	val_out <= 16'h0f25;
             14'h26a 	:	val_out <= 16'h0f2b;
             14'h26b 	:	val_out <= 16'h0f32;
             14'h26c 	:	val_out <= 16'h0f38;
             14'h26d 	:	val_out <= 16'h0f3e;
             14'h26e 	:	val_out <= 16'h0f44;
             14'h26f 	:	val_out <= 16'h0f4b;
             14'h270 	:	val_out <= 16'h0f51;
             14'h271 	:	val_out <= 16'h0f57;
             14'h272 	:	val_out <= 16'h0f5e;
             14'h273 	:	val_out <= 16'h0f64;
             14'h274 	:	val_out <= 16'h0f6a;
             14'h275 	:	val_out <= 16'h0f70;
             14'h276 	:	val_out <= 16'h0f77;
             14'h277 	:	val_out <= 16'h0f7d;
             14'h278 	:	val_out <= 16'h0f83;
             14'h279 	:	val_out <= 16'h0f89;
             14'h27a 	:	val_out <= 16'h0f90;
             14'h27b 	:	val_out <= 16'h0f96;
             14'h27c 	:	val_out <= 16'h0f9c;
             14'h27d 	:	val_out <= 16'h0fa3;
             14'h27e 	:	val_out <= 16'h0fa9;
             14'h27f 	:	val_out <= 16'h0faf;
             14'h280 	:	val_out <= 16'h0fb5;
             14'h281 	:	val_out <= 16'h0fbc;
             14'h282 	:	val_out <= 16'h0fc2;
             14'h283 	:	val_out <= 16'h0fc8;
             14'h284 	:	val_out <= 16'h0fce;
             14'h285 	:	val_out <= 16'h0fd5;
             14'h286 	:	val_out <= 16'h0fdb;
             14'h287 	:	val_out <= 16'h0fe1;
             14'h288 	:	val_out <= 16'h0fe8;
             14'h289 	:	val_out <= 16'h0fee;
             14'h28a 	:	val_out <= 16'h0ff4;
             14'h28b 	:	val_out <= 16'h0ffa;
             14'h28c 	:	val_out <= 16'h1001;
             14'h28d 	:	val_out <= 16'h1007;
             14'h28e 	:	val_out <= 16'h100d;
             14'h28f 	:	val_out <= 16'h1013;
             14'h290 	:	val_out <= 16'h101a;
             14'h291 	:	val_out <= 16'h1020;
             14'h292 	:	val_out <= 16'h1026;
             14'h293 	:	val_out <= 16'h102d;
             14'h294 	:	val_out <= 16'h1033;
             14'h295 	:	val_out <= 16'h1039;
             14'h296 	:	val_out <= 16'h103f;
             14'h297 	:	val_out <= 16'h1046;
             14'h298 	:	val_out <= 16'h104c;
             14'h299 	:	val_out <= 16'h1052;
             14'h29a 	:	val_out <= 16'h1058;
             14'h29b 	:	val_out <= 16'h105f;
             14'h29c 	:	val_out <= 16'h1065;
             14'h29d 	:	val_out <= 16'h106b;
             14'h29e 	:	val_out <= 16'h1071;
             14'h29f 	:	val_out <= 16'h1078;
             14'h2a0 	:	val_out <= 16'h107e;
             14'h2a1 	:	val_out <= 16'h1084;
             14'h2a2 	:	val_out <= 16'h108b;
             14'h2a3 	:	val_out <= 16'h1091;
             14'h2a4 	:	val_out <= 16'h1097;
             14'h2a5 	:	val_out <= 16'h109d;
             14'h2a6 	:	val_out <= 16'h10a4;
             14'h2a7 	:	val_out <= 16'h10aa;
             14'h2a8 	:	val_out <= 16'h10b0;
             14'h2a9 	:	val_out <= 16'h10b6;
             14'h2aa 	:	val_out <= 16'h10bd;
             14'h2ab 	:	val_out <= 16'h10c3;
             14'h2ac 	:	val_out <= 16'h10c9;
             14'h2ad 	:	val_out <= 16'h10d0;
             14'h2ae 	:	val_out <= 16'h10d6;
             14'h2af 	:	val_out <= 16'h10dc;
             14'h2b0 	:	val_out <= 16'h10e2;
             14'h2b1 	:	val_out <= 16'h10e9;
             14'h2b2 	:	val_out <= 16'h10ef;
             14'h2b3 	:	val_out <= 16'h10f5;
             14'h2b4 	:	val_out <= 16'h10fb;
             14'h2b5 	:	val_out <= 16'h1102;
             14'h2b6 	:	val_out <= 16'h1108;
             14'h2b7 	:	val_out <= 16'h110e;
             14'h2b8 	:	val_out <= 16'h1114;
             14'h2b9 	:	val_out <= 16'h111b;
             14'h2ba 	:	val_out <= 16'h1121;
             14'h2bb 	:	val_out <= 16'h1127;
             14'h2bc 	:	val_out <= 16'h112e;
             14'h2bd 	:	val_out <= 16'h1134;
             14'h2be 	:	val_out <= 16'h113a;
             14'h2bf 	:	val_out <= 16'h1140;
             14'h2c0 	:	val_out <= 16'h1147;
             14'h2c1 	:	val_out <= 16'h114d;
             14'h2c2 	:	val_out <= 16'h1153;
             14'h2c3 	:	val_out <= 16'h1159;
             14'h2c4 	:	val_out <= 16'h1160;
             14'h2c5 	:	val_out <= 16'h1166;
             14'h2c6 	:	val_out <= 16'h116c;
             14'h2c7 	:	val_out <= 16'h1173;
             14'h2c8 	:	val_out <= 16'h1179;
             14'h2c9 	:	val_out <= 16'h117f;
             14'h2ca 	:	val_out <= 16'h1185;
             14'h2cb 	:	val_out <= 16'h118c;
             14'h2cc 	:	val_out <= 16'h1192;
             14'h2cd 	:	val_out <= 16'h1198;
             14'h2ce 	:	val_out <= 16'h119e;
             14'h2cf 	:	val_out <= 16'h11a5;
             14'h2d0 	:	val_out <= 16'h11ab;
             14'h2d1 	:	val_out <= 16'h11b1;
             14'h2d2 	:	val_out <= 16'h11b7;
             14'h2d3 	:	val_out <= 16'h11be;
             14'h2d4 	:	val_out <= 16'h11c4;
             14'h2d5 	:	val_out <= 16'h11ca;
             14'h2d6 	:	val_out <= 16'h11d1;
             14'h2d7 	:	val_out <= 16'h11d7;
             14'h2d8 	:	val_out <= 16'h11dd;
             14'h2d9 	:	val_out <= 16'h11e3;
             14'h2da 	:	val_out <= 16'h11ea;
             14'h2db 	:	val_out <= 16'h11f0;
             14'h2dc 	:	val_out <= 16'h11f6;
             14'h2dd 	:	val_out <= 16'h11fc;
             14'h2de 	:	val_out <= 16'h1203;
             14'h2df 	:	val_out <= 16'h1209;
             14'h2e0 	:	val_out <= 16'h120f;
             14'h2e1 	:	val_out <= 16'h1215;
             14'h2e2 	:	val_out <= 16'h121c;
             14'h2e3 	:	val_out <= 16'h1222;
             14'h2e4 	:	val_out <= 16'h1228;
             14'h2e5 	:	val_out <= 16'h122f;
             14'h2e6 	:	val_out <= 16'h1235;
             14'h2e7 	:	val_out <= 16'h123b;
             14'h2e8 	:	val_out <= 16'h1241;
             14'h2e9 	:	val_out <= 16'h1248;
             14'h2ea 	:	val_out <= 16'h124e;
             14'h2eb 	:	val_out <= 16'h1254;
             14'h2ec 	:	val_out <= 16'h125a;
             14'h2ed 	:	val_out <= 16'h1261;
             14'h2ee 	:	val_out <= 16'h1267;
             14'h2ef 	:	val_out <= 16'h126d;
             14'h2f0 	:	val_out <= 16'h1273;
             14'h2f1 	:	val_out <= 16'h127a;
             14'h2f2 	:	val_out <= 16'h1280;
             14'h2f3 	:	val_out <= 16'h1286;
             14'h2f4 	:	val_out <= 16'h128d;
             14'h2f5 	:	val_out <= 16'h1293;
             14'h2f6 	:	val_out <= 16'h1299;
             14'h2f7 	:	val_out <= 16'h129f;
             14'h2f8 	:	val_out <= 16'h12a6;
             14'h2f9 	:	val_out <= 16'h12ac;
             14'h2fa 	:	val_out <= 16'h12b2;
             14'h2fb 	:	val_out <= 16'h12b8;
             14'h2fc 	:	val_out <= 16'h12bf;
             14'h2fd 	:	val_out <= 16'h12c5;
             14'h2fe 	:	val_out <= 16'h12cb;
             14'h2ff 	:	val_out <= 16'h12d1;
             14'h300 	:	val_out <= 16'h12d8;
             14'h301 	:	val_out <= 16'h12de;
             14'h302 	:	val_out <= 16'h12e4;
             14'h303 	:	val_out <= 16'h12eb;
             14'h304 	:	val_out <= 16'h12f1;
             14'h305 	:	val_out <= 16'h12f7;
             14'h306 	:	val_out <= 16'h12fd;
             14'h307 	:	val_out <= 16'h1304;
             14'h308 	:	val_out <= 16'h130a;
             14'h309 	:	val_out <= 16'h1310;
             14'h30a 	:	val_out <= 16'h1316;
             14'h30b 	:	val_out <= 16'h131d;
             14'h30c 	:	val_out <= 16'h1323;
             14'h30d 	:	val_out <= 16'h1329;
             14'h30e 	:	val_out <= 16'h132f;
             14'h30f 	:	val_out <= 16'h1336;
             14'h310 	:	val_out <= 16'h133c;
             14'h311 	:	val_out <= 16'h1342;
             14'h312 	:	val_out <= 16'h1349;
             14'h313 	:	val_out <= 16'h134f;
             14'h314 	:	val_out <= 16'h1355;
             14'h315 	:	val_out <= 16'h135b;
             14'h316 	:	val_out <= 16'h1362;
             14'h317 	:	val_out <= 16'h1368;
             14'h318 	:	val_out <= 16'h136e;
             14'h319 	:	val_out <= 16'h1374;
             14'h31a 	:	val_out <= 16'h137b;
             14'h31b 	:	val_out <= 16'h1381;
             14'h31c 	:	val_out <= 16'h1387;
             14'h31d 	:	val_out <= 16'h138d;
             14'h31e 	:	val_out <= 16'h1394;
             14'h31f 	:	val_out <= 16'h139a;
             14'h320 	:	val_out <= 16'h13a0;
             14'h321 	:	val_out <= 16'h13a7;
             14'h322 	:	val_out <= 16'h13ad;
             14'h323 	:	val_out <= 16'h13b3;
             14'h324 	:	val_out <= 16'h13b9;
             14'h325 	:	val_out <= 16'h13c0;
             14'h326 	:	val_out <= 16'h13c6;
             14'h327 	:	val_out <= 16'h13cc;
             14'h328 	:	val_out <= 16'h13d2;
             14'h329 	:	val_out <= 16'h13d9;
             14'h32a 	:	val_out <= 16'h13df;
             14'h32b 	:	val_out <= 16'h13e5;
             14'h32c 	:	val_out <= 16'h13eb;
             14'h32d 	:	val_out <= 16'h13f2;
             14'h32e 	:	val_out <= 16'h13f8;
             14'h32f 	:	val_out <= 16'h13fe;
             14'h330 	:	val_out <= 16'h1404;
             14'h331 	:	val_out <= 16'h140b;
             14'h332 	:	val_out <= 16'h1411;
             14'h333 	:	val_out <= 16'h1417;
             14'h334 	:	val_out <= 16'h141e;
             14'h335 	:	val_out <= 16'h1424;
             14'h336 	:	val_out <= 16'h142a;
             14'h337 	:	val_out <= 16'h1430;
             14'h338 	:	val_out <= 16'h1437;
             14'h339 	:	val_out <= 16'h143d;
             14'h33a 	:	val_out <= 16'h1443;
             14'h33b 	:	val_out <= 16'h1449;
             14'h33c 	:	val_out <= 16'h1450;
             14'h33d 	:	val_out <= 16'h1456;
             14'h33e 	:	val_out <= 16'h145c;
             14'h33f 	:	val_out <= 16'h1462;
             14'h340 	:	val_out <= 16'h1469;
             14'h341 	:	val_out <= 16'h146f;
             14'h342 	:	val_out <= 16'h1475;
             14'h343 	:	val_out <= 16'h147b;
             14'h344 	:	val_out <= 16'h1482;
             14'h345 	:	val_out <= 16'h1488;
             14'h346 	:	val_out <= 16'h148e;
             14'h347 	:	val_out <= 16'h1495;
             14'h348 	:	val_out <= 16'h149b;
             14'h349 	:	val_out <= 16'h14a1;
             14'h34a 	:	val_out <= 16'h14a7;
             14'h34b 	:	val_out <= 16'h14ae;
             14'h34c 	:	val_out <= 16'h14b4;
             14'h34d 	:	val_out <= 16'h14ba;
             14'h34e 	:	val_out <= 16'h14c0;
             14'h34f 	:	val_out <= 16'h14c7;
             14'h350 	:	val_out <= 16'h14cd;
             14'h351 	:	val_out <= 16'h14d3;
             14'h352 	:	val_out <= 16'h14d9;
             14'h353 	:	val_out <= 16'h14e0;
             14'h354 	:	val_out <= 16'h14e6;
             14'h355 	:	val_out <= 16'h14ec;
             14'h356 	:	val_out <= 16'h14f2;
             14'h357 	:	val_out <= 16'h14f9;
             14'h358 	:	val_out <= 16'h14ff;
             14'h359 	:	val_out <= 16'h1505;
             14'h35a 	:	val_out <= 16'h150c;
             14'h35b 	:	val_out <= 16'h1512;
             14'h35c 	:	val_out <= 16'h1518;
             14'h35d 	:	val_out <= 16'h151e;
             14'h35e 	:	val_out <= 16'h1525;
             14'h35f 	:	val_out <= 16'h152b;
             14'h360 	:	val_out <= 16'h1531;
             14'h361 	:	val_out <= 16'h1537;
             14'h362 	:	val_out <= 16'h153e;
             14'h363 	:	val_out <= 16'h1544;
             14'h364 	:	val_out <= 16'h154a;
             14'h365 	:	val_out <= 16'h1550;
             14'h366 	:	val_out <= 16'h1557;
             14'h367 	:	val_out <= 16'h155d;
             14'h368 	:	val_out <= 16'h1563;
             14'h369 	:	val_out <= 16'h1569;
             14'h36a 	:	val_out <= 16'h1570;
             14'h36b 	:	val_out <= 16'h1576;
             14'h36c 	:	val_out <= 16'h157c;
             14'h36d 	:	val_out <= 16'h1582;
             14'h36e 	:	val_out <= 16'h1589;
             14'h36f 	:	val_out <= 16'h158f;
             14'h370 	:	val_out <= 16'h1595;
             14'h371 	:	val_out <= 16'h159c;
             14'h372 	:	val_out <= 16'h15a2;
             14'h373 	:	val_out <= 16'h15a8;
             14'h374 	:	val_out <= 16'h15ae;
             14'h375 	:	val_out <= 16'h15b5;
             14'h376 	:	val_out <= 16'h15bb;
             14'h377 	:	val_out <= 16'h15c1;
             14'h378 	:	val_out <= 16'h15c7;
             14'h379 	:	val_out <= 16'h15ce;
             14'h37a 	:	val_out <= 16'h15d4;
             14'h37b 	:	val_out <= 16'h15da;
             14'h37c 	:	val_out <= 16'h15e0;
             14'h37d 	:	val_out <= 16'h15e7;
             14'h37e 	:	val_out <= 16'h15ed;
             14'h37f 	:	val_out <= 16'h15f3;
             14'h380 	:	val_out <= 16'h15f9;
             14'h381 	:	val_out <= 16'h1600;
             14'h382 	:	val_out <= 16'h1606;
             14'h383 	:	val_out <= 16'h160c;
             14'h384 	:	val_out <= 16'h1612;
             14'h385 	:	val_out <= 16'h1619;
             14'h386 	:	val_out <= 16'h161f;
             14'h387 	:	val_out <= 16'h1625;
             14'h388 	:	val_out <= 16'h162c;
             14'h389 	:	val_out <= 16'h1632;
             14'h38a 	:	val_out <= 16'h1638;
             14'h38b 	:	val_out <= 16'h163e;
             14'h38c 	:	val_out <= 16'h1645;
             14'h38d 	:	val_out <= 16'h164b;
             14'h38e 	:	val_out <= 16'h1651;
             14'h38f 	:	val_out <= 16'h1657;
             14'h390 	:	val_out <= 16'h165e;
             14'h391 	:	val_out <= 16'h1664;
             14'h392 	:	val_out <= 16'h166a;
             14'h393 	:	val_out <= 16'h1670;
             14'h394 	:	val_out <= 16'h1677;
             14'h395 	:	val_out <= 16'h167d;
             14'h396 	:	val_out <= 16'h1683;
             14'h397 	:	val_out <= 16'h1689;
             14'h398 	:	val_out <= 16'h1690;
             14'h399 	:	val_out <= 16'h1696;
             14'h39a 	:	val_out <= 16'h169c;
             14'h39b 	:	val_out <= 16'h16a2;
             14'h39c 	:	val_out <= 16'h16a9;
             14'h39d 	:	val_out <= 16'h16af;
             14'h39e 	:	val_out <= 16'h16b5;
             14'h39f 	:	val_out <= 16'h16bb;
             14'h3a0 	:	val_out <= 16'h16c2;
             14'h3a1 	:	val_out <= 16'h16c8;
             14'h3a2 	:	val_out <= 16'h16ce;
             14'h3a3 	:	val_out <= 16'h16d5;
             14'h3a4 	:	val_out <= 16'h16db;
             14'h3a5 	:	val_out <= 16'h16e1;
             14'h3a6 	:	val_out <= 16'h16e7;
             14'h3a7 	:	val_out <= 16'h16ee;
             14'h3a8 	:	val_out <= 16'h16f4;
             14'h3a9 	:	val_out <= 16'h16fa;
             14'h3aa 	:	val_out <= 16'h1700;
             14'h3ab 	:	val_out <= 16'h1707;
             14'h3ac 	:	val_out <= 16'h170d;
             14'h3ad 	:	val_out <= 16'h1713;
             14'h3ae 	:	val_out <= 16'h1719;
             14'h3af 	:	val_out <= 16'h1720;
             14'h3b0 	:	val_out <= 16'h1726;
             14'h3b1 	:	val_out <= 16'h172c;
             14'h3b2 	:	val_out <= 16'h1732;
             14'h3b3 	:	val_out <= 16'h1739;
             14'h3b4 	:	val_out <= 16'h173f;
             14'h3b5 	:	val_out <= 16'h1745;
             14'h3b6 	:	val_out <= 16'h174b;
             14'h3b7 	:	val_out <= 16'h1752;
             14'h3b8 	:	val_out <= 16'h1758;
             14'h3b9 	:	val_out <= 16'h175e;
             14'h3ba 	:	val_out <= 16'h1764;
             14'h3bb 	:	val_out <= 16'h176b;
             14'h3bc 	:	val_out <= 16'h1771;
             14'h3bd 	:	val_out <= 16'h1777;
             14'h3be 	:	val_out <= 16'h177d;
             14'h3bf 	:	val_out <= 16'h1784;
             14'h3c0 	:	val_out <= 16'h178a;
             14'h3c1 	:	val_out <= 16'h1790;
             14'h3c2 	:	val_out <= 16'h1796;
             14'h3c3 	:	val_out <= 16'h179d;
             14'h3c4 	:	val_out <= 16'h17a3;
             14'h3c5 	:	val_out <= 16'h17a9;
             14'h3c6 	:	val_out <= 16'h17b0;
             14'h3c7 	:	val_out <= 16'h17b6;
             14'h3c8 	:	val_out <= 16'h17bc;
             14'h3c9 	:	val_out <= 16'h17c2;
             14'h3ca 	:	val_out <= 16'h17c9;
             14'h3cb 	:	val_out <= 16'h17cf;
             14'h3cc 	:	val_out <= 16'h17d5;
             14'h3cd 	:	val_out <= 16'h17db;
             14'h3ce 	:	val_out <= 16'h17e2;
             14'h3cf 	:	val_out <= 16'h17e8;
             14'h3d0 	:	val_out <= 16'h17ee;
             14'h3d1 	:	val_out <= 16'h17f4;
             14'h3d2 	:	val_out <= 16'h17fb;
             14'h3d3 	:	val_out <= 16'h1801;
             14'h3d4 	:	val_out <= 16'h1807;
             14'h3d5 	:	val_out <= 16'h180d;
             14'h3d6 	:	val_out <= 16'h1814;
             14'h3d7 	:	val_out <= 16'h181a;
             14'h3d8 	:	val_out <= 16'h1820;
             14'h3d9 	:	val_out <= 16'h1826;
             14'h3da 	:	val_out <= 16'h182d;
             14'h3db 	:	val_out <= 16'h1833;
             14'h3dc 	:	val_out <= 16'h1839;
             14'h3dd 	:	val_out <= 16'h183f;
             14'h3de 	:	val_out <= 16'h1846;
             14'h3df 	:	val_out <= 16'h184c;
             14'h3e0 	:	val_out <= 16'h1852;
             14'h3e1 	:	val_out <= 16'h1858;
             14'h3e2 	:	val_out <= 16'h185f;
             14'h3e3 	:	val_out <= 16'h1865;
             14'h3e4 	:	val_out <= 16'h186b;
             14'h3e5 	:	val_out <= 16'h1871;
             14'h3e6 	:	val_out <= 16'h1878;
             14'h3e7 	:	val_out <= 16'h187e;
             14'h3e8 	:	val_out <= 16'h1884;
             14'h3e9 	:	val_out <= 16'h188a;
             14'h3ea 	:	val_out <= 16'h1891;
             14'h3eb 	:	val_out <= 16'h1897;
             14'h3ec 	:	val_out <= 16'h189d;
             14'h3ed 	:	val_out <= 16'h18a3;
             14'h3ee 	:	val_out <= 16'h18aa;
             14'h3ef 	:	val_out <= 16'h18b0;
             14'h3f0 	:	val_out <= 16'h18b6;
             14'h3f1 	:	val_out <= 16'h18bc;
             14'h3f2 	:	val_out <= 16'h18c3;
             14'h3f3 	:	val_out <= 16'h18c9;
             14'h3f4 	:	val_out <= 16'h18cf;
             14'h3f5 	:	val_out <= 16'h18d5;
             14'h3f6 	:	val_out <= 16'h18dc;
             14'h3f7 	:	val_out <= 16'h18e2;
             14'h3f8 	:	val_out <= 16'h18e8;
             14'h3f9 	:	val_out <= 16'h18ef;
             14'h3fa 	:	val_out <= 16'h18f5;
             14'h3fb 	:	val_out <= 16'h18fb;
             14'h3fc 	:	val_out <= 16'h1901;
             14'h3fd 	:	val_out <= 16'h1908;
             14'h3fe 	:	val_out <= 16'h190e;
             14'h3ff 	:	val_out <= 16'h1914;
             14'h400 	:	val_out <= 16'h191a;
             14'h401 	:	val_out <= 16'h1921;
             14'h402 	:	val_out <= 16'h1927;
             14'h403 	:	val_out <= 16'h192d;
             14'h404 	:	val_out <= 16'h1933;
             14'h405 	:	val_out <= 16'h193a;
             14'h406 	:	val_out <= 16'h1940;
             14'h407 	:	val_out <= 16'h1946;
             14'h408 	:	val_out <= 16'h194c;
             14'h409 	:	val_out <= 16'h1953;
             14'h40a 	:	val_out <= 16'h1959;
             14'h40b 	:	val_out <= 16'h195f;
             14'h40c 	:	val_out <= 16'h1965;
             14'h40d 	:	val_out <= 16'h196c;
             14'h40e 	:	val_out <= 16'h1972;
             14'h40f 	:	val_out <= 16'h1978;
             14'h410 	:	val_out <= 16'h197e;
             14'h411 	:	val_out <= 16'h1985;
             14'h412 	:	val_out <= 16'h198b;
             14'h413 	:	val_out <= 16'h1991;
             14'h414 	:	val_out <= 16'h1997;
             14'h415 	:	val_out <= 16'h199e;
             14'h416 	:	val_out <= 16'h19a4;
             14'h417 	:	val_out <= 16'h19aa;
             14'h418 	:	val_out <= 16'h19b0;
             14'h419 	:	val_out <= 16'h19b7;
             14'h41a 	:	val_out <= 16'h19bd;
             14'h41b 	:	val_out <= 16'h19c3;
             14'h41c 	:	val_out <= 16'h19c9;
             14'h41d 	:	val_out <= 16'h19d0;
             14'h41e 	:	val_out <= 16'h19d6;
             14'h41f 	:	val_out <= 16'h19dc;
             14'h420 	:	val_out <= 16'h19e2;
             14'h421 	:	val_out <= 16'h19e9;
             14'h422 	:	val_out <= 16'h19ef;
             14'h423 	:	val_out <= 16'h19f5;
             14'h424 	:	val_out <= 16'h19fb;
             14'h425 	:	val_out <= 16'h1a02;
             14'h426 	:	val_out <= 16'h1a08;
             14'h427 	:	val_out <= 16'h1a0e;
             14'h428 	:	val_out <= 16'h1a14;
             14'h429 	:	val_out <= 16'h1a1b;
             14'h42a 	:	val_out <= 16'h1a21;
             14'h42b 	:	val_out <= 16'h1a27;
             14'h42c 	:	val_out <= 16'h1a2d;
             14'h42d 	:	val_out <= 16'h1a34;
             14'h42e 	:	val_out <= 16'h1a3a;
             14'h42f 	:	val_out <= 16'h1a40;
             14'h430 	:	val_out <= 16'h1a46;
             14'h431 	:	val_out <= 16'h1a4d;
             14'h432 	:	val_out <= 16'h1a53;
             14'h433 	:	val_out <= 16'h1a59;
             14'h434 	:	val_out <= 16'h1a5f;
             14'h435 	:	val_out <= 16'h1a66;
             14'h436 	:	val_out <= 16'h1a6c;
             14'h437 	:	val_out <= 16'h1a72;
             14'h438 	:	val_out <= 16'h1a78;
             14'h439 	:	val_out <= 16'h1a7f;
             14'h43a 	:	val_out <= 16'h1a85;
             14'h43b 	:	val_out <= 16'h1a8b;
             14'h43c 	:	val_out <= 16'h1a91;
             14'h43d 	:	val_out <= 16'h1a98;
             14'h43e 	:	val_out <= 16'h1a9e;
             14'h43f 	:	val_out <= 16'h1aa4;
             14'h440 	:	val_out <= 16'h1aaa;
             14'h441 	:	val_out <= 16'h1ab1;
             14'h442 	:	val_out <= 16'h1ab7;
             14'h443 	:	val_out <= 16'h1abd;
             14'h444 	:	val_out <= 16'h1ac3;
             14'h445 	:	val_out <= 16'h1aca;
             14'h446 	:	val_out <= 16'h1ad0;
             14'h447 	:	val_out <= 16'h1ad6;
             14'h448 	:	val_out <= 16'h1adc;
             14'h449 	:	val_out <= 16'h1ae3;
             14'h44a 	:	val_out <= 16'h1ae9;
             14'h44b 	:	val_out <= 16'h1aef;
             14'h44c 	:	val_out <= 16'h1af5;
             14'h44d 	:	val_out <= 16'h1afc;
             14'h44e 	:	val_out <= 16'h1b02;
             14'h44f 	:	val_out <= 16'h1b08;
             14'h450 	:	val_out <= 16'h1b0e;
             14'h451 	:	val_out <= 16'h1b15;
             14'h452 	:	val_out <= 16'h1b1b;
             14'h453 	:	val_out <= 16'h1b21;
             14'h454 	:	val_out <= 16'h1b27;
             14'h455 	:	val_out <= 16'h1b2e;
             14'h456 	:	val_out <= 16'h1b34;
             14'h457 	:	val_out <= 16'h1b3a;
             14'h458 	:	val_out <= 16'h1b40;
             14'h459 	:	val_out <= 16'h1b47;
             14'h45a 	:	val_out <= 16'h1b4d;
             14'h45b 	:	val_out <= 16'h1b53;
             14'h45c 	:	val_out <= 16'h1b59;
             14'h45d 	:	val_out <= 16'h1b60;
             14'h45e 	:	val_out <= 16'h1b66;
             14'h45f 	:	val_out <= 16'h1b6c;
             14'h460 	:	val_out <= 16'h1b72;
             14'h461 	:	val_out <= 16'h1b79;
             14'h462 	:	val_out <= 16'h1b7f;
             14'h463 	:	val_out <= 16'h1b85;
             14'h464 	:	val_out <= 16'h1b8b;
             14'h465 	:	val_out <= 16'h1b92;
             14'h466 	:	val_out <= 16'h1b98;
             14'h467 	:	val_out <= 16'h1b9e;
             14'h468 	:	val_out <= 16'h1ba4;
             14'h469 	:	val_out <= 16'h1baa;
             14'h46a 	:	val_out <= 16'h1bb1;
             14'h46b 	:	val_out <= 16'h1bb7;
             14'h46c 	:	val_out <= 16'h1bbd;
             14'h46d 	:	val_out <= 16'h1bc3;
             14'h46e 	:	val_out <= 16'h1bca;
             14'h46f 	:	val_out <= 16'h1bd0;
             14'h470 	:	val_out <= 16'h1bd6;
             14'h471 	:	val_out <= 16'h1bdc;
             14'h472 	:	val_out <= 16'h1be3;
             14'h473 	:	val_out <= 16'h1be9;
             14'h474 	:	val_out <= 16'h1bef;
             14'h475 	:	val_out <= 16'h1bf5;
             14'h476 	:	val_out <= 16'h1bfc;
             14'h477 	:	val_out <= 16'h1c02;
             14'h478 	:	val_out <= 16'h1c08;
             14'h479 	:	val_out <= 16'h1c0e;
             14'h47a 	:	val_out <= 16'h1c15;
             14'h47b 	:	val_out <= 16'h1c1b;
             14'h47c 	:	val_out <= 16'h1c21;
             14'h47d 	:	val_out <= 16'h1c27;
             14'h47e 	:	val_out <= 16'h1c2e;
             14'h47f 	:	val_out <= 16'h1c34;
             14'h480 	:	val_out <= 16'h1c3a;
             14'h481 	:	val_out <= 16'h1c40;
             14'h482 	:	val_out <= 16'h1c47;
             14'h483 	:	val_out <= 16'h1c4d;
             14'h484 	:	val_out <= 16'h1c53;
             14'h485 	:	val_out <= 16'h1c59;
             14'h486 	:	val_out <= 16'h1c60;
             14'h487 	:	val_out <= 16'h1c66;
             14'h488 	:	val_out <= 16'h1c6c;
             14'h489 	:	val_out <= 16'h1c72;
             14'h48a 	:	val_out <= 16'h1c79;
             14'h48b 	:	val_out <= 16'h1c7f;
             14'h48c 	:	val_out <= 16'h1c85;
             14'h48d 	:	val_out <= 16'h1c8b;
             14'h48e 	:	val_out <= 16'h1c92;
             14'h48f 	:	val_out <= 16'h1c98;
             14'h490 	:	val_out <= 16'h1c9e;
             14'h491 	:	val_out <= 16'h1ca4;
             14'h492 	:	val_out <= 16'h1cab;
             14'h493 	:	val_out <= 16'h1cb1;
             14'h494 	:	val_out <= 16'h1cb7;
             14'h495 	:	val_out <= 16'h1cbd;
             14'h496 	:	val_out <= 16'h1cc4;
             14'h497 	:	val_out <= 16'h1cca;
             14'h498 	:	val_out <= 16'h1cd0;
             14'h499 	:	val_out <= 16'h1cd6;
             14'h49a 	:	val_out <= 16'h1cdc;
             14'h49b 	:	val_out <= 16'h1ce3;
             14'h49c 	:	val_out <= 16'h1ce9;
             14'h49d 	:	val_out <= 16'h1cef;
             14'h49e 	:	val_out <= 16'h1cf5;
             14'h49f 	:	val_out <= 16'h1cfc;
             14'h4a0 	:	val_out <= 16'h1d02;
             14'h4a1 	:	val_out <= 16'h1d08;
             14'h4a2 	:	val_out <= 16'h1d0e;
             14'h4a3 	:	val_out <= 16'h1d15;
             14'h4a4 	:	val_out <= 16'h1d1b;
             14'h4a5 	:	val_out <= 16'h1d21;
             14'h4a6 	:	val_out <= 16'h1d27;
             14'h4a7 	:	val_out <= 16'h1d2e;
             14'h4a8 	:	val_out <= 16'h1d34;
             14'h4a9 	:	val_out <= 16'h1d3a;
             14'h4aa 	:	val_out <= 16'h1d40;
             14'h4ab 	:	val_out <= 16'h1d47;
             14'h4ac 	:	val_out <= 16'h1d4d;
             14'h4ad 	:	val_out <= 16'h1d53;
             14'h4ae 	:	val_out <= 16'h1d59;
             14'h4af 	:	val_out <= 16'h1d60;
             14'h4b0 	:	val_out <= 16'h1d66;
             14'h4b1 	:	val_out <= 16'h1d6c;
             14'h4b2 	:	val_out <= 16'h1d72;
             14'h4b3 	:	val_out <= 16'h1d79;
             14'h4b4 	:	val_out <= 16'h1d7f;
             14'h4b5 	:	val_out <= 16'h1d85;
             14'h4b6 	:	val_out <= 16'h1d8b;
             14'h4b7 	:	val_out <= 16'h1d92;
             14'h4b8 	:	val_out <= 16'h1d98;
             14'h4b9 	:	val_out <= 16'h1d9e;
             14'h4ba 	:	val_out <= 16'h1da4;
             14'h4bb 	:	val_out <= 16'h1daa;
             14'h4bc 	:	val_out <= 16'h1db1;
             14'h4bd 	:	val_out <= 16'h1db7;
             14'h4be 	:	val_out <= 16'h1dbd;
             14'h4bf 	:	val_out <= 16'h1dc3;
             14'h4c0 	:	val_out <= 16'h1dca;
             14'h4c1 	:	val_out <= 16'h1dd0;
             14'h4c2 	:	val_out <= 16'h1dd6;
             14'h4c3 	:	val_out <= 16'h1ddc;
             14'h4c4 	:	val_out <= 16'h1de3;
             14'h4c5 	:	val_out <= 16'h1de9;
             14'h4c6 	:	val_out <= 16'h1def;
             14'h4c7 	:	val_out <= 16'h1df5;
             14'h4c8 	:	val_out <= 16'h1dfc;
             14'h4c9 	:	val_out <= 16'h1e02;
             14'h4ca 	:	val_out <= 16'h1e08;
             14'h4cb 	:	val_out <= 16'h1e0e;
             14'h4cc 	:	val_out <= 16'h1e15;
             14'h4cd 	:	val_out <= 16'h1e1b;
             14'h4ce 	:	val_out <= 16'h1e21;
             14'h4cf 	:	val_out <= 16'h1e27;
             14'h4d0 	:	val_out <= 16'h1e2e;
             14'h4d1 	:	val_out <= 16'h1e34;
             14'h4d2 	:	val_out <= 16'h1e3a;
             14'h4d3 	:	val_out <= 16'h1e40;
             14'h4d4 	:	val_out <= 16'h1e46;
             14'h4d5 	:	val_out <= 16'h1e4d;
             14'h4d6 	:	val_out <= 16'h1e53;
             14'h4d7 	:	val_out <= 16'h1e59;
             14'h4d8 	:	val_out <= 16'h1e5f;
             14'h4d9 	:	val_out <= 16'h1e66;
             14'h4da 	:	val_out <= 16'h1e6c;
             14'h4db 	:	val_out <= 16'h1e72;
             14'h4dc 	:	val_out <= 16'h1e78;
             14'h4dd 	:	val_out <= 16'h1e7f;
             14'h4de 	:	val_out <= 16'h1e85;
             14'h4df 	:	val_out <= 16'h1e8b;
             14'h4e0 	:	val_out <= 16'h1e91;
             14'h4e1 	:	val_out <= 16'h1e98;
             14'h4e2 	:	val_out <= 16'h1e9e;
             14'h4e3 	:	val_out <= 16'h1ea4;
             14'h4e4 	:	val_out <= 16'h1eaa;
             14'h4e5 	:	val_out <= 16'h1eb1;
             14'h4e6 	:	val_out <= 16'h1eb7;
             14'h4e7 	:	val_out <= 16'h1ebd;
             14'h4e8 	:	val_out <= 16'h1ec3;
             14'h4e9 	:	val_out <= 16'h1ec9;
             14'h4ea 	:	val_out <= 16'h1ed0;
             14'h4eb 	:	val_out <= 16'h1ed6;
             14'h4ec 	:	val_out <= 16'h1edc;
             14'h4ed 	:	val_out <= 16'h1ee2;
             14'h4ee 	:	val_out <= 16'h1ee9;
             14'h4ef 	:	val_out <= 16'h1eef;
             14'h4f0 	:	val_out <= 16'h1ef5;
             14'h4f1 	:	val_out <= 16'h1efb;
             14'h4f2 	:	val_out <= 16'h1f02;
             14'h4f3 	:	val_out <= 16'h1f08;
             14'h4f4 	:	val_out <= 16'h1f0e;
             14'h4f5 	:	val_out <= 16'h1f14;
             14'h4f6 	:	val_out <= 16'h1f1b;
             14'h4f7 	:	val_out <= 16'h1f21;
             14'h4f8 	:	val_out <= 16'h1f27;
             14'h4f9 	:	val_out <= 16'h1f2d;
             14'h4fa 	:	val_out <= 16'h1f34;
             14'h4fb 	:	val_out <= 16'h1f3a;
             14'h4fc 	:	val_out <= 16'h1f40;
             14'h4fd 	:	val_out <= 16'h1f46;
             14'h4fe 	:	val_out <= 16'h1f4c;
             14'h4ff 	:	val_out <= 16'h1f53;
             14'h500 	:	val_out <= 16'h1f59;
             14'h501 	:	val_out <= 16'h1f5f;
             14'h502 	:	val_out <= 16'h1f65;
             14'h503 	:	val_out <= 16'h1f6c;
             14'h504 	:	val_out <= 16'h1f72;
             14'h505 	:	val_out <= 16'h1f78;
             14'h506 	:	val_out <= 16'h1f7e;
             14'h507 	:	val_out <= 16'h1f85;
             14'h508 	:	val_out <= 16'h1f8b;
             14'h509 	:	val_out <= 16'h1f91;
             14'h50a 	:	val_out <= 16'h1f97;
             14'h50b 	:	val_out <= 16'h1f9e;
             14'h50c 	:	val_out <= 16'h1fa4;
             14'h50d 	:	val_out <= 16'h1faa;
             14'h50e 	:	val_out <= 16'h1fb0;
             14'h50f 	:	val_out <= 16'h1fb6;
             14'h510 	:	val_out <= 16'h1fbd;
             14'h511 	:	val_out <= 16'h1fc3;
             14'h512 	:	val_out <= 16'h1fc9;
             14'h513 	:	val_out <= 16'h1fcf;
             14'h514 	:	val_out <= 16'h1fd6;
             14'h515 	:	val_out <= 16'h1fdc;
             14'h516 	:	val_out <= 16'h1fe2;
             14'h517 	:	val_out <= 16'h1fe8;
             14'h518 	:	val_out <= 16'h1fef;
             14'h519 	:	val_out <= 16'h1ff5;
             14'h51a 	:	val_out <= 16'h1ffb;
             14'h51b 	:	val_out <= 16'h2001;
             14'h51c 	:	val_out <= 16'h2007;
             14'h51d 	:	val_out <= 16'h200e;
             14'h51e 	:	val_out <= 16'h2014;
             14'h51f 	:	val_out <= 16'h201a;
             14'h520 	:	val_out <= 16'h2020;
             14'h521 	:	val_out <= 16'h2027;
             14'h522 	:	val_out <= 16'h202d;
             14'h523 	:	val_out <= 16'h2033;
             14'h524 	:	val_out <= 16'h2039;
             14'h525 	:	val_out <= 16'h2040;
             14'h526 	:	val_out <= 16'h2046;
             14'h527 	:	val_out <= 16'h204c;
             14'h528 	:	val_out <= 16'h2052;
             14'h529 	:	val_out <= 16'h2059;
             14'h52a 	:	val_out <= 16'h205f;
             14'h52b 	:	val_out <= 16'h2065;
             14'h52c 	:	val_out <= 16'h206b;
             14'h52d 	:	val_out <= 16'h2071;
             14'h52e 	:	val_out <= 16'h2078;
             14'h52f 	:	val_out <= 16'h207e;
             14'h530 	:	val_out <= 16'h2084;
             14'h531 	:	val_out <= 16'h208a;
             14'h532 	:	val_out <= 16'h2091;
             14'h533 	:	val_out <= 16'h2097;
             14'h534 	:	val_out <= 16'h209d;
             14'h535 	:	val_out <= 16'h20a3;
             14'h536 	:	val_out <= 16'h20aa;
             14'h537 	:	val_out <= 16'h20b0;
             14'h538 	:	val_out <= 16'h20b6;
             14'h539 	:	val_out <= 16'h20bc;
             14'h53a 	:	val_out <= 16'h20c2;
             14'h53b 	:	val_out <= 16'h20c9;
             14'h53c 	:	val_out <= 16'h20cf;
             14'h53d 	:	val_out <= 16'h20d5;
             14'h53e 	:	val_out <= 16'h20db;
             14'h53f 	:	val_out <= 16'h20e2;
             14'h540 	:	val_out <= 16'h20e8;
             14'h541 	:	val_out <= 16'h20ee;
             14'h542 	:	val_out <= 16'h20f4;
             14'h543 	:	val_out <= 16'h20fb;
             14'h544 	:	val_out <= 16'h2101;
             14'h545 	:	val_out <= 16'h2107;
             14'h546 	:	val_out <= 16'h210d;
             14'h547 	:	val_out <= 16'h2113;
             14'h548 	:	val_out <= 16'h211a;
             14'h549 	:	val_out <= 16'h2120;
             14'h54a 	:	val_out <= 16'h2126;
             14'h54b 	:	val_out <= 16'h212c;
             14'h54c 	:	val_out <= 16'h2133;
             14'h54d 	:	val_out <= 16'h2139;
             14'h54e 	:	val_out <= 16'h213f;
             14'h54f 	:	val_out <= 16'h2145;
             14'h550 	:	val_out <= 16'h214c;
             14'h551 	:	val_out <= 16'h2152;
             14'h552 	:	val_out <= 16'h2158;
             14'h553 	:	val_out <= 16'h215e;
             14'h554 	:	val_out <= 16'h2164;
             14'h555 	:	val_out <= 16'h216b;
             14'h556 	:	val_out <= 16'h2171;
             14'h557 	:	val_out <= 16'h2177;
             14'h558 	:	val_out <= 16'h217d;
             14'h559 	:	val_out <= 16'h2184;
             14'h55a 	:	val_out <= 16'h218a;
             14'h55b 	:	val_out <= 16'h2190;
             14'h55c 	:	val_out <= 16'h2196;
             14'h55d 	:	val_out <= 16'h219d;
             14'h55e 	:	val_out <= 16'h21a3;
             14'h55f 	:	val_out <= 16'h21a9;
             14'h560 	:	val_out <= 16'h21af;
             14'h561 	:	val_out <= 16'h21b5;
             14'h562 	:	val_out <= 16'h21bc;
             14'h563 	:	val_out <= 16'h21c2;
             14'h564 	:	val_out <= 16'h21c8;
             14'h565 	:	val_out <= 16'h21ce;
             14'h566 	:	val_out <= 16'h21d5;
             14'h567 	:	val_out <= 16'h21db;
             14'h568 	:	val_out <= 16'h21e1;
             14'h569 	:	val_out <= 16'h21e7;
             14'h56a 	:	val_out <= 16'h21ee;
             14'h56b 	:	val_out <= 16'h21f4;
             14'h56c 	:	val_out <= 16'h21fa;
             14'h56d 	:	val_out <= 16'h2200;
             14'h56e 	:	val_out <= 16'h2206;
             14'h56f 	:	val_out <= 16'h220d;
             14'h570 	:	val_out <= 16'h2213;
             14'h571 	:	val_out <= 16'h2219;
             14'h572 	:	val_out <= 16'h221f;
             14'h573 	:	val_out <= 16'h2226;
             14'h574 	:	val_out <= 16'h222c;
             14'h575 	:	val_out <= 16'h2232;
             14'h576 	:	val_out <= 16'h2238;
             14'h577 	:	val_out <= 16'h223e;
             14'h578 	:	val_out <= 16'h2245;
             14'h579 	:	val_out <= 16'h224b;
             14'h57a 	:	val_out <= 16'h2251;
             14'h57b 	:	val_out <= 16'h2257;
             14'h57c 	:	val_out <= 16'h225e;
             14'h57d 	:	val_out <= 16'h2264;
             14'h57e 	:	val_out <= 16'h226a;
             14'h57f 	:	val_out <= 16'h2270;
             14'h580 	:	val_out <= 16'h2276;
             14'h581 	:	val_out <= 16'h227d;
             14'h582 	:	val_out <= 16'h2283;
             14'h583 	:	val_out <= 16'h2289;
             14'h584 	:	val_out <= 16'h228f;
             14'h585 	:	val_out <= 16'h2296;
             14'h586 	:	val_out <= 16'h229c;
             14'h587 	:	val_out <= 16'h22a2;
             14'h588 	:	val_out <= 16'h22a8;
             14'h589 	:	val_out <= 16'h22af;
             14'h58a 	:	val_out <= 16'h22b5;
             14'h58b 	:	val_out <= 16'h22bb;
             14'h58c 	:	val_out <= 16'h22c1;
             14'h58d 	:	val_out <= 16'h22c7;
             14'h58e 	:	val_out <= 16'h22ce;
             14'h58f 	:	val_out <= 16'h22d4;
             14'h590 	:	val_out <= 16'h22da;
             14'h591 	:	val_out <= 16'h22e0;
             14'h592 	:	val_out <= 16'h22e7;
             14'h593 	:	val_out <= 16'h22ed;
             14'h594 	:	val_out <= 16'h22f3;
             14'h595 	:	val_out <= 16'h22f9;
             14'h596 	:	val_out <= 16'h22ff;
             14'h597 	:	val_out <= 16'h2306;
             14'h598 	:	val_out <= 16'h230c;
             14'h599 	:	val_out <= 16'h2312;
             14'h59a 	:	val_out <= 16'h2318;
             14'h59b 	:	val_out <= 16'h231f;
             14'h59c 	:	val_out <= 16'h2325;
             14'h59d 	:	val_out <= 16'h232b;
             14'h59e 	:	val_out <= 16'h2331;
             14'h59f 	:	val_out <= 16'h2337;
             14'h5a0 	:	val_out <= 16'h233e;
             14'h5a1 	:	val_out <= 16'h2344;
             14'h5a2 	:	val_out <= 16'h234a;
             14'h5a3 	:	val_out <= 16'h2350;
             14'h5a4 	:	val_out <= 16'h2357;
             14'h5a5 	:	val_out <= 16'h235d;
             14'h5a6 	:	val_out <= 16'h2363;
             14'h5a7 	:	val_out <= 16'h2369;
             14'h5a8 	:	val_out <= 16'h236f;
             14'h5a9 	:	val_out <= 16'h2376;
             14'h5aa 	:	val_out <= 16'h237c;
             14'h5ab 	:	val_out <= 16'h2382;
             14'h5ac 	:	val_out <= 16'h2388;
             14'h5ad 	:	val_out <= 16'h238f;
             14'h5ae 	:	val_out <= 16'h2395;
             14'h5af 	:	val_out <= 16'h239b;
             14'h5b0 	:	val_out <= 16'h23a1;
             14'h5b1 	:	val_out <= 16'h23a7;
             14'h5b2 	:	val_out <= 16'h23ae;
             14'h5b3 	:	val_out <= 16'h23b4;
             14'h5b4 	:	val_out <= 16'h23ba;
             14'h5b5 	:	val_out <= 16'h23c0;
             14'h5b6 	:	val_out <= 16'h23c7;
             14'h5b7 	:	val_out <= 16'h23cd;
             14'h5b8 	:	val_out <= 16'h23d3;
             14'h5b9 	:	val_out <= 16'h23d9;
             14'h5ba 	:	val_out <= 16'h23df;
             14'h5bb 	:	val_out <= 16'h23e6;
             14'h5bc 	:	val_out <= 16'h23ec;
             14'h5bd 	:	val_out <= 16'h23f2;
             14'h5be 	:	val_out <= 16'h23f8;
             14'h5bf 	:	val_out <= 16'h23ff;
             14'h5c0 	:	val_out <= 16'h2405;
             14'h5c1 	:	val_out <= 16'h240b;
             14'h5c2 	:	val_out <= 16'h2411;
             14'h5c3 	:	val_out <= 16'h2417;
             14'h5c4 	:	val_out <= 16'h241e;
             14'h5c5 	:	val_out <= 16'h2424;
             14'h5c6 	:	val_out <= 16'h242a;
             14'h5c7 	:	val_out <= 16'h2430;
             14'h5c8 	:	val_out <= 16'h2437;
             14'h5c9 	:	val_out <= 16'h243d;
             14'h5ca 	:	val_out <= 16'h2443;
             14'h5cb 	:	val_out <= 16'h2449;
             14'h5cc 	:	val_out <= 16'h244f;
             14'h5cd 	:	val_out <= 16'h2456;
             14'h5ce 	:	val_out <= 16'h245c;
             14'h5cf 	:	val_out <= 16'h2462;
             14'h5d0 	:	val_out <= 16'h2468;
             14'h5d1 	:	val_out <= 16'h246f;
             14'h5d2 	:	val_out <= 16'h2475;
             14'h5d3 	:	val_out <= 16'h247b;
             14'h5d4 	:	val_out <= 16'h2481;
             14'h5d5 	:	val_out <= 16'h2487;
             14'h5d6 	:	val_out <= 16'h248e;
             14'h5d7 	:	val_out <= 16'h2494;
             14'h5d8 	:	val_out <= 16'h249a;
             14'h5d9 	:	val_out <= 16'h24a0;
             14'h5da 	:	val_out <= 16'h24a6;
             14'h5db 	:	val_out <= 16'h24ad;
             14'h5dc 	:	val_out <= 16'h24b3;
             14'h5dd 	:	val_out <= 16'h24b9;
             14'h5de 	:	val_out <= 16'h24bf;
             14'h5df 	:	val_out <= 16'h24c6;
             14'h5e0 	:	val_out <= 16'h24cc;
             14'h5e1 	:	val_out <= 16'h24d2;
             14'h5e2 	:	val_out <= 16'h24d8;
             14'h5e3 	:	val_out <= 16'h24de;
             14'h5e4 	:	val_out <= 16'h24e5;
             14'h5e5 	:	val_out <= 16'h24eb;
             14'h5e6 	:	val_out <= 16'h24f1;
             14'h5e7 	:	val_out <= 16'h24f7;
             14'h5e8 	:	val_out <= 16'h24fe;
             14'h5e9 	:	val_out <= 16'h2504;
             14'h5ea 	:	val_out <= 16'h250a;
             14'h5eb 	:	val_out <= 16'h2510;
             14'h5ec 	:	val_out <= 16'h2516;
             14'h5ed 	:	val_out <= 16'h251d;
             14'h5ee 	:	val_out <= 16'h2523;
             14'h5ef 	:	val_out <= 16'h2529;
             14'h5f0 	:	val_out <= 16'h252f;
             14'h5f1 	:	val_out <= 16'h2535;
             14'h5f2 	:	val_out <= 16'h253c;
             14'h5f3 	:	val_out <= 16'h2542;
             14'h5f4 	:	val_out <= 16'h2548;
             14'h5f5 	:	val_out <= 16'h254e;
             14'h5f6 	:	val_out <= 16'h2555;
             14'h5f7 	:	val_out <= 16'h255b;
             14'h5f8 	:	val_out <= 16'h2561;
             14'h5f9 	:	val_out <= 16'h2567;
             14'h5fa 	:	val_out <= 16'h256d;
             14'h5fb 	:	val_out <= 16'h2574;
             14'h5fc 	:	val_out <= 16'h257a;
             14'h5fd 	:	val_out <= 16'h2580;
             14'h5fe 	:	val_out <= 16'h2586;
             14'h5ff 	:	val_out <= 16'h258d;
             14'h600 	:	val_out <= 16'h2593;
             14'h601 	:	val_out <= 16'h2599;
             14'h602 	:	val_out <= 16'h259f;
             14'h603 	:	val_out <= 16'h25a5;
             14'h604 	:	val_out <= 16'h25ac;
             14'h605 	:	val_out <= 16'h25b2;
             14'h606 	:	val_out <= 16'h25b8;
             14'h607 	:	val_out <= 16'h25be;
             14'h608 	:	val_out <= 16'h25c4;
             14'h609 	:	val_out <= 16'h25cb;
             14'h60a 	:	val_out <= 16'h25d1;
             14'h60b 	:	val_out <= 16'h25d7;
             14'h60c 	:	val_out <= 16'h25dd;
             14'h60d 	:	val_out <= 16'h25e4;
             14'h60e 	:	val_out <= 16'h25ea;
             14'h60f 	:	val_out <= 16'h25f0;
             14'h610 	:	val_out <= 16'h25f6;
             14'h611 	:	val_out <= 16'h25fc;
             14'h612 	:	val_out <= 16'h2603;
             14'h613 	:	val_out <= 16'h2609;
             14'h614 	:	val_out <= 16'h260f;
             14'h615 	:	val_out <= 16'h2615;
             14'h616 	:	val_out <= 16'h261b;
             14'h617 	:	val_out <= 16'h2622;
             14'h618 	:	val_out <= 16'h2628;
             14'h619 	:	val_out <= 16'h262e;
             14'h61a 	:	val_out <= 16'h2634;
             14'h61b 	:	val_out <= 16'h263b;
             14'h61c 	:	val_out <= 16'h2641;
             14'h61d 	:	val_out <= 16'h2647;
             14'h61e 	:	val_out <= 16'h264d;
             14'h61f 	:	val_out <= 16'h2653;
             14'h620 	:	val_out <= 16'h265a;
             14'h621 	:	val_out <= 16'h2660;
             14'h622 	:	val_out <= 16'h2666;
             14'h623 	:	val_out <= 16'h266c;
             14'h624 	:	val_out <= 16'h2672;
             14'h625 	:	val_out <= 16'h2679;
             14'h626 	:	val_out <= 16'h267f;
             14'h627 	:	val_out <= 16'h2685;
             14'h628 	:	val_out <= 16'h268b;
             14'h629 	:	val_out <= 16'h2691;
             14'h62a 	:	val_out <= 16'h2698;
             14'h62b 	:	val_out <= 16'h269e;
             14'h62c 	:	val_out <= 16'h26a4;
             14'h62d 	:	val_out <= 16'h26aa;
             14'h62e 	:	val_out <= 16'h26b1;
             14'h62f 	:	val_out <= 16'h26b7;
             14'h630 	:	val_out <= 16'h26bd;
             14'h631 	:	val_out <= 16'h26c3;
             14'h632 	:	val_out <= 16'h26c9;
             14'h633 	:	val_out <= 16'h26d0;
             14'h634 	:	val_out <= 16'h26d6;
             14'h635 	:	val_out <= 16'h26dc;
             14'h636 	:	val_out <= 16'h26e2;
             14'h637 	:	val_out <= 16'h26e8;
             14'h638 	:	val_out <= 16'h26ef;
             14'h639 	:	val_out <= 16'h26f5;
             14'h63a 	:	val_out <= 16'h26fb;
             14'h63b 	:	val_out <= 16'h2701;
             14'h63c 	:	val_out <= 16'h2707;
             14'h63d 	:	val_out <= 16'h270e;
             14'h63e 	:	val_out <= 16'h2714;
             14'h63f 	:	val_out <= 16'h271a;
             14'h640 	:	val_out <= 16'h2720;
             14'h641 	:	val_out <= 16'h2727;
             14'h642 	:	val_out <= 16'h272d;
             14'h643 	:	val_out <= 16'h2733;
             14'h644 	:	val_out <= 16'h2739;
             14'h645 	:	val_out <= 16'h273f;
             14'h646 	:	val_out <= 16'h2746;
             14'h647 	:	val_out <= 16'h274c;
             14'h648 	:	val_out <= 16'h2752;
             14'h649 	:	val_out <= 16'h2758;
             14'h64a 	:	val_out <= 16'h275e;
             14'h64b 	:	val_out <= 16'h2765;
             14'h64c 	:	val_out <= 16'h276b;
             14'h64d 	:	val_out <= 16'h2771;
             14'h64e 	:	val_out <= 16'h2777;
             14'h64f 	:	val_out <= 16'h277d;
             14'h650 	:	val_out <= 16'h2784;
             14'h651 	:	val_out <= 16'h278a;
             14'h652 	:	val_out <= 16'h2790;
             14'h653 	:	val_out <= 16'h2796;
             14'h654 	:	val_out <= 16'h279c;
             14'h655 	:	val_out <= 16'h27a3;
             14'h656 	:	val_out <= 16'h27a9;
             14'h657 	:	val_out <= 16'h27af;
             14'h658 	:	val_out <= 16'h27b5;
             14'h659 	:	val_out <= 16'h27bc;
             14'h65a 	:	val_out <= 16'h27c2;
             14'h65b 	:	val_out <= 16'h27c8;
             14'h65c 	:	val_out <= 16'h27ce;
             14'h65d 	:	val_out <= 16'h27d4;
             14'h65e 	:	val_out <= 16'h27db;
             14'h65f 	:	val_out <= 16'h27e1;
             14'h660 	:	val_out <= 16'h27e7;
             14'h661 	:	val_out <= 16'h27ed;
             14'h662 	:	val_out <= 16'h27f3;
             14'h663 	:	val_out <= 16'h27fa;
             14'h664 	:	val_out <= 16'h2800;
             14'h665 	:	val_out <= 16'h2806;
             14'h666 	:	val_out <= 16'h280c;
             14'h667 	:	val_out <= 16'h2812;
             14'h668 	:	val_out <= 16'h2819;
             14'h669 	:	val_out <= 16'h281f;
             14'h66a 	:	val_out <= 16'h2825;
             14'h66b 	:	val_out <= 16'h282b;
             14'h66c 	:	val_out <= 16'h2831;
             14'h66d 	:	val_out <= 16'h2838;
             14'h66e 	:	val_out <= 16'h283e;
             14'h66f 	:	val_out <= 16'h2844;
             14'h670 	:	val_out <= 16'h284a;
             14'h671 	:	val_out <= 16'h2850;
             14'h672 	:	val_out <= 16'h2857;
             14'h673 	:	val_out <= 16'h285d;
             14'h674 	:	val_out <= 16'h2863;
             14'h675 	:	val_out <= 16'h2869;
             14'h676 	:	val_out <= 16'h286f;
             14'h677 	:	val_out <= 16'h2876;
             14'h678 	:	val_out <= 16'h287c;
             14'h679 	:	val_out <= 16'h2882;
             14'h67a 	:	val_out <= 16'h2888;
             14'h67b 	:	val_out <= 16'h288f;
             14'h67c 	:	val_out <= 16'h2895;
             14'h67d 	:	val_out <= 16'h289b;
             14'h67e 	:	val_out <= 16'h28a1;
             14'h67f 	:	val_out <= 16'h28a7;
             14'h680 	:	val_out <= 16'h28ae;
             14'h681 	:	val_out <= 16'h28b4;
             14'h682 	:	val_out <= 16'h28ba;
             14'h683 	:	val_out <= 16'h28c0;
             14'h684 	:	val_out <= 16'h28c6;
             14'h685 	:	val_out <= 16'h28cd;
             14'h686 	:	val_out <= 16'h28d3;
             14'h687 	:	val_out <= 16'h28d9;
             14'h688 	:	val_out <= 16'h28df;
             14'h689 	:	val_out <= 16'h28e5;
             14'h68a 	:	val_out <= 16'h28ec;
             14'h68b 	:	val_out <= 16'h28f2;
             14'h68c 	:	val_out <= 16'h28f8;
             14'h68d 	:	val_out <= 16'h28fe;
             14'h68e 	:	val_out <= 16'h2904;
             14'h68f 	:	val_out <= 16'h290b;
             14'h690 	:	val_out <= 16'h2911;
             14'h691 	:	val_out <= 16'h2917;
             14'h692 	:	val_out <= 16'h291d;
             14'h693 	:	val_out <= 16'h2923;
             14'h694 	:	val_out <= 16'h292a;
             14'h695 	:	val_out <= 16'h2930;
             14'h696 	:	val_out <= 16'h2936;
             14'h697 	:	val_out <= 16'h293c;
             14'h698 	:	val_out <= 16'h2942;
             14'h699 	:	val_out <= 16'h2949;
             14'h69a 	:	val_out <= 16'h294f;
             14'h69b 	:	val_out <= 16'h2955;
             14'h69c 	:	val_out <= 16'h295b;
             14'h69d 	:	val_out <= 16'h2961;
             14'h69e 	:	val_out <= 16'h2968;
             14'h69f 	:	val_out <= 16'h296e;
             14'h6a0 	:	val_out <= 16'h2974;
             14'h6a1 	:	val_out <= 16'h297a;
             14'h6a2 	:	val_out <= 16'h2980;
             14'h6a3 	:	val_out <= 16'h2987;
             14'h6a4 	:	val_out <= 16'h298d;
             14'h6a5 	:	val_out <= 16'h2993;
             14'h6a6 	:	val_out <= 16'h2999;
             14'h6a7 	:	val_out <= 16'h299f;
             14'h6a8 	:	val_out <= 16'h29a6;
             14'h6a9 	:	val_out <= 16'h29ac;
             14'h6aa 	:	val_out <= 16'h29b2;
             14'h6ab 	:	val_out <= 16'h29b8;
             14'h6ac 	:	val_out <= 16'h29be;
             14'h6ad 	:	val_out <= 16'h29c5;
             14'h6ae 	:	val_out <= 16'h29cb;
             14'h6af 	:	val_out <= 16'h29d1;
             14'h6b0 	:	val_out <= 16'h29d7;
             14'h6b1 	:	val_out <= 16'h29dd;
             14'h6b2 	:	val_out <= 16'h29e4;
             14'h6b3 	:	val_out <= 16'h29ea;
             14'h6b4 	:	val_out <= 16'h29f0;
             14'h6b5 	:	val_out <= 16'h29f6;
             14'h6b6 	:	val_out <= 16'h29fc;
             14'h6b7 	:	val_out <= 16'h2a03;
             14'h6b8 	:	val_out <= 16'h2a09;
             14'h6b9 	:	val_out <= 16'h2a0f;
             14'h6ba 	:	val_out <= 16'h2a15;
             14'h6bb 	:	val_out <= 16'h2a1b;
             14'h6bc 	:	val_out <= 16'h2a22;
             14'h6bd 	:	val_out <= 16'h2a28;
             14'h6be 	:	val_out <= 16'h2a2e;
             14'h6bf 	:	val_out <= 16'h2a34;
             14'h6c0 	:	val_out <= 16'h2a3a;
             14'h6c1 	:	val_out <= 16'h2a41;
             14'h6c2 	:	val_out <= 16'h2a47;
             14'h6c3 	:	val_out <= 16'h2a4d;
             14'h6c4 	:	val_out <= 16'h2a53;
             14'h6c5 	:	val_out <= 16'h2a59;
             14'h6c6 	:	val_out <= 16'h2a60;
             14'h6c7 	:	val_out <= 16'h2a66;
             14'h6c8 	:	val_out <= 16'h2a6c;
             14'h6c9 	:	val_out <= 16'h2a72;
             14'h6ca 	:	val_out <= 16'h2a78;
             14'h6cb 	:	val_out <= 16'h2a7f;
             14'h6cc 	:	val_out <= 16'h2a85;
             14'h6cd 	:	val_out <= 16'h2a8b;
             14'h6ce 	:	val_out <= 16'h2a91;
             14'h6cf 	:	val_out <= 16'h2a97;
             14'h6d0 	:	val_out <= 16'h2a9d;
             14'h6d1 	:	val_out <= 16'h2aa4;
             14'h6d2 	:	val_out <= 16'h2aaa;
             14'h6d3 	:	val_out <= 16'h2ab0;
             14'h6d4 	:	val_out <= 16'h2ab6;
             14'h6d5 	:	val_out <= 16'h2abc;
             14'h6d6 	:	val_out <= 16'h2ac3;
             14'h6d7 	:	val_out <= 16'h2ac9;
             14'h6d8 	:	val_out <= 16'h2acf;
             14'h6d9 	:	val_out <= 16'h2ad5;
             14'h6da 	:	val_out <= 16'h2adb;
             14'h6db 	:	val_out <= 16'h2ae2;
             14'h6dc 	:	val_out <= 16'h2ae8;
             14'h6dd 	:	val_out <= 16'h2aee;
             14'h6de 	:	val_out <= 16'h2af4;
             14'h6df 	:	val_out <= 16'h2afa;
             14'h6e0 	:	val_out <= 16'h2b01;
             14'h6e1 	:	val_out <= 16'h2b07;
             14'h6e2 	:	val_out <= 16'h2b0d;
             14'h6e3 	:	val_out <= 16'h2b13;
             14'h6e4 	:	val_out <= 16'h2b19;
             14'h6e5 	:	val_out <= 16'h2b20;
             14'h6e6 	:	val_out <= 16'h2b26;
             14'h6e7 	:	val_out <= 16'h2b2c;
             14'h6e8 	:	val_out <= 16'h2b32;
             14'h6e9 	:	val_out <= 16'h2b38;
             14'h6ea 	:	val_out <= 16'h2b3f;
             14'h6eb 	:	val_out <= 16'h2b45;
             14'h6ec 	:	val_out <= 16'h2b4b;
             14'h6ed 	:	val_out <= 16'h2b51;
             14'h6ee 	:	val_out <= 16'h2b57;
             14'h6ef 	:	val_out <= 16'h2b5d;
             14'h6f0 	:	val_out <= 16'h2b64;
             14'h6f1 	:	val_out <= 16'h2b6a;
             14'h6f2 	:	val_out <= 16'h2b70;
             14'h6f3 	:	val_out <= 16'h2b76;
             14'h6f4 	:	val_out <= 16'h2b7c;
             14'h6f5 	:	val_out <= 16'h2b83;
             14'h6f6 	:	val_out <= 16'h2b89;
             14'h6f7 	:	val_out <= 16'h2b8f;
             14'h6f8 	:	val_out <= 16'h2b95;
             14'h6f9 	:	val_out <= 16'h2b9b;
             14'h6fa 	:	val_out <= 16'h2ba2;
             14'h6fb 	:	val_out <= 16'h2ba8;
             14'h6fc 	:	val_out <= 16'h2bae;
             14'h6fd 	:	val_out <= 16'h2bb4;
             14'h6fe 	:	val_out <= 16'h2bba;
             14'h6ff 	:	val_out <= 16'h2bc1;
             14'h700 	:	val_out <= 16'h2bc7;
             14'h701 	:	val_out <= 16'h2bcd;
             14'h702 	:	val_out <= 16'h2bd3;
             14'h703 	:	val_out <= 16'h2bd9;
             14'h704 	:	val_out <= 16'h2be0;
             14'h705 	:	val_out <= 16'h2be6;
             14'h706 	:	val_out <= 16'h2bec;
             14'h707 	:	val_out <= 16'h2bf2;
             14'h708 	:	val_out <= 16'h2bf8;
             14'h709 	:	val_out <= 16'h2bfe;
             14'h70a 	:	val_out <= 16'h2c05;
             14'h70b 	:	val_out <= 16'h2c0b;
             14'h70c 	:	val_out <= 16'h2c11;
             14'h70d 	:	val_out <= 16'h2c17;
             14'h70e 	:	val_out <= 16'h2c1d;
             14'h70f 	:	val_out <= 16'h2c24;
             14'h710 	:	val_out <= 16'h2c2a;
             14'h711 	:	val_out <= 16'h2c30;
             14'h712 	:	val_out <= 16'h2c36;
             14'h713 	:	val_out <= 16'h2c3c;
             14'h714 	:	val_out <= 16'h2c43;
             14'h715 	:	val_out <= 16'h2c49;
             14'h716 	:	val_out <= 16'h2c4f;
             14'h717 	:	val_out <= 16'h2c55;
             14'h718 	:	val_out <= 16'h2c5b;
             14'h719 	:	val_out <= 16'h2c61;
             14'h71a 	:	val_out <= 16'h2c68;
             14'h71b 	:	val_out <= 16'h2c6e;
             14'h71c 	:	val_out <= 16'h2c74;
             14'h71d 	:	val_out <= 16'h2c7a;
             14'h71e 	:	val_out <= 16'h2c80;
             14'h71f 	:	val_out <= 16'h2c87;
             14'h720 	:	val_out <= 16'h2c8d;
             14'h721 	:	val_out <= 16'h2c93;
             14'h722 	:	val_out <= 16'h2c99;
             14'h723 	:	val_out <= 16'h2c9f;
             14'h724 	:	val_out <= 16'h2ca6;
             14'h725 	:	val_out <= 16'h2cac;
             14'h726 	:	val_out <= 16'h2cb2;
             14'h727 	:	val_out <= 16'h2cb8;
             14'h728 	:	val_out <= 16'h2cbe;
             14'h729 	:	val_out <= 16'h2cc4;
             14'h72a 	:	val_out <= 16'h2ccb;
             14'h72b 	:	val_out <= 16'h2cd1;
             14'h72c 	:	val_out <= 16'h2cd7;
             14'h72d 	:	val_out <= 16'h2cdd;
             14'h72e 	:	val_out <= 16'h2ce3;
             14'h72f 	:	val_out <= 16'h2cea;
             14'h730 	:	val_out <= 16'h2cf0;
             14'h731 	:	val_out <= 16'h2cf6;
             14'h732 	:	val_out <= 16'h2cfc;
             14'h733 	:	val_out <= 16'h2d02;
             14'h734 	:	val_out <= 16'h2d09;
             14'h735 	:	val_out <= 16'h2d0f;
             14'h736 	:	val_out <= 16'h2d15;
             14'h737 	:	val_out <= 16'h2d1b;
             14'h738 	:	val_out <= 16'h2d21;
             14'h739 	:	val_out <= 16'h2d27;
             14'h73a 	:	val_out <= 16'h2d2e;
             14'h73b 	:	val_out <= 16'h2d34;
             14'h73c 	:	val_out <= 16'h2d3a;
             14'h73d 	:	val_out <= 16'h2d40;
             14'h73e 	:	val_out <= 16'h2d46;
             14'h73f 	:	val_out <= 16'h2d4d;
             14'h740 	:	val_out <= 16'h2d53;
             14'h741 	:	val_out <= 16'h2d59;
             14'h742 	:	val_out <= 16'h2d5f;
             14'h743 	:	val_out <= 16'h2d65;
             14'h744 	:	val_out <= 16'h2d6b;
             14'h745 	:	val_out <= 16'h2d72;
             14'h746 	:	val_out <= 16'h2d78;
             14'h747 	:	val_out <= 16'h2d7e;
             14'h748 	:	val_out <= 16'h2d84;
             14'h749 	:	val_out <= 16'h2d8a;
             14'h74a 	:	val_out <= 16'h2d91;
             14'h74b 	:	val_out <= 16'h2d97;
             14'h74c 	:	val_out <= 16'h2d9d;
             14'h74d 	:	val_out <= 16'h2da3;
             14'h74e 	:	val_out <= 16'h2da9;
             14'h74f 	:	val_out <= 16'h2daf;
             14'h750 	:	val_out <= 16'h2db6;
             14'h751 	:	val_out <= 16'h2dbc;
             14'h752 	:	val_out <= 16'h2dc2;
             14'h753 	:	val_out <= 16'h2dc8;
             14'h754 	:	val_out <= 16'h2dce;
             14'h755 	:	val_out <= 16'h2dd5;
             14'h756 	:	val_out <= 16'h2ddb;
             14'h757 	:	val_out <= 16'h2de1;
             14'h758 	:	val_out <= 16'h2de7;
             14'h759 	:	val_out <= 16'h2ded;
             14'h75a 	:	val_out <= 16'h2df3;
             14'h75b 	:	val_out <= 16'h2dfa;
             14'h75c 	:	val_out <= 16'h2e00;
             14'h75d 	:	val_out <= 16'h2e06;
             14'h75e 	:	val_out <= 16'h2e0c;
             14'h75f 	:	val_out <= 16'h2e12;
             14'h760 	:	val_out <= 16'h2e19;
             14'h761 	:	val_out <= 16'h2e1f;
             14'h762 	:	val_out <= 16'h2e25;
             14'h763 	:	val_out <= 16'h2e2b;
             14'h764 	:	val_out <= 16'h2e31;
             14'h765 	:	val_out <= 16'h2e37;
             14'h766 	:	val_out <= 16'h2e3e;
             14'h767 	:	val_out <= 16'h2e44;
             14'h768 	:	val_out <= 16'h2e4a;
             14'h769 	:	val_out <= 16'h2e50;
             14'h76a 	:	val_out <= 16'h2e56;
             14'h76b 	:	val_out <= 16'h2e5d;
             14'h76c 	:	val_out <= 16'h2e63;
             14'h76d 	:	val_out <= 16'h2e69;
             14'h76e 	:	val_out <= 16'h2e6f;
             14'h76f 	:	val_out <= 16'h2e75;
             14'h770 	:	val_out <= 16'h2e7b;
             14'h771 	:	val_out <= 16'h2e82;
             14'h772 	:	val_out <= 16'h2e88;
             14'h773 	:	val_out <= 16'h2e8e;
             14'h774 	:	val_out <= 16'h2e94;
             14'h775 	:	val_out <= 16'h2e9a;
             14'h776 	:	val_out <= 16'h2ea1;
             14'h777 	:	val_out <= 16'h2ea7;
             14'h778 	:	val_out <= 16'h2ead;
             14'h779 	:	val_out <= 16'h2eb3;
             14'h77a 	:	val_out <= 16'h2eb9;
             14'h77b 	:	val_out <= 16'h2ebf;
             14'h77c 	:	val_out <= 16'h2ec6;
             14'h77d 	:	val_out <= 16'h2ecc;
             14'h77e 	:	val_out <= 16'h2ed2;
             14'h77f 	:	val_out <= 16'h2ed8;
             14'h780 	:	val_out <= 16'h2ede;
             14'h781 	:	val_out <= 16'h2ee4;
             14'h782 	:	val_out <= 16'h2eeb;
             14'h783 	:	val_out <= 16'h2ef1;
             14'h784 	:	val_out <= 16'h2ef7;
             14'h785 	:	val_out <= 16'h2efd;
             14'h786 	:	val_out <= 16'h2f03;
             14'h787 	:	val_out <= 16'h2f0a;
             14'h788 	:	val_out <= 16'h2f10;
             14'h789 	:	val_out <= 16'h2f16;
             14'h78a 	:	val_out <= 16'h2f1c;
             14'h78b 	:	val_out <= 16'h2f22;
             14'h78c 	:	val_out <= 16'h2f28;
             14'h78d 	:	val_out <= 16'h2f2f;
             14'h78e 	:	val_out <= 16'h2f35;
             14'h78f 	:	val_out <= 16'h2f3b;
             14'h790 	:	val_out <= 16'h2f41;
             14'h791 	:	val_out <= 16'h2f47;
             14'h792 	:	val_out <= 16'h2f4d;
             14'h793 	:	val_out <= 16'h2f54;
             14'h794 	:	val_out <= 16'h2f5a;
             14'h795 	:	val_out <= 16'h2f60;
             14'h796 	:	val_out <= 16'h2f66;
             14'h797 	:	val_out <= 16'h2f6c;
             14'h798 	:	val_out <= 16'h2f73;
             14'h799 	:	val_out <= 16'h2f79;
             14'h79a 	:	val_out <= 16'h2f7f;
             14'h79b 	:	val_out <= 16'h2f85;
             14'h79c 	:	val_out <= 16'h2f8b;
             14'h79d 	:	val_out <= 16'h2f91;
             14'h79e 	:	val_out <= 16'h2f98;
             14'h79f 	:	val_out <= 16'h2f9e;
             14'h7a0 	:	val_out <= 16'h2fa4;
             14'h7a1 	:	val_out <= 16'h2faa;
             14'h7a2 	:	val_out <= 16'h2fb0;
             14'h7a3 	:	val_out <= 16'h2fb6;
             14'h7a4 	:	val_out <= 16'h2fbd;
             14'h7a5 	:	val_out <= 16'h2fc3;
             14'h7a6 	:	val_out <= 16'h2fc9;
             14'h7a7 	:	val_out <= 16'h2fcf;
             14'h7a8 	:	val_out <= 16'h2fd5;
             14'h7a9 	:	val_out <= 16'h2fdb;
             14'h7aa 	:	val_out <= 16'h2fe2;
             14'h7ab 	:	val_out <= 16'h2fe8;
             14'h7ac 	:	val_out <= 16'h2fee;
             14'h7ad 	:	val_out <= 16'h2ff4;
             14'h7ae 	:	val_out <= 16'h2ffa;
             14'h7af 	:	val_out <= 16'h3000;
             14'h7b0 	:	val_out <= 16'h3007;
             14'h7b1 	:	val_out <= 16'h300d;
             14'h7b2 	:	val_out <= 16'h3013;
             14'h7b3 	:	val_out <= 16'h3019;
             14'h7b4 	:	val_out <= 16'h301f;
             14'h7b5 	:	val_out <= 16'h3026;
             14'h7b6 	:	val_out <= 16'h302c;
             14'h7b7 	:	val_out <= 16'h3032;
             14'h7b8 	:	val_out <= 16'h3038;
             14'h7b9 	:	val_out <= 16'h303e;
             14'h7ba 	:	val_out <= 16'h3044;
             14'h7bb 	:	val_out <= 16'h304b;
             14'h7bc 	:	val_out <= 16'h3051;
             14'h7bd 	:	val_out <= 16'h3057;
             14'h7be 	:	val_out <= 16'h305d;
             14'h7bf 	:	val_out <= 16'h3063;
             14'h7c0 	:	val_out <= 16'h3069;
             14'h7c1 	:	val_out <= 16'h3070;
             14'h7c2 	:	val_out <= 16'h3076;
             14'h7c3 	:	val_out <= 16'h307c;
             14'h7c4 	:	val_out <= 16'h3082;
             14'h7c5 	:	val_out <= 16'h3088;
             14'h7c6 	:	val_out <= 16'h308e;
             14'h7c7 	:	val_out <= 16'h3095;
             14'h7c8 	:	val_out <= 16'h309b;
             14'h7c9 	:	val_out <= 16'h30a1;
             14'h7ca 	:	val_out <= 16'h30a7;
             14'h7cb 	:	val_out <= 16'h30ad;
             14'h7cc 	:	val_out <= 16'h30b3;
             14'h7cd 	:	val_out <= 16'h30ba;
             14'h7ce 	:	val_out <= 16'h30c0;
             14'h7cf 	:	val_out <= 16'h30c6;
             14'h7d0 	:	val_out <= 16'h30cc;
             14'h7d1 	:	val_out <= 16'h30d2;
             14'h7d2 	:	val_out <= 16'h30d8;
             14'h7d3 	:	val_out <= 16'h30df;
             14'h7d4 	:	val_out <= 16'h30e5;
             14'h7d5 	:	val_out <= 16'h30eb;
             14'h7d6 	:	val_out <= 16'h30f1;
             14'h7d7 	:	val_out <= 16'h30f7;
             14'h7d8 	:	val_out <= 16'h30fd;
             14'h7d9 	:	val_out <= 16'h3104;
             14'h7da 	:	val_out <= 16'h310a;
             14'h7db 	:	val_out <= 16'h3110;
             14'h7dc 	:	val_out <= 16'h3116;
             14'h7dd 	:	val_out <= 16'h311c;
             14'h7de 	:	val_out <= 16'h3122;
             14'h7df 	:	val_out <= 16'h3129;
             14'h7e0 	:	val_out <= 16'h312f;
             14'h7e1 	:	val_out <= 16'h3135;
             14'h7e2 	:	val_out <= 16'h313b;
             14'h7e3 	:	val_out <= 16'h3141;
             14'h7e4 	:	val_out <= 16'h3147;
             14'h7e5 	:	val_out <= 16'h314e;
             14'h7e6 	:	val_out <= 16'h3154;
             14'h7e7 	:	val_out <= 16'h315a;
             14'h7e8 	:	val_out <= 16'h3160;
             14'h7e9 	:	val_out <= 16'h3166;
             14'h7ea 	:	val_out <= 16'h316c;
             14'h7eb 	:	val_out <= 16'h3173;
             14'h7ec 	:	val_out <= 16'h3179;
             14'h7ed 	:	val_out <= 16'h317f;
             14'h7ee 	:	val_out <= 16'h3185;
             14'h7ef 	:	val_out <= 16'h318b;
             14'h7f0 	:	val_out <= 16'h3191;
             14'h7f1 	:	val_out <= 16'h3198;
             14'h7f2 	:	val_out <= 16'h319e;
             14'h7f3 	:	val_out <= 16'h31a4;
             14'h7f4 	:	val_out <= 16'h31aa;
             14'h7f5 	:	val_out <= 16'h31b0;
             14'h7f6 	:	val_out <= 16'h31b6;
             14'h7f7 	:	val_out <= 16'h31bd;
             14'h7f8 	:	val_out <= 16'h31c3;
             14'h7f9 	:	val_out <= 16'h31c9;
             14'h7fa 	:	val_out <= 16'h31cf;
             14'h7fb 	:	val_out <= 16'h31d5;
             14'h7fc 	:	val_out <= 16'h31db;
             14'h7fd 	:	val_out <= 16'h31e2;
             14'h7fe 	:	val_out <= 16'h31e8;
             14'h7ff 	:	val_out <= 16'h31ee;
             14'h800 	:	val_out <= 16'h31f4;
             14'h801 	:	val_out <= 16'h31fa;
             14'h802 	:	val_out <= 16'h3200;
             14'h803 	:	val_out <= 16'h3207;
             14'h804 	:	val_out <= 16'h320d;
             14'h805 	:	val_out <= 16'h3213;
             14'h806 	:	val_out <= 16'h3219;
             14'h807 	:	val_out <= 16'h321f;
             14'h808 	:	val_out <= 16'h3225;
             14'h809 	:	val_out <= 16'h322b;
             14'h80a 	:	val_out <= 16'h3232;
             14'h80b 	:	val_out <= 16'h3238;
             14'h80c 	:	val_out <= 16'h323e;
             14'h80d 	:	val_out <= 16'h3244;
             14'h80e 	:	val_out <= 16'h324a;
             14'h80f 	:	val_out <= 16'h3250;
             14'h810 	:	val_out <= 16'h3257;
             14'h811 	:	val_out <= 16'h325d;
             14'h812 	:	val_out <= 16'h3263;
             14'h813 	:	val_out <= 16'h3269;
             14'h814 	:	val_out <= 16'h326f;
             14'h815 	:	val_out <= 16'h3275;
             14'h816 	:	val_out <= 16'h327c;
             14'h817 	:	val_out <= 16'h3282;
             14'h818 	:	val_out <= 16'h3288;
             14'h819 	:	val_out <= 16'h328e;
             14'h81a 	:	val_out <= 16'h3294;
             14'h81b 	:	val_out <= 16'h329a;
             14'h81c 	:	val_out <= 16'h32a1;
             14'h81d 	:	val_out <= 16'h32a7;
             14'h81e 	:	val_out <= 16'h32ad;
             14'h81f 	:	val_out <= 16'h32b3;
             14'h820 	:	val_out <= 16'h32b9;
             14'h821 	:	val_out <= 16'h32bf;
             14'h822 	:	val_out <= 16'h32c5;
             14'h823 	:	val_out <= 16'h32cc;
             14'h824 	:	val_out <= 16'h32d2;
             14'h825 	:	val_out <= 16'h32d8;
             14'h826 	:	val_out <= 16'h32de;
             14'h827 	:	val_out <= 16'h32e4;
             14'h828 	:	val_out <= 16'h32ea;
             14'h829 	:	val_out <= 16'h32f1;
             14'h82a 	:	val_out <= 16'h32f7;
             14'h82b 	:	val_out <= 16'h32fd;
             14'h82c 	:	val_out <= 16'h3303;
             14'h82d 	:	val_out <= 16'h3309;
             14'h82e 	:	val_out <= 16'h330f;
             14'h82f 	:	val_out <= 16'h3316;
             14'h830 	:	val_out <= 16'h331c;
             14'h831 	:	val_out <= 16'h3322;
             14'h832 	:	val_out <= 16'h3328;
             14'h833 	:	val_out <= 16'h332e;
             14'h834 	:	val_out <= 16'h3334;
             14'h835 	:	val_out <= 16'h333a;
             14'h836 	:	val_out <= 16'h3341;
             14'h837 	:	val_out <= 16'h3347;
             14'h838 	:	val_out <= 16'h334d;
             14'h839 	:	val_out <= 16'h3353;
             14'h83a 	:	val_out <= 16'h3359;
             14'h83b 	:	val_out <= 16'h335f;
             14'h83c 	:	val_out <= 16'h3366;
             14'h83d 	:	val_out <= 16'h336c;
             14'h83e 	:	val_out <= 16'h3372;
             14'h83f 	:	val_out <= 16'h3378;
             14'h840 	:	val_out <= 16'h337e;
             14'h841 	:	val_out <= 16'h3384;
             14'h842 	:	val_out <= 16'h338a;
             14'h843 	:	val_out <= 16'h3391;
             14'h844 	:	val_out <= 16'h3397;
             14'h845 	:	val_out <= 16'h339d;
             14'h846 	:	val_out <= 16'h33a3;
             14'h847 	:	val_out <= 16'h33a9;
             14'h848 	:	val_out <= 16'h33af;
             14'h849 	:	val_out <= 16'h33b6;
             14'h84a 	:	val_out <= 16'h33bc;
             14'h84b 	:	val_out <= 16'h33c2;
             14'h84c 	:	val_out <= 16'h33c8;
             14'h84d 	:	val_out <= 16'h33ce;
             14'h84e 	:	val_out <= 16'h33d4;
             14'h84f 	:	val_out <= 16'h33da;
             14'h850 	:	val_out <= 16'h33e1;
             14'h851 	:	val_out <= 16'h33e7;
             14'h852 	:	val_out <= 16'h33ed;
             14'h853 	:	val_out <= 16'h33f3;
             14'h854 	:	val_out <= 16'h33f9;
             14'h855 	:	val_out <= 16'h33ff;
             14'h856 	:	val_out <= 16'h3406;
             14'h857 	:	val_out <= 16'h340c;
             14'h858 	:	val_out <= 16'h3412;
             14'h859 	:	val_out <= 16'h3418;
             14'h85a 	:	val_out <= 16'h341e;
             14'h85b 	:	val_out <= 16'h3424;
             14'h85c 	:	val_out <= 16'h342a;
             14'h85d 	:	val_out <= 16'h3431;
             14'h85e 	:	val_out <= 16'h3437;
             14'h85f 	:	val_out <= 16'h343d;
             14'h860 	:	val_out <= 16'h3443;
             14'h861 	:	val_out <= 16'h3449;
             14'h862 	:	val_out <= 16'h344f;
             14'h863 	:	val_out <= 16'h3456;
             14'h864 	:	val_out <= 16'h345c;
             14'h865 	:	val_out <= 16'h3462;
             14'h866 	:	val_out <= 16'h3468;
             14'h867 	:	val_out <= 16'h346e;
             14'h868 	:	val_out <= 16'h3474;
             14'h869 	:	val_out <= 16'h347a;
             14'h86a 	:	val_out <= 16'h3481;
             14'h86b 	:	val_out <= 16'h3487;
             14'h86c 	:	val_out <= 16'h348d;
             14'h86d 	:	val_out <= 16'h3493;
             14'h86e 	:	val_out <= 16'h3499;
             14'h86f 	:	val_out <= 16'h349f;
             14'h870 	:	val_out <= 16'h34a5;
             14'h871 	:	val_out <= 16'h34ac;
             14'h872 	:	val_out <= 16'h34b2;
             14'h873 	:	val_out <= 16'h34b8;
             14'h874 	:	val_out <= 16'h34be;
             14'h875 	:	val_out <= 16'h34c4;
             14'h876 	:	val_out <= 16'h34ca;
             14'h877 	:	val_out <= 16'h34d0;
             14'h878 	:	val_out <= 16'h34d7;
             14'h879 	:	val_out <= 16'h34dd;
             14'h87a 	:	val_out <= 16'h34e3;
             14'h87b 	:	val_out <= 16'h34e9;
             14'h87c 	:	val_out <= 16'h34ef;
             14'h87d 	:	val_out <= 16'h34f5;
             14'h87e 	:	val_out <= 16'h34fc;
             14'h87f 	:	val_out <= 16'h3502;
             14'h880 	:	val_out <= 16'h3508;
             14'h881 	:	val_out <= 16'h350e;
             14'h882 	:	val_out <= 16'h3514;
             14'h883 	:	val_out <= 16'h351a;
             14'h884 	:	val_out <= 16'h3520;
             14'h885 	:	val_out <= 16'h3527;
             14'h886 	:	val_out <= 16'h352d;
             14'h887 	:	val_out <= 16'h3533;
             14'h888 	:	val_out <= 16'h3539;
             14'h889 	:	val_out <= 16'h353f;
             14'h88a 	:	val_out <= 16'h3545;
             14'h88b 	:	val_out <= 16'h354b;
             14'h88c 	:	val_out <= 16'h3552;
             14'h88d 	:	val_out <= 16'h3558;
             14'h88e 	:	val_out <= 16'h355e;
             14'h88f 	:	val_out <= 16'h3564;
             14'h890 	:	val_out <= 16'h356a;
             14'h891 	:	val_out <= 16'h3570;
             14'h892 	:	val_out <= 16'h3576;
             14'h893 	:	val_out <= 16'h357d;
             14'h894 	:	val_out <= 16'h3583;
             14'h895 	:	val_out <= 16'h3589;
             14'h896 	:	val_out <= 16'h358f;
             14'h897 	:	val_out <= 16'h3595;
             14'h898 	:	val_out <= 16'h359b;
             14'h899 	:	val_out <= 16'h35a1;
             14'h89a 	:	val_out <= 16'h35a8;
             14'h89b 	:	val_out <= 16'h35ae;
             14'h89c 	:	val_out <= 16'h35b4;
             14'h89d 	:	val_out <= 16'h35ba;
             14'h89e 	:	val_out <= 16'h35c0;
             14'h89f 	:	val_out <= 16'h35c6;
             14'h8a0 	:	val_out <= 16'h35cc;
             14'h8a1 	:	val_out <= 16'h35d3;
             14'h8a2 	:	val_out <= 16'h35d9;
             14'h8a3 	:	val_out <= 16'h35df;
             14'h8a4 	:	val_out <= 16'h35e5;
             14'h8a5 	:	val_out <= 16'h35eb;
             14'h8a6 	:	val_out <= 16'h35f1;
             14'h8a7 	:	val_out <= 16'h35f7;
             14'h8a8 	:	val_out <= 16'h35fe;
             14'h8a9 	:	val_out <= 16'h3604;
             14'h8aa 	:	val_out <= 16'h360a;
             14'h8ab 	:	val_out <= 16'h3610;
             14'h8ac 	:	val_out <= 16'h3616;
             14'h8ad 	:	val_out <= 16'h361c;
             14'h8ae 	:	val_out <= 16'h3622;
             14'h8af 	:	val_out <= 16'h3629;
             14'h8b0 	:	val_out <= 16'h362f;
             14'h8b1 	:	val_out <= 16'h3635;
             14'h8b2 	:	val_out <= 16'h363b;
             14'h8b3 	:	val_out <= 16'h3641;
             14'h8b4 	:	val_out <= 16'h3647;
             14'h8b5 	:	val_out <= 16'h364d;
             14'h8b6 	:	val_out <= 16'h3654;
             14'h8b7 	:	val_out <= 16'h365a;
             14'h8b8 	:	val_out <= 16'h3660;
             14'h8b9 	:	val_out <= 16'h3666;
             14'h8ba 	:	val_out <= 16'h366c;
             14'h8bb 	:	val_out <= 16'h3672;
             14'h8bc 	:	val_out <= 16'h3678;
             14'h8bd 	:	val_out <= 16'h367f;
             14'h8be 	:	val_out <= 16'h3685;
             14'h8bf 	:	val_out <= 16'h368b;
             14'h8c0 	:	val_out <= 16'h3691;
             14'h8c1 	:	val_out <= 16'h3697;
             14'h8c2 	:	val_out <= 16'h369d;
             14'h8c3 	:	val_out <= 16'h36a3;
             14'h8c4 	:	val_out <= 16'h36aa;
             14'h8c5 	:	val_out <= 16'h36b0;
             14'h8c6 	:	val_out <= 16'h36b6;
             14'h8c7 	:	val_out <= 16'h36bc;
             14'h8c8 	:	val_out <= 16'h36c2;
             14'h8c9 	:	val_out <= 16'h36c8;
             14'h8ca 	:	val_out <= 16'h36ce;
             14'h8cb 	:	val_out <= 16'h36d4;
             14'h8cc 	:	val_out <= 16'h36db;
             14'h8cd 	:	val_out <= 16'h36e1;
             14'h8ce 	:	val_out <= 16'h36e7;
             14'h8cf 	:	val_out <= 16'h36ed;
             14'h8d0 	:	val_out <= 16'h36f3;
             14'h8d1 	:	val_out <= 16'h36f9;
             14'h8d2 	:	val_out <= 16'h36ff;
             14'h8d3 	:	val_out <= 16'h3706;
             14'h8d4 	:	val_out <= 16'h370c;
             14'h8d5 	:	val_out <= 16'h3712;
             14'h8d6 	:	val_out <= 16'h3718;
             14'h8d7 	:	val_out <= 16'h371e;
             14'h8d8 	:	val_out <= 16'h3724;
             14'h8d9 	:	val_out <= 16'h372a;
             14'h8da 	:	val_out <= 16'h3731;
             14'h8db 	:	val_out <= 16'h3737;
             14'h8dc 	:	val_out <= 16'h373d;
             14'h8dd 	:	val_out <= 16'h3743;
             14'h8de 	:	val_out <= 16'h3749;
             14'h8df 	:	val_out <= 16'h374f;
             14'h8e0 	:	val_out <= 16'h3755;
             14'h8e1 	:	val_out <= 16'h375b;
             14'h8e2 	:	val_out <= 16'h3762;
             14'h8e3 	:	val_out <= 16'h3768;
             14'h8e4 	:	val_out <= 16'h376e;
             14'h8e5 	:	val_out <= 16'h3774;
             14'h8e6 	:	val_out <= 16'h377a;
             14'h8e7 	:	val_out <= 16'h3780;
             14'h8e8 	:	val_out <= 16'h3786;
             14'h8e9 	:	val_out <= 16'h378d;
             14'h8ea 	:	val_out <= 16'h3793;
             14'h8eb 	:	val_out <= 16'h3799;
             14'h8ec 	:	val_out <= 16'h379f;
             14'h8ed 	:	val_out <= 16'h37a5;
             14'h8ee 	:	val_out <= 16'h37ab;
             14'h8ef 	:	val_out <= 16'h37b1;
             14'h8f0 	:	val_out <= 16'h37b7;
             14'h8f1 	:	val_out <= 16'h37be;
             14'h8f2 	:	val_out <= 16'h37c4;
             14'h8f3 	:	val_out <= 16'h37ca;
             14'h8f4 	:	val_out <= 16'h37d0;
             14'h8f5 	:	val_out <= 16'h37d6;
             14'h8f6 	:	val_out <= 16'h37dc;
             14'h8f7 	:	val_out <= 16'h37e2;
             14'h8f8 	:	val_out <= 16'h37e9;
             14'h8f9 	:	val_out <= 16'h37ef;
             14'h8fa 	:	val_out <= 16'h37f5;
             14'h8fb 	:	val_out <= 16'h37fb;
             14'h8fc 	:	val_out <= 16'h3801;
             14'h8fd 	:	val_out <= 16'h3807;
             14'h8fe 	:	val_out <= 16'h380d;
             14'h8ff 	:	val_out <= 16'h3813;
             14'h900 	:	val_out <= 16'h381a;
             14'h901 	:	val_out <= 16'h3820;
             14'h902 	:	val_out <= 16'h3826;
             14'h903 	:	val_out <= 16'h382c;
             14'h904 	:	val_out <= 16'h3832;
             14'h905 	:	val_out <= 16'h3838;
             14'h906 	:	val_out <= 16'h383e;
             14'h907 	:	val_out <= 16'h3844;
             14'h908 	:	val_out <= 16'h384b;
             14'h909 	:	val_out <= 16'h3851;
             14'h90a 	:	val_out <= 16'h3857;
             14'h90b 	:	val_out <= 16'h385d;
             14'h90c 	:	val_out <= 16'h3863;
             14'h90d 	:	val_out <= 16'h3869;
             14'h90e 	:	val_out <= 16'h386f;
             14'h90f 	:	val_out <= 16'h3876;
             14'h910 	:	val_out <= 16'h387c;
             14'h911 	:	val_out <= 16'h3882;
             14'h912 	:	val_out <= 16'h3888;
             14'h913 	:	val_out <= 16'h388e;
             14'h914 	:	val_out <= 16'h3894;
             14'h915 	:	val_out <= 16'h389a;
             14'h916 	:	val_out <= 16'h38a0;
             14'h917 	:	val_out <= 16'h38a7;
             14'h918 	:	val_out <= 16'h38ad;
             14'h919 	:	val_out <= 16'h38b3;
             14'h91a 	:	val_out <= 16'h38b9;
             14'h91b 	:	val_out <= 16'h38bf;
             14'h91c 	:	val_out <= 16'h38c5;
             14'h91d 	:	val_out <= 16'h38cb;
             14'h91e 	:	val_out <= 16'h38d1;
             14'h91f 	:	val_out <= 16'h38d8;
             14'h920 	:	val_out <= 16'h38de;
             14'h921 	:	val_out <= 16'h38e4;
             14'h922 	:	val_out <= 16'h38ea;
             14'h923 	:	val_out <= 16'h38f0;
             14'h924 	:	val_out <= 16'h38f6;
             14'h925 	:	val_out <= 16'h38fc;
             14'h926 	:	val_out <= 16'h3902;
             14'h927 	:	val_out <= 16'h3909;
             14'h928 	:	val_out <= 16'h390f;
             14'h929 	:	val_out <= 16'h3915;
             14'h92a 	:	val_out <= 16'h391b;
             14'h92b 	:	val_out <= 16'h3921;
             14'h92c 	:	val_out <= 16'h3927;
             14'h92d 	:	val_out <= 16'h392d;
             14'h92e 	:	val_out <= 16'h3933;
             14'h92f 	:	val_out <= 16'h393a;
             14'h930 	:	val_out <= 16'h3940;
             14'h931 	:	val_out <= 16'h3946;
             14'h932 	:	val_out <= 16'h394c;
             14'h933 	:	val_out <= 16'h3952;
             14'h934 	:	val_out <= 16'h3958;
             14'h935 	:	val_out <= 16'h395e;
             14'h936 	:	val_out <= 16'h3964;
             14'h937 	:	val_out <= 16'h396b;
             14'h938 	:	val_out <= 16'h3971;
             14'h939 	:	val_out <= 16'h3977;
             14'h93a 	:	val_out <= 16'h397d;
             14'h93b 	:	val_out <= 16'h3983;
             14'h93c 	:	val_out <= 16'h3989;
             14'h93d 	:	val_out <= 16'h398f;
             14'h93e 	:	val_out <= 16'h3995;
             14'h93f 	:	val_out <= 16'h399c;
             14'h940 	:	val_out <= 16'h39a2;
             14'h941 	:	val_out <= 16'h39a8;
             14'h942 	:	val_out <= 16'h39ae;
             14'h943 	:	val_out <= 16'h39b4;
             14'h944 	:	val_out <= 16'h39ba;
             14'h945 	:	val_out <= 16'h39c0;
             14'h946 	:	val_out <= 16'h39c6;
             14'h947 	:	val_out <= 16'h39cd;
             14'h948 	:	val_out <= 16'h39d3;
             14'h949 	:	val_out <= 16'h39d9;
             14'h94a 	:	val_out <= 16'h39df;
             14'h94b 	:	val_out <= 16'h39e5;
             14'h94c 	:	val_out <= 16'h39eb;
             14'h94d 	:	val_out <= 16'h39f1;
             14'h94e 	:	val_out <= 16'h39f7;
             14'h94f 	:	val_out <= 16'h39fd;
             14'h950 	:	val_out <= 16'h3a04;
             14'h951 	:	val_out <= 16'h3a0a;
             14'h952 	:	val_out <= 16'h3a10;
             14'h953 	:	val_out <= 16'h3a16;
             14'h954 	:	val_out <= 16'h3a1c;
             14'h955 	:	val_out <= 16'h3a22;
             14'h956 	:	val_out <= 16'h3a28;
             14'h957 	:	val_out <= 16'h3a2e;
             14'h958 	:	val_out <= 16'h3a35;
             14'h959 	:	val_out <= 16'h3a3b;
             14'h95a 	:	val_out <= 16'h3a41;
             14'h95b 	:	val_out <= 16'h3a47;
             14'h95c 	:	val_out <= 16'h3a4d;
             14'h95d 	:	val_out <= 16'h3a53;
             14'h95e 	:	val_out <= 16'h3a59;
             14'h95f 	:	val_out <= 16'h3a5f;
             14'h960 	:	val_out <= 16'h3a65;
             14'h961 	:	val_out <= 16'h3a6c;
             14'h962 	:	val_out <= 16'h3a72;
             14'h963 	:	val_out <= 16'h3a78;
             14'h964 	:	val_out <= 16'h3a7e;
             14'h965 	:	val_out <= 16'h3a84;
             14'h966 	:	val_out <= 16'h3a8a;
             14'h967 	:	val_out <= 16'h3a90;
             14'h968 	:	val_out <= 16'h3a96;
             14'h969 	:	val_out <= 16'h3a9d;
             14'h96a 	:	val_out <= 16'h3aa3;
             14'h96b 	:	val_out <= 16'h3aa9;
             14'h96c 	:	val_out <= 16'h3aaf;
             14'h96d 	:	val_out <= 16'h3ab5;
             14'h96e 	:	val_out <= 16'h3abb;
             14'h96f 	:	val_out <= 16'h3ac1;
             14'h970 	:	val_out <= 16'h3ac7;
             14'h971 	:	val_out <= 16'h3acd;
             14'h972 	:	val_out <= 16'h3ad4;
             14'h973 	:	val_out <= 16'h3ada;
             14'h974 	:	val_out <= 16'h3ae0;
             14'h975 	:	val_out <= 16'h3ae6;
             14'h976 	:	val_out <= 16'h3aec;
             14'h977 	:	val_out <= 16'h3af2;
             14'h978 	:	val_out <= 16'h3af8;
             14'h979 	:	val_out <= 16'h3afe;
             14'h97a 	:	val_out <= 16'h3b04;
             14'h97b 	:	val_out <= 16'h3b0b;
             14'h97c 	:	val_out <= 16'h3b11;
             14'h97d 	:	val_out <= 16'h3b17;
             14'h97e 	:	val_out <= 16'h3b1d;
             14'h97f 	:	val_out <= 16'h3b23;
             14'h980 	:	val_out <= 16'h3b29;
             14'h981 	:	val_out <= 16'h3b2f;
             14'h982 	:	val_out <= 16'h3b35;
             14'h983 	:	val_out <= 16'h3b3c;
             14'h984 	:	val_out <= 16'h3b42;
             14'h985 	:	val_out <= 16'h3b48;
             14'h986 	:	val_out <= 16'h3b4e;
             14'h987 	:	val_out <= 16'h3b54;
             14'h988 	:	val_out <= 16'h3b5a;
             14'h989 	:	val_out <= 16'h3b60;
             14'h98a 	:	val_out <= 16'h3b66;
             14'h98b 	:	val_out <= 16'h3b6c;
             14'h98c 	:	val_out <= 16'h3b73;
             14'h98d 	:	val_out <= 16'h3b79;
             14'h98e 	:	val_out <= 16'h3b7f;
             14'h98f 	:	val_out <= 16'h3b85;
             14'h990 	:	val_out <= 16'h3b8b;
             14'h991 	:	val_out <= 16'h3b91;
             14'h992 	:	val_out <= 16'h3b97;
             14'h993 	:	val_out <= 16'h3b9d;
             14'h994 	:	val_out <= 16'h3ba3;
             14'h995 	:	val_out <= 16'h3baa;
             14'h996 	:	val_out <= 16'h3bb0;
             14'h997 	:	val_out <= 16'h3bb6;
             14'h998 	:	val_out <= 16'h3bbc;
             14'h999 	:	val_out <= 16'h3bc2;
             14'h99a 	:	val_out <= 16'h3bc8;
             14'h99b 	:	val_out <= 16'h3bce;
             14'h99c 	:	val_out <= 16'h3bd4;
             14'h99d 	:	val_out <= 16'h3bda;
             14'h99e 	:	val_out <= 16'h3be1;
             14'h99f 	:	val_out <= 16'h3be7;
             14'h9a0 	:	val_out <= 16'h3bed;
             14'h9a1 	:	val_out <= 16'h3bf3;
             14'h9a2 	:	val_out <= 16'h3bf9;
             14'h9a3 	:	val_out <= 16'h3bff;
             14'h9a4 	:	val_out <= 16'h3c05;
             14'h9a5 	:	val_out <= 16'h3c0b;
             14'h9a6 	:	val_out <= 16'h3c11;
             14'h9a7 	:	val_out <= 16'h3c17;
             14'h9a8 	:	val_out <= 16'h3c1e;
             14'h9a9 	:	val_out <= 16'h3c24;
             14'h9aa 	:	val_out <= 16'h3c2a;
             14'h9ab 	:	val_out <= 16'h3c30;
             14'h9ac 	:	val_out <= 16'h3c36;
             14'h9ad 	:	val_out <= 16'h3c3c;
             14'h9ae 	:	val_out <= 16'h3c42;
             14'h9af 	:	val_out <= 16'h3c48;
             14'h9b0 	:	val_out <= 16'h3c4e;
             14'h9b1 	:	val_out <= 16'h3c55;
             14'h9b2 	:	val_out <= 16'h3c5b;
             14'h9b3 	:	val_out <= 16'h3c61;
             14'h9b4 	:	val_out <= 16'h3c67;
             14'h9b5 	:	val_out <= 16'h3c6d;
             14'h9b6 	:	val_out <= 16'h3c73;
             14'h9b7 	:	val_out <= 16'h3c79;
             14'h9b8 	:	val_out <= 16'h3c7f;
             14'h9b9 	:	val_out <= 16'h3c85;
             14'h9ba 	:	val_out <= 16'h3c8c;
             14'h9bb 	:	val_out <= 16'h3c92;
             14'h9bc 	:	val_out <= 16'h3c98;
             14'h9bd 	:	val_out <= 16'h3c9e;
             14'h9be 	:	val_out <= 16'h3ca4;
             14'h9bf 	:	val_out <= 16'h3caa;
             14'h9c0 	:	val_out <= 16'h3cb0;
             14'h9c1 	:	val_out <= 16'h3cb6;
             14'h9c2 	:	val_out <= 16'h3cbc;
             14'h9c3 	:	val_out <= 16'h3cc2;
             14'h9c4 	:	val_out <= 16'h3cc9;
             14'h9c5 	:	val_out <= 16'h3ccf;
             14'h9c6 	:	val_out <= 16'h3cd5;
             14'h9c7 	:	val_out <= 16'h3cdb;
             14'h9c8 	:	val_out <= 16'h3ce1;
             14'h9c9 	:	val_out <= 16'h3ce7;
             14'h9ca 	:	val_out <= 16'h3ced;
             14'h9cb 	:	val_out <= 16'h3cf3;
             14'h9cc 	:	val_out <= 16'h3cf9;
             14'h9cd 	:	val_out <= 16'h3cff;
             14'h9ce 	:	val_out <= 16'h3d06;
             14'h9cf 	:	val_out <= 16'h3d0c;
             14'h9d0 	:	val_out <= 16'h3d12;
             14'h9d1 	:	val_out <= 16'h3d18;
             14'h9d2 	:	val_out <= 16'h3d1e;
             14'h9d3 	:	val_out <= 16'h3d24;
             14'h9d4 	:	val_out <= 16'h3d2a;
             14'h9d5 	:	val_out <= 16'h3d30;
             14'h9d6 	:	val_out <= 16'h3d36;
             14'h9d7 	:	val_out <= 16'h3d3c;
             14'h9d8 	:	val_out <= 16'h3d43;
             14'h9d9 	:	val_out <= 16'h3d49;
             14'h9da 	:	val_out <= 16'h3d4f;
             14'h9db 	:	val_out <= 16'h3d55;
             14'h9dc 	:	val_out <= 16'h3d5b;
             14'h9dd 	:	val_out <= 16'h3d61;
             14'h9de 	:	val_out <= 16'h3d67;
             14'h9df 	:	val_out <= 16'h3d6d;
             14'h9e0 	:	val_out <= 16'h3d73;
             14'h9e1 	:	val_out <= 16'h3d79;
             14'h9e2 	:	val_out <= 16'h3d80;
             14'h9e3 	:	val_out <= 16'h3d86;
             14'h9e4 	:	val_out <= 16'h3d8c;
             14'h9e5 	:	val_out <= 16'h3d92;
             14'h9e6 	:	val_out <= 16'h3d98;
             14'h9e7 	:	val_out <= 16'h3d9e;
             14'h9e8 	:	val_out <= 16'h3da4;
             14'h9e9 	:	val_out <= 16'h3daa;
             14'h9ea 	:	val_out <= 16'h3db0;
             14'h9eb 	:	val_out <= 16'h3db6;
             14'h9ec 	:	val_out <= 16'h3dbd;
             14'h9ed 	:	val_out <= 16'h3dc3;
             14'h9ee 	:	val_out <= 16'h3dc9;
             14'h9ef 	:	val_out <= 16'h3dcf;
             14'h9f0 	:	val_out <= 16'h3dd5;
             14'h9f1 	:	val_out <= 16'h3ddb;
             14'h9f2 	:	val_out <= 16'h3de1;
             14'h9f3 	:	val_out <= 16'h3de7;
             14'h9f4 	:	val_out <= 16'h3ded;
             14'h9f5 	:	val_out <= 16'h3df3;
             14'h9f6 	:	val_out <= 16'h3dfa;
             14'h9f7 	:	val_out <= 16'h3e00;
             14'h9f8 	:	val_out <= 16'h3e06;
             14'h9f9 	:	val_out <= 16'h3e0c;
             14'h9fa 	:	val_out <= 16'h3e12;
             14'h9fb 	:	val_out <= 16'h3e18;
             14'h9fc 	:	val_out <= 16'h3e1e;
             14'h9fd 	:	val_out <= 16'h3e24;
             14'h9fe 	:	val_out <= 16'h3e2a;
             14'h9ff 	:	val_out <= 16'h3e30;
             14'ha00 	:	val_out <= 16'h3e36;
             14'ha01 	:	val_out <= 16'h3e3d;
             14'ha02 	:	val_out <= 16'h3e43;
             14'ha03 	:	val_out <= 16'h3e49;
             14'ha04 	:	val_out <= 16'h3e4f;
             14'ha05 	:	val_out <= 16'h3e55;
             14'ha06 	:	val_out <= 16'h3e5b;
             14'ha07 	:	val_out <= 16'h3e61;
             14'ha08 	:	val_out <= 16'h3e67;
             14'ha09 	:	val_out <= 16'h3e6d;
             14'ha0a 	:	val_out <= 16'h3e73;
             14'ha0b 	:	val_out <= 16'h3e7a;
             14'ha0c 	:	val_out <= 16'h3e80;
             14'ha0d 	:	val_out <= 16'h3e86;
             14'ha0e 	:	val_out <= 16'h3e8c;
             14'ha0f 	:	val_out <= 16'h3e92;
             14'ha10 	:	val_out <= 16'h3e98;
             14'ha11 	:	val_out <= 16'h3e9e;
             14'ha12 	:	val_out <= 16'h3ea4;
             14'ha13 	:	val_out <= 16'h3eaa;
             14'ha14 	:	val_out <= 16'h3eb0;
             14'ha15 	:	val_out <= 16'h3eb6;
             14'ha16 	:	val_out <= 16'h3ebd;
             14'ha17 	:	val_out <= 16'h3ec3;
             14'ha18 	:	val_out <= 16'h3ec9;
             14'ha19 	:	val_out <= 16'h3ecf;
             14'ha1a 	:	val_out <= 16'h3ed5;
             14'ha1b 	:	val_out <= 16'h3edb;
             14'ha1c 	:	val_out <= 16'h3ee1;
             14'ha1d 	:	val_out <= 16'h3ee7;
             14'ha1e 	:	val_out <= 16'h3eed;
             14'ha1f 	:	val_out <= 16'h3ef3;
             14'ha20 	:	val_out <= 16'h3ef9;
             14'ha21 	:	val_out <= 16'h3f00;
             14'ha22 	:	val_out <= 16'h3f06;
             14'ha23 	:	val_out <= 16'h3f0c;
             14'ha24 	:	val_out <= 16'h3f12;
             14'ha25 	:	val_out <= 16'h3f18;
             14'ha26 	:	val_out <= 16'h3f1e;
             14'ha27 	:	val_out <= 16'h3f24;
             14'ha28 	:	val_out <= 16'h3f2a;
             14'ha29 	:	val_out <= 16'h3f30;
             14'ha2a 	:	val_out <= 16'h3f36;
             14'ha2b 	:	val_out <= 16'h3f3c;
             14'ha2c 	:	val_out <= 16'h3f43;
             14'ha2d 	:	val_out <= 16'h3f49;
             14'ha2e 	:	val_out <= 16'h3f4f;
             14'ha2f 	:	val_out <= 16'h3f55;
             14'ha30 	:	val_out <= 16'h3f5b;
             14'ha31 	:	val_out <= 16'h3f61;
             14'ha32 	:	val_out <= 16'h3f67;
             14'ha33 	:	val_out <= 16'h3f6d;
             14'ha34 	:	val_out <= 16'h3f73;
             14'ha35 	:	val_out <= 16'h3f79;
             14'ha36 	:	val_out <= 16'h3f7f;
             14'ha37 	:	val_out <= 16'h3f85;
             14'ha38 	:	val_out <= 16'h3f8c;
             14'ha39 	:	val_out <= 16'h3f92;
             14'ha3a 	:	val_out <= 16'h3f98;
             14'ha3b 	:	val_out <= 16'h3f9e;
             14'ha3c 	:	val_out <= 16'h3fa4;
             14'ha3d 	:	val_out <= 16'h3faa;
             14'ha3e 	:	val_out <= 16'h3fb0;
             14'ha3f 	:	val_out <= 16'h3fb6;
             14'ha40 	:	val_out <= 16'h3fbc;
             14'ha41 	:	val_out <= 16'h3fc2;
             14'ha42 	:	val_out <= 16'h3fc8;
             14'ha43 	:	val_out <= 16'h3fcf;
             14'ha44 	:	val_out <= 16'h3fd5;
             14'ha45 	:	val_out <= 16'h3fdb;
             14'ha46 	:	val_out <= 16'h3fe1;
             14'ha47 	:	val_out <= 16'h3fe7;
             14'ha48 	:	val_out <= 16'h3fed;
             14'ha49 	:	val_out <= 16'h3ff3;
             14'ha4a 	:	val_out <= 16'h3ff9;
             14'ha4b 	:	val_out <= 16'h3fff;
             14'ha4c 	:	val_out <= 16'h4005;
             14'ha4d 	:	val_out <= 16'h400b;
             14'ha4e 	:	val_out <= 16'h4011;
             14'ha4f 	:	val_out <= 16'h4018;
             14'ha50 	:	val_out <= 16'h401e;
             14'ha51 	:	val_out <= 16'h4024;
             14'ha52 	:	val_out <= 16'h402a;
             14'ha53 	:	val_out <= 16'h4030;
             14'ha54 	:	val_out <= 16'h4036;
             14'ha55 	:	val_out <= 16'h403c;
             14'ha56 	:	val_out <= 16'h4042;
             14'ha57 	:	val_out <= 16'h4048;
             14'ha58 	:	val_out <= 16'h404e;
             14'ha59 	:	val_out <= 16'h4054;
             14'ha5a 	:	val_out <= 16'h405a;
             14'ha5b 	:	val_out <= 16'h4061;
             14'ha5c 	:	val_out <= 16'h4067;
             14'ha5d 	:	val_out <= 16'h406d;
             14'ha5e 	:	val_out <= 16'h4073;
             14'ha5f 	:	val_out <= 16'h4079;
             14'ha60 	:	val_out <= 16'h407f;
             14'ha61 	:	val_out <= 16'h4085;
             14'ha62 	:	val_out <= 16'h408b;
             14'ha63 	:	val_out <= 16'h4091;
             14'ha64 	:	val_out <= 16'h4097;
             14'ha65 	:	val_out <= 16'h409d;
             14'ha66 	:	val_out <= 16'h40a3;
             14'ha67 	:	val_out <= 16'h40a9;
             14'ha68 	:	val_out <= 16'h40b0;
             14'ha69 	:	val_out <= 16'h40b6;
             14'ha6a 	:	val_out <= 16'h40bc;
             14'ha6b 	:	val_out <= 16'h40c2;
             14'ha6c 	:	val_out <= 16'h40c8;
             14'ha6d 	:	val_out <= 16'h40ce;
             14'ha6e 	:	val_out <= 16'h40d4;
             14'ha6f 	:	val_out <= 16'h40da;
             14'ha70 	:	val_out <= 16'h40e0;
             14'ha71 	:	val_out <= 16'h40e6;
             14'ha72 	:	val_out <= 16'h40ec;
             14'ha73 	:	val_out <= 16'h40f2;
             14'ha74 	:	val_out <= 16'h40f8;
             14'ha75 	:	val_out <= 16'h40ff;
             14'ha76 	:	val_out <= 16'h4105;
             14'ha77 	:	val_out <= 16'h410b;
             14'ha78 	:	val_out <= 16'h4111;
             14'ha79 	:	val_out <= 16'h4117;
             14'ha7a 	:	val_out <= 16'h411d;
             14'ha7b 	:	val_out <= 16'h4123;
             14'ha7c 	:	val_out <= 16'h4129;
             14'ha7d 	:	val_out <= 16'h412f;
             14'ha7e 	:	val_out <= 16'h4135;
             14'ha7f 	:	val_out <= 16'h413b;
             14'ha80 	:	val_out <= 16'h4141;
             14'ha81 	:	val_out <= 16'h4147;
             14'ha82 	:	val_out <= 16'h414e;
             14'ha83 	:	val_out <= 16'h4154;
             14'ha84 	:	val_out <= 16'h415a;
             14'ha85 	:	val_out <= 16'h4160;
             14'ha86 	:	val_out <= 16'h4166;
             14'ha87 	:	val_out <= 16'h416c;
             14'ha88 	:	val_out <= 16'h4172;
             14'ha89 	:	val_out <= 16'h4178;
             14'ha8a 	:	val_out <= 16'h417e;
             14'ha8b 	:	val_out <= 16'h4184;
             14'ha8c 	:	val_out <= 16'h418a;
             14'ha8d 	:	val_out <= 16'h4190;
             14'ha8e 	:	val_out <= 16'h4196;
             14'ha8f 	:	val_out <= 16'h419d;
             14'ha90 	:	val_out <= 16'h41a3;
             14'ha91 	:	val_out <= 16'h41a9;
             14'ha92 	:	val_out <= 16'h41af;
             14'ha93 	:	val_out <= 16'h41b5;
             14'ha94 	:	val_out <= 16'h41bb;
             14'ha95 	:	val_out <= 16'h41c1;
             14'ha96 	:	val_out <= 16'h41c7;
             14'ha97 	:	val_out <= 16'h41cd;
             14'ha98 	:	val_out <= 16'h41d3;
             14'ha99 	:	val_out <= 16'h41d9;
             14'ha9a 	:	val_out <= 16'h41df;
             14'ha9b 	:	val_out <= 16'h41e5;
             14'ha9c 	:	val_out <= 16'h41eb;
             14'ha9d 	:	val_out <= 16'h41f2;
             14'ha9e 	:	val_out <= 16'h41f8;
             14'ha9f 	:	val_out <= 16'h41fe;
             14'haa0 	:	val_out <= 16'h4204;
             14'haa1 	:	val_out <= 16'h420a;
             14'haa2 	:	val_out <= 16'h4210;
             14'haa3 	:	val_out <= 16'h4216;
             14'haa4 	:	val_out <= 16'h421c;
             14'haa5 	:	val_out <= 16'h4222;
             14'haa6 	:	val_out <= 16'h4228;
             14'haa7 	:	val_out <= 16'h422e;
             14'haa8 	:	val_out <= 16'h4234;
             14'haa9 	:	val_out <= 16'h423a;
             14'haaa 	:	val_out <= 16'h4240;
             14'haab 	:	val_out <= 16'h4247;
             14'haac 	:	val_out <= 16'h424d;
             14'haad 	:	val_out <= 16'h4253;
             14'haae 	:	val_out <= 16'h4259;
             14'haaf 	:	val_out <= 16'h425f;
             14'hab0 	:	val_out <= 16'h4265;
             14'hab1 	:	val_out <= 16'h426b;
             14'hab2 	:	val_out <= 16'h4271;
             14'hab3 	:	val_out <= 16'h4277;
             14'hab4 	:	val_out <= 16'h427d;
             14'hab5 	:	val_out <= 16'h4283;
             14'hab6 	:	val_out <= 16'h4289;
             14'hab7 	:	val_out <= 16'h428f;
             14'hab8 	:	val_out <= 16'h4295;
             14'hab9 	:	val_out <= 16'h429b;
             14'haba 	:	val_out <= 16'h42a2;
             14'habb 	:	val_out <= 16'h42a8;
             14'habc 	:	val_out <= 16'h42ae;
             14'habd 	:	val_out <= 16'h42b4;
             14'habe 	:	val_out <= 16'h42ba;
             14'habf 	:	val_out <= 16'h42c0;
             14'hac0 	:	val_out <= 16'h42c6;
             14'hac1 	:	val_out <= 16'h42cc;
             14'hac2 	:	val_out <= 16'h42d2;
             14'hac3 	:	val_out <= 16'h42d8;
             14'hac4 	:	val_out <= 16'h42de;
             14'hac5 	:	val_out <= 16'h42e4;
             14'hac6 	:	val_out <= 16'h42ea;
             14'hac7 	:	val_out <= 16'h42f0;
             14'hac8 	:	val_out <= 16'h42f6;
             14'hac9 	:	val_out <= 16'h42fd;
             14'haca 	:	val_out <= 16'h4303;
             14'hacb 	:	val_out <= 16'h4309;
             14'hacc 	:	val_out <= 16'h430f;
             14'hacd 	:	val_out <= 16'h4315;
             14'hace 	:	val_out <= 16'h431b;
             14'hacf 	:	val_out <= 16'h4321;
             14'had0 	:	val_out <= 16'h4327;
             14'had1 	:	val_out <= 16'h432d;
             14'had2 	:	val_out <= 16'h4333;
             14'had3 	:	val_out <= 16'h4339;
             14'had4 	:	val_out <= 16'h433f;
             14'had5 	:	val_out <= 16'h4345;
             14'had6 	:	val_out <= 16'h434b;
             14'had7 	:	val_out <= 16'h4351;
             14'had8 	:	val_out <= 16'h4357;
             14'had9 	:	val_out <= 16'h435e;
             14'hada 	:	val_out <= 16'h4364;
             14'hadb 	:	val_out <= 16'h436a;
             14'hadc 	:	val_out <= 16'h4370;
             14'hadd 	:	val_out <= 16'h4376;
             14'hade 	:	val_out <= 16'h437c;
             14'hadf 	:	val_out <= 16'h4382;
             14'hae0 	:	val_out <= 16'h4388;
             14'hae1 	:	val_out <= 16'h438e;
             14'hae2 	:	val_out <= 16'h4394;
             14'hae3 	:	val_out <= 16'h439a;
             14'hae4 	:	val_out <= 16'h43a0;
             14'hae5 	:	val_out <= 16'h43a6;
             14'hae6 	:	val_out <= 16'h43ac;
             14'hae7 	:	val_out <= 16'h43b2;
             14'hae8 	:	val_out <= 16'h43b8;
             14'hae9 	:	val_out <= 16'h43be;
             14'haea 	:	val_out <= 16'h43c5;
             14'haeb 	:	val_out <= 16'h43cb;
             14'haec 	:	val_out <= 16'h43d1;
             14'haed 	:	val_out <= 16'h43d7;
             14'haee 	:	val_out <= 16'h43dd;
             14'haef 	:	val_out <= 16'h43e3;
             14'haf0 	:	val_out <= 16'h43e9;
             14'haf1 	:	val_out <= 16'h43ef;
             14'haf2 	:	val_out <= 16'h43f5;
             14'haf3 	:	val_out <= 16'h43fb;
             14'haf4 	:	val_out <= 16'h4401;
             14'haf5 	:	val_out <= 16'h4407;
             14'haf6 	:	val_out <= 16'h440d;
             14'haf7 	:	val_out <= 16'h4413;
             14'haf8 	:	val_out <= 16'h4419;
             14'haf9 	:	val_out <= 16'h441f;
             14'hafa 	:	val_out <= 16'h4425;
             14'hafb 	:	val_out <= 16'h442c;
             14'hafc 	:	val_out <= 16'h4432;
             14'hafd 	:	val_out <= 16'h4438;
             14'hafe 	:	val_out <= 16'h443e;
             14'haff 	:	val_out <= 16'h4444;
             14'hb00 	:	val_out <= 16'h444a;
             14'hb01 	:	val_out <= 16'h4450;
             14'hb02 	:	val_out <= 16'h4456;
             14'hb03 	:	val_out <= 16'h445c;
             14'hb04 	:	val_out <= 16'h4462;
             14'hb05 	:	val_out <= 16'h4468;
             14'hb06 	:	val_out <= 16'h446e;
             14'hb07 	:	val_out <= 16'h4474;
             14'hb08 	:	val_out <= 16'h447a;
             14'hb09 	:	val_out <= 16'h4480;
             14'hb0a 	:	val_out <= 16'h4486;
             14'hb0b 	:	val_out <= 16'h448c;
             14'hb0c 	:	val_out <= 16'h4492;
             14'hb0d 	:	val_out <= 16'h4499;
             14'hb0e 	:	val_out <= 16'h449f;
             14'hb0f 	:	val_out <= 16'h44a5;
             14'hb10 	:	val_out <= 16'h44ab;
             14'hb11 	:	val_out <= 16'h44b1;
             14'hb12 	:	val_out <= 16'h44b7;
             14'hb13 	:	val_out <= 16'h44bd;
             14'hb14 	:	val_out <= 16'h44c3;
             14'hb15 	:	val_out <= 16'h44c9;
             14'hb16 	:	val_out <= 16'h44cf;
             14'hb17 	:	val_out <= 16'h44d5;
             14'hb18 	:	val_out <= 16'h44db;
             14'hb19 	:	val_out <= 16'h44e1;
             14'hb1a 	:	val_out <= 16'h44e7;
             14'hb1b 	:	val_out <= 16'h44ed;
             14'hb1c 	:	val_out <= 16'h44f3;
             14'hb1d 	:	val_out <= 16'h44f9;
             14'hb1e 	:	val_out <= 16'h44ff;
             14'hb1f 	:	val_out <= 16'h4505;
             14'hb20 	:	val_out <= 16'h450c;
             14'hb21 	:	val_out <= 16'h4512;
             14'hb22 	:	val_out <= 16'h4518;
             14'hb23 	:	val_out <= 16'h451e;
             14'hb24 	:	val_out <= 16'h4524;
             14'hb25 	:	val_out <= 16'h452a;
             14'hb26 	:	val_out <= 16'h4530;
             14'hb27 	:	val_out <= 16'h4536;
             14'hb28 	:	val_out <= 16'h453c;
             14'hb29 	:	val_out <= 16'h4542;
             14'hb2a 	:	val_out <= 16'h4548;
             14'hb2b 	:	val_out <= 16'h454e;
             14'hb2c 	:	val_out <= 16'h4554;
             14'hb2d 	:	val_out <= 16'h455a;
             14'hb2e 	:	val_out <= 16'h4560;
             14'hb2f 	:	val_out <= 16'h4566;
             14'hb30 	:	val_out <= 16'h456c;
             14'hb31 	:	val_out <= 16'h4572;
             14'hb32 	:	val_out <= 16'h4578;
             14'hb33 	:	val_out <= 16'h457e;
             14'hb34 	:	val_out <= 16'h4584;
             14'hb35 	:	val_out <= 16'h458b;
             14'hb36 	:	val_out <= 16'h4591;
             14'hb37 	:	val_out <= 16'h4597;
             14'hb38 	:	val_out <= 16'h459d;
             14'hb39 	:	val_out <= 16'h45a3;
             14'hb3a 	:	val_out <= 16'h45a9;
             14'hb3b 	:	val_out <= 16'h45af;
             14'hb3c 	:	val_out <= 16'h45b5;
             14'hb3d 	:	val_out <= 16'h45bb;
             14'hb3e 	:	val_out <= 16'h45c1;
             14'hb3f 	:	val_out <= 16'h45c7;
             14'hb40 	:	val_out <= 16'h45cd;
             14'hb41 	:	val_out <= 16'h45d3;
             14'hb42 	:	val_out <= 16'h45d9;
             14'hb43 	:	val_out <= 16'h45df;
             14'hb44 	:	val_out <= 16'h45e5;
             14'hb45 	:	val_out <= 16'h45eb;
             14'hb46 	:	val_out <= 16'h45f1;
             14'hb47 	:	val_out <= 16'h45f7;
             14'hb48 	:	val_out <= 16'h45fd;
             14'hb49 	:	val_out <= 16'h4603;
             14'hb4a 	:	val_out <= 16'h4609;
             14'hb4b 	:	val_out <= 16'h4610;
             14'hb4c 	:	val_out <= 16'h4616;
             14'hb4d 	:	val_out <= 16'h461c;
             14'hb4e 	:	val_out <= 16'h4622;
             14'hb4f 	:	val_out <= 16'h4628;
             14'hb50 	:	val_out <= 16'h462e;
             14'hb51 	:	val_out <= 16'h4634;
             14'hb52 	:	val_out <= 16'h463a;
             14'hb53 	:	val_out <= 16'h4640;
             14'hb54 	:	val_out <= 16'h4646;
             14'hb55 	:	val_out <= 16'h464c;
             14'hb56 	:	val_out <= 16'h4652;
             14'hb57 	:	val_out <= 16'h4658;
             14'hb58 	:	val_out <= 16'h465e;
             14'hb59 	:	val_out <= 16'h4664;
             14'hb5a 	:	val_out <= 16'h466a;
             14'hb5b 	:	val_out <= 16'h4670;
             14'hb5c 	:	val_out <= 16'h4676;
             14'hb5d 	:	val_out <= 16'h467c;
             14'hb5e 	:	val_out <= 16'h4682;
             14'hb5f 	:	val_out <= 16'h4688;
             14'hb60 	:	val_out <= 16'h468e;
             14'hb61 	:	val_out <= 16'h4694;
             14'hb62 	:	val_out <= 16'h469a;
             14'hb63 	:	val_out <= 16'h46a1;
             14'hb64 	:	val_out <= 16'h46a7;
             14'hb65 	:	val_out <= 16'h46ad;
             14'hb66 	:	val_out <= 16'h46b3;
             14'hb67 	:	val_out <= 16'h46b9;
             14'hb68 	:	val_out <= 16'h46bf;
             14'hb69 	:	val_out <= 16'h46c5;
             14'hb6a 	:	val_out <= 16'h46cb;
             14'hb6b 	:	val_out <= 16'h46d1;
             14'hb6c 	:	val_out <= 16'h46d7;
             14'hb6d 	:	val_out <= 16'h46dd;
             14'hb6e 	:	val_out <= 16'h46e3;
             14'hb6f 	:	val_out <= 16'h46e9;
             14'hb70 	:	val_out <= 16'h46ef;
             14'hb71 	:	val_out <= 16'h46f5;
             14'hb72 	:	val_out <= 16'h46fb;
             14'hb73 	:	val_out <= 16'h4701;
             14'hb74 	:	val_out <= 16'h4707;
             14'hb75 	:	val_out <= 16'h470d;
             14'hb76 	:	val_out <= 16'h4713;
             14'hb77 	:	val_out <= 16'h4719;
             14'hb78 	:	val_out <= 16'h471f;
             14'hb79 	:	val_out <= 16'h4725;
             14'hb7a 	:	val_out <= 16'h472b;
             14'hb7b 	:	val_out <= 16'h4731;
             14'hb7c 	:	val_out <= 16'h4737;
             14'hb7d 	:	val_out <= 16'h473d;
             14'hb7e 	:	val_out <= 16'h4744;
             14'hb7f 	:	val_out <= 16'h474a;
             14'hb80 	:	val_out <= 16'h4750;
             14'hb81 	:	val_out <= 16'h4756;
             14'hb82 	:	val_out <= 16'h475c;
             14'hb83 	:	val_out <= 16'h4762;
             14'hb84 	:	val_out <= 16'h4768;
             14'hb85 	:	val_out <= 16'h476e;
             14'hb86 	:	val_out <= 16'h4774;
             14'hb87 	:	val_out <= 16'h477a;
             14'hb88 	:	val_out <= 16'h4780;
             14'hb89 	:	val_out <= 16'h4786;
             14'hb8a 	:	val_out <= 16'h478c;
             14'hb8b 	:	val_out <= 16'h4792;
             14'hb8c 	:	val_out <= 16'h4798;
             14'hb8d 	:	val_out <= 16'h479e;
             14'hb8e 	:	val_out <= 16'h47a4;
             14'hb8f 	:	val_out <= 16'h47aa;
             14'hb90 	:	val_out <= 16'h47b0;
             14'hb91 	:	val_out <= 16'h47b6;
             14'hb92 	:	val_out <= 16'h47bc;
             14'hb93 	:	val_out <= 16'h47c2;
             14'hb94 	:	val_out <= 16'h47c8;
             14'hb95 	:	val_out <= 16'h47ce;
             14'hb96 	:	val_out <= 16'h47d4;
             14'hb97 	:	val_out <= 16'h47da;
             14'hb98 	:	val_out <= 16'h47e0;
             14'hb99 	:	val_out <= 16'h47e6;
             14'hb9a 	:	val_out <= 16'h47ec;
             14'hb9b 	:	val_out <= 16'h47f2;
             14'hb9c 	:	val_out <= 16'h47f8;
             14'hb9d 	:	val_out <= 16'h47ff;
             14'hb9e 	:	val_out <= 16'h4805;
             14'hb9f 	:	val_out <= 16'h480b;
             14'hba0 	:	val_out <= 16'h4811;
             14'hba1 	:	val_out <= 16'h4817;
             14'hba2 	:	val_out <= 16'h481d;
             14'hba3 	:	val_out <= 16'h4823;
             14'hba4 	:	val_out <= 16'h4829;
             14'hba5 	:	val_out <= 16'h482f;
             14'hba6 	:	val_out <= 16'h4835;
             14'hba7 	:	val_out <= 16'h483b;
             14'hba8 	:	val_out <= 16'h4841;
             14'hba9 	:	val_out <= 16'h4847;
             14'hbaa 	:	val_out <= 16'h484d;
             14'hbab 	:	val_out <= 16'h4853;
             14'hbac 	:	val_out <= 16'h4859;
             14'hbad 	:	val_out <= 16'h485f;
             14'hbae 	:	val_out <= 16'h4865;
             14'hbaf 	:	val_out <= 16'h486b;
             14'hbb0 	:	val_out <= 16'h4871;
             14'hbb1 	:	val_out <= 16'h4877;
             14'hbb2 	:	val_out <= 16'h487d;
             14'hbb3 	:	val_out <= 16'h4883;
             14'hbb4 	:	val_out <= 16'h4889;
             14'hbb5 	:	val_out <= 16'h488f;
             14'hbb6 	:	val_out <= 16'h4895;
             14'hbb7 	:	val_out <= 16'h489b;
             14'hbb8 	:	val_out <= 16'h48a1;
             14'hbb9 	:	val_out <= 16'h48a7;
             14'hbba 	:	val_out <= 16'h48ad;
             14'hbbb 	:	val_out <= 16'h48b3;
             14'hbbc 	:	val_out <= 16'h48b9;
             14'hbbd 	:	val_out <= 16'h48bf;
             14'hbbe 	:	val_out <= 16'h48c5;
             14'hbbf 	:	val_out <= 16'h48cb;
             14'hbc0 	:	val_out <= 16'h48d1;
             14'hbc1 	:	val_out <= 16'h48d7;
             14'hbc2 	:	val_out <= 16'h48dd;
             14'hbc3 	:	val_out <= 16'h48e4;
             14'hbc4 	:	val_out <= 16'h48ea;
             14'hbc5 	:	val_out <= 16'h48f0;
             14'hbc6 	:	val_out <= 16'h48f6;
             14'hbc7 	:	val_out <= 16'h48fc;
             14'hbc8 	:	val_out <= 16'h4902;
             14'hbc9 	:	val_out <= 16'h4908;
             14'hbca 	:	val_out <= 16'h490e;
             14'hbcb 	:	val_out <= 16'h4914;
             14'hbcc 	:	val_out <= 16'h491a;
             14'hbcd 	:	val_out <= 16'h4920;
             14'hbce 	:	val_out <= 16'h4926;
             14'hbcf 	:	val_out <= 16'h492c;
             14'hbd0 	:	val_out <= 16'h4932;
             14'hbd1 	:	val_out <= 16'h4938;
             14'hbd2 	:	val_out <= 16'h493e;
             14'hbd3 	:	val_out <= 16'h4944;
             14'hbd4 	:	val_out <= 16'h494a;
             14'hbd5 	:	val_out <= 16'h4950;
             14'hbd6 	:	val_out <= 16'h4956;
             14'hbd7 	:	val_out <= 16'h495c;
             14'hbd8 	:	val_out <= 16'h4962;
             14'hbd9 	:	val_out <= 16'h4968;
             14'hbda 	:	val_out <= 16'h496e;
             14'hbdb 	:	val_out <= 16'h4974;
             14'hbdc 	:	val_out <= 16'h497a;
             14'hbdd 	:	val_out <= 16'h4980;
             14'hbde 	:	val_out <= 16'h4986;
             14'hbdf 	:	val_out <= 16'h498c;
             14'hbe0 	:	val_out <= 16'h4992;
             14'hbe1 	:	val_out <= 16'h4998;
             14'hbe2 	:	val_out <= 16'h499e;
             14'hbe3 	:	val_out <= 16'h49a4;
             14'hbe4 	:	val_out <= 16'h49aa;
             14'hbe5 	:	val_out <= 16'h49b0;
             14'hbe6 	:	val_out <= 16'h49b6;
             14'hbe7 	:	val_out <= 16'h49bc;
             14'hbe8 	:	val_out <= 16'h49c2;
             14'hbe9 	:	val_out <= 16'h49c8;
             14'hbea 	:	val_out <= 16'h49ce;
             14'hbeb 	:	val_out <= 16'h49d4;
             14'hbec 	:	val_out <= 16'h49da;
             14'hbed 	:	val_out <= 16'h49e0;
             14'hbee 	:	val_out <= 16'h49e6;
             14'hbef 	:	val_out <= 16'h49ec;
             14'hbf0 	:	val_out <= 16'h49f2;
             14'hbf1 	:	val_out <= 16'h49f8;
             14'hbf2 	:	val_out <= 16'h49fe;
             14'hbf3 	:	val_out <= 16'h4a04;
             14'hbf4 	:	val_out <= 16'h4a0a;
             14'hbf5 	:	val_out <= 16'h4a10;
             14'hbf6 	:	val_out <= 16'h4a16;
             14'hbf7 	:	val_out <= 16'h4a1c;
             14'hbf8 	:	val_out <= 16'h4a22;
             14'hbf9 	:	val_out <= 16'h4a29;
             14'hbfa 	:	val_out <= 16'h4a2f;
             14'hbfb 	:	val_out <= 16'h4a35;
             14'hbfc 	:	val_out <= 16'h4a3b;
             14'hbfd 	:	val_out <= 16'h4a41;
             14'hbfe 	:	val_out <= 16'h4a47;
             14'hbff 	:	val_out <= 16'h4a4d;
             14'hc00 	:	val_out <= 16'h4a53;
             14'hc01 	:	val_out <= 16'h4a59;
             14'hc02 	:	val_out <= 16'h4a5f;
             14'hc03 	:	val_out <= 16'h4a65;
             14'hc04 	:	val_out <= 16'h4a6b;
             14'hc05 	:	val_out <= 16'h4a71;
             14'hc06 	:	val_out <= 16'h4a77;
             14'hc07 	:	val_out <= 16'h4a7d;
             14'hc08 	:	val_out <= 16'h4a83;
             14'hc09 	:	val_out <= 16'h4a89;
             14'hc0a 	:	val_out <= 16'h4a8f;
             14'hc0b 	:	val_out <= 16'h4a95;
             14'hc0c 	:	val_out <= 16'h4a9b;
             14'hc0d 	:	val_out <= 16'h4aa1;
             14'hc0e 	:	val_out <= 16'h4aa7;
             14'hc0f 	:	val_out <= 16'h4aad;
             14'hc10 	:	val_out <= 16'h4ab3;
             14'hc11 	:	val_out <= 16'h4ab9;
             14'hc12 	:	val_out <= 16'h4abf;
             14'hc13 	:	val_out <= 16'h4ac5;
             14'hc14 	:	val_out <= 16'h4acb;
             14'hc15 	:	val_out <= 16'h4ad1;
             14'hc16 	:	val_out <= 16'h4ad7;
             14'hc17 	:	val_out <= 16'h4add;
             14'hc18 	:	val_out <= 16'h4ae3;
             14'hc19 	:	val_out <= 16'h4ae9;
             14'hc1a 	:	val_out <= 16'h4aef;
             14'hc1b 	:	val_out <= 16'h4af5;
             14'hc1c 	:	val_out <= 16'h4afb;
             14'hc1d 	:	val_out <= 16'h4b01;
             14'hc1e 	:	val_out <= 16'h4b07;
             14'hc1f 	:	val_out <= 16'h4b0d;
             14'hc20 	:	val_out <= 16'h4b13;
             14'hc21 	:	val_out <= 16'h4b19;
             14'hc22 	:	val_out <= 16'h4b1f;
             14'hc23 	:	val_out <= 16'h4b25;
             14'hc24 	:	val_out <= 16'h4b2b;
             14'hc25 	:	val_out <= 16'h4b31;
             14'hc26 	:	val_out <= 16'h4b37;
             14'hc27 	:	val_out <= 16'h4b3d;
             14'hc28 	:	val_out <= 16'h4b43;
             14'hc29 	:	val_out <= 16'h4b49;
             14'hc2a 	:	val_out <= 16'h4b4f;
             14'hc2b 	:	val_out <= 16'h4b55;
             14'hc2c 	:	val_out <= 16'h4b5b;
             14'hc2d 	:	val_out <= 16'h4b61;
             14'hc2e 	:	val_out <= 16'h4b67;
             14'hc2f 	:	val_out <= 16'h4b6d;
             14'hc30 	:	val_out <= 16'h4b73;
             14'hc31 	:	val_out <= 16'h4b79;
             14'hc32 	:	val_out <= 16'h4b7f;
             14'hc33 	:	val_out <= 16'h4b85;
             14'hc34 	:	val_out <= 16'h4b8b;
             14'hc35 	:	val_out <= 16'h4b91;
             14'hc36 	:	val_out <= 16'h4b97;
             14'hc37 	:	val_out <= 16'h4b9d;
             14'hc38 	:	val_out <= 16'h4ba3;
             14'hc39 	:	val_out <= 16'h4ba9;
             14'hc3a 	:	val_out <= 16'h4baf;
             14'hc3b 	:	val_out <= 16'h4bb5;
             14'hc3c 	:	val_out <= 16'h4bbb;
             14'hc3d 	:	val_out <= 16'h4bc1;
             14'hc3e 	:	val_out <= 16'h4bc7;
             14'hc3f 	:	val_out <= 16'h4bcd;
             14'hc40 	:	val_out <= 16'h4bd3;
             14'hc41 	:	val_out <= 16'h4bd9;
             14'hc42 	:	val_out <= 16'h4bdf;
             14'hc43 	:	val_out <= 16'h4be5;
             14'hc44 	:	val_out <= 16'h4beb;
             14'hc45 	:	val_out <= 16'h4bf1;
             14'hc46 	:	val_out <= 16'h4bf7;
             14'hc47 	:	val_out <= 16'h4bfd;
             14'hc48 	:	val_out <= 16'h4c03;
             14'hc49 	:	val_out <= 16'h4c09;
             14'hc4a 	:	val_out <= 16'h4c0f;
             14'hc4b 	:	val_out <= 16'h4c15;
             14'hc4c 	:	val_out <= 16'h4c1b;
             14'hc4d 	:	val_out <= 16'h4c21;
             14'hc4e 	:	val_out <= 16'h4c27;
             14'hc4f 	:	val_out <= 16'h4c2d;
             14'hc50 	:	val_out <= 16'h4c33;
             14'hc51 	:	val_out <= 16'h4c39;
             14'hc52 	:	val_out <= 16'h4c3f;
             14'hc53 	:	val_out <= 16'h4c45;
             14'hc54 	:	val_out <= 16'h4c4b;
             14'hc55 	:	val_out <= 16'h4c51;
             14'hc56 	:	val_out <= 16'h4c57;
             14'hc57 	:	val_out <= 16'h4c5d;
             14'hc58 	:	val_out <= 16'h4c63;
             14'hc59 	:	val_out <= 16'h4c69;
             14'hc5a 	:	val_out <= 16'h4c6f;
             14'hc5b 	:	val_out <= 16'h4c75;
             14'hc5c 	:	val_out <= 16'h4c7b;
             14'hc5d 	:	val_out <= 16'h4c81;
             14'hc5e 	:	val_out <= 16'h4c87;
             14'hc5f 	:	val_out <= 16'h4c8d;
             14'hc60 	:	val_out <= 16'h4c93;
             14'hc61 	:	val_out <= 16'h4c99;
             14'hc62 	:	val_out <= 16'h4c9f;
             14'hc63 	:	val_out <= 16'h4ca5;
             14'hc64 	:	val_out <= 16'h4cab;
             14'hc65 	:	val_out <= 16'h4cb1;
             14'hc66 	:	val_out <= 16'h4cb7;
             14'hc67 	:	val_out <= 16'h4cbd;
             14'hc68 	:	val_out <= 16'h4cc3;
             14'hc69 	:	val_out <= 16'h4cc9;
             14'hc6a 	:	val_out <= 16'h4ccf;
             14'hc6b 	:	val_out <= 16'h4cd5;
             14'hc6c 	:	val_out <= 16'h4cdb;
             14'hc6d 	:	val_out <= 16'h4ce1;
             14'hc6e 	:	val_out <= 16'h4ce7;
             14'hc6f 	:	val_out <= 16'h4ced;
             14'hc70 	:	val_out <= 16'h4cf3;
             14'hc71 	:	val_out <= 16'h4cf9;
             14'hc72 	:	val_out <= 16'h4cff;
             14'hc73 	:	val_out <= 16'h4d05;
             14'hc74 	:	val_out <= 16'h4d0b;
             14'hc75 	:	val_out <= 16'h4d11;
             14'hc76 	:	val_out <= 16'h4d17;
             14'hc77 	:	val_out <= 16'h4d1d;
             14'hc78 	:	val_out <= 16'h4d23;
             14'hc79 	:	val_out <= 16'h4d29;
             14'hc7a 	:	val_out <= 16'h4d2f;
             14'hc7b 	:	val_out <= 16'h4d35;
             14'hc7c 	:	val_out <= 16'h4d3b;
             14'hc7d 	:	val_out <= 16'h4d41;
             14'hc7e 	:	val_out <= 16'h4d47;
             14'hc7f 	:	val_out <= 16'h4d4d;
             14'hc80 	:	val_out <= 16'h4d53;
             14'hc81 	:	val_out <= 16'h4d59;
             14'hc82 	:	val_out <= 16'h4d5f;
             14'hc83 	:	val_out <= 16'h4d65;
             14'hc84 	:	val_out <= 16'h4d6b;
             14'hc85 	:	val_out <= 16'h4d71;
             14'hc86 	:	val_out <= 16'h4d77;
             14'hc87 	:	val_out <= 16'h4d7d;
             14'hc88 	:	val_out <= 16'h4d83;
             14'hc89 	:	val_out <= 16'h4d89;
             14'hc8a 	:	val_out <= 16'h4d8f;
             14'hc8b 	:	val_out <= 16'h4d95;
             14'hc8c 	:	val_out <= 16'h4d9b;
             14'hc8d 	:	val_out <= 16'h4da1;
             14'hc8e 	:	val_out <= 16'h4da7;
             14'hc8f 	:	val_out <= 16'h4dad;
             14'hc90 	:	val_out <= 16'h4db3;
             14'hc91 	:	val_out <= 16'h4db9;
             14'hc92 	:	val_out <= 16'h4dbf;
             14'hc93 	:	val_out <= 16'h4dc5;
             14'hc94 	:	val_out <= 16'h4dcb;
             14'hc95 	:	val_out <= 16'h4dd1;
             14'hc96 	:	val_out <= 16'h4dd6;
             14'hc97 	:	val_out <= 16'h4ddc;
             14'hc98 	:	val_out <= 16'h4de2;
             14'hc99 	:	val_out <= 16'h4de8;
             14'hc9a 	:	val_out <= 16'h4dee;
             14'hc9b 	:	val_out <= 16'h4df4;
             14'hc9c 	:	val_out <= 16'h4dfa;
             14'hc9d 	:	val_out <= 16'h4e00;
             14'hc9e 	:	val_out <= 16'h4e06;
             14'hc9f 	:	val_out <= 16'h4e0c;
             14'hca0 	:	val_out <= 16'h4e12;
             14'hca1 	:	val_out <= 16'h4e18;
             14'hca2 	:	val_out <= 16'h4e1e;
             14'hca3 	:	val_out <= 16'h4e24;
             14'hca4 	:	val_out <= 16'h4e2a;
             14'hca5 	:	val_out <= 16'h4e30;
             14'hca6 	:	val_out <= 16'h4e36;
             14'hca7 	:	val_out <= 16'h4e3c;
             14'hca8 	:	val_out <= 16'h4e42;
             14'hca9 	:	val_out <= 16'h4e48;
             14'hcaa 	:	val_out <= 16'h4e4e;
             14'hcab 	:	val_out <= 16'h4e54;
             14'hcac 	:	val_out <= 16'h4e5a;
             14'hcad 	:	val_out <= 16'h4e60;
             14'hcae 	:	val_out <= 16'h4e66;
             14'hcaf 	:	val_out <= 16'h4e6c;
             14'hcb0 	:	val_out <= 16'h4e72;
             14'hcb1 	:	val_out <= 16'h4e78;
             14'hcb2 	:	val_out <= 16'h4e7e;
             14'hcb3 	:	val_out <= 16'h4e84;
             14'hcb4 	:	val_out <= 16'h4e8a;
             14'hcb5 	:	val_out <= 16'h4e90;
             14'hcb6 	:	val_out <= 16'h4e96;
             14'hcb7 	:	val_out <= 16'h4e9c;
             14'hcb8 	:	val_out <= 16'h4ea2;
             14'hcb9 	:	val_out <= 16'h4ea8;
             14'hcba 	:	val_out <= 16'h4eae;
             14'hcbb 	:	val_out <= 16'h4eb4;
             14'hcbc 	:	val_out <= 16'h4eba;
             14'hcbd 	:	val_out <= 16'h4ec0;
             14'hcbe 	:	val_out <= 16'h4ec6;
             14'hcbf 	:	val_out <= 16'h4ecc;
             14'hcc0 	:	val_out <= 16'h4ed2;
             14'hcc1 	:	val_out <= 16'h4ed8;
             14'hcc2 	:	val_out <= 16'h4ede;
             14'hcc3 	:	val_out <= 16'h4ee4;
             14'hcc4 	:	val_out <= 16'h4eea;
             14'hcc5 	:	val_out <= 16'h4ef0;
             14'hcc6 	:	val_out <= 16'h4ef6;
             14'hcc7 	:	val_out <= 16'h4efc;
             14'hcc8 	:	val_out <= 16'h4f02;
             14'hcc9 	:	val_out <= 16'h4f08;
             14'hcca 	:	val_out <= 16'h4f0d;
             14'hccb 	:	val_out <= 16'h4f13;
             14'hccc 	:	val_out <= 16'h4f19;
             14'hccd 	:	val_out <= 16'h4f1f;
             14'hcce 	:	val_out <= 16'h4f25;
             14'hccf 	:	val_out <= 16'h4f2b;
             14'hcd0 	:	val_out <= 16'h4f31;
             14'hcd1 	:	val_out <= 16'h4f37;
             14'hcd2 	:	val_out <= 16'h4f3d;
             14'hcd3 	:	val_out <= 16'h4f43;
             14'hcd4 	:	val_out <= 16'h4f49;
             14'hcd5 	:	val_out <= 16'h4f4f;
             14'hcd6 	:	val_out <= 16'h4f55;
             14'hcd7 	:	val_out <= 16'h4f5b;
             14'hcd8 	:	val_out <= 16'h4f61;
             14'hcd9 	:	val_out <= 16'h4f67;
             14'hcda 	:	val_out <= 16'h4f6d;
             14'hcdb 	:	val_out <= 16'h4f73;
             14'hcdc 	:	val_out <= 16'h4f79;
             14'hcdd 	:	val_out <= 16'h4f7f;
             14'hcde 	:	val_out <= 16'h4f85;
             14'hcdf 	:	val_out <= 16'h4f8b;
             14'hce0 	:	val_out <= 16'h4f91;
             14'hce1 	:	val_out <= 16'h4f97;
             14'hce2 	:	val_out <= 16'h4f9d;
             14'hce3 	:	val_out <= 16'h4fa3;
             14'hce4 	:	val_out <= 16'h4fa9;
             14'hce5 	:	val_out <= 16'h4faf;
             14'hce6 	:	val_out <= 16'h4fb5;
             14'hce7 	:	val_out <= 16'h4fbb;
             14'hce8 	:	val_out <= 16'h4fc1;
             14'hce9 	:	val_out <= 16'h4fc7;
             14'hcea 	:	val_out <= 16'h4fcd;
             14'hceb 	:	val_out <= 16'h4fd3;
             14'hcec 	:	val_out <= 16'h4fd9;
             14'hced 	:	val_out <= 16'h4fdf;
             14'hcee 	:	val_out <= 16'h4fe5;
             14'hcef 	:	val_out <= 16'h4fea;
             14'hcf0 	:	val_out <= 16'h4ff0;
             14'hcf1 	:	val_out <= 16'h4ff6;
             14'hcf2 	:	val_out <= 16'h4ffc;
             14'hcf3 	:	val_out <= 16'h5002;
             14'hcf4 	:	val_out <= 16'h5008;
             14'hcf5 	:	val_out <= 16'h500e;
             14'hcf6 	:	val_out <= 16'h5014;
             14'hcf7 	:	val_out <= 16'h501a;
             14'hcf8 	:	val_out <= 16'h5020;
             14'hcf9 	:	val_out <= 16'h5026;
             14'hcfa 	:	val_out <= 16'h502c;
             14'hcfb 	:	val_out <= 16'h5032;
             14'hcfc 	:	val_out <= 16'h5038;
             14'hcfd 	:	val_out <= 16'h503e;
             14'hcfe 	:	val_out <= 16'h5044;
             14'hcff 	:	val_out <= 16'h504a;
             14'hd00 	:	val_out <= 16'h5050;
             14'hd01 	:	val_out <= 16'h5056;
             14'hd02 	:	val_out <= 16'h505c;
             14'hd03 	:	val_out <= 16'h5062;
             14'hd04 	:	val_out <= 16'h5068;
             14'hd05 	:	val_out <= 16'h506e;
             14'hd06 	:	val_out <= 16'h5074;
             14'hd07 	:	val_out <= 16'h507a;
             14'hd08 	:	val_out <= 16'h5080;
             14'hd09 	:	val_out <= 16'h5086;
             14'hd0a 	:	val_out <= 16'h508c;
             14'hd0b 	:	val_out <= 16'h5092;
             14'hd0c 	:	val_out <= 16'h5098;
             14'hd0d 	:	val_out <= 16'h509d;
             14'hd0e 	:	val_out <= 16'h50a3;
             14'hd0f 	:	val_out <= 16'h50a9;
             14'hd10 	:	val_out <= 16'h50af;
             14'hd11 	:	val_out <= 16'h50b5;
             14'hd12 	:	val_out <= 16'h50bb;
             14'hd13 	:	val_out <= 16'h50c1;
             14'hd14 	:	val_out <= 16'h50c7;
             14'hd15 	:	val_out <= 16'h50cd;
             14'hd16 	:	val_out <= 16'h50d3;
             14'hd17 	:	val_out <= 16'h50d9;
             14'hd18 	:	val_out <= 16'h50df;
             14'hd19 	:	val_out <= 16'h50e5;
             14'hd1a 	:	val_out <= 16'h50eb;
             14'hd1b 	:	val_out <= 16'h50f1;
             14'hd1c 	:	val_out <= 16'h50f7;
             14'hd1d 	:	val_out <= 16'h50fd;
             14'hd1e 	:	val_out <= 16'h5103;
             14'hd1f 	:	val_out <= 16'h5109;
             14'hd20 	:	val_out <= 16'h510f;
             14'hd21 	:	val_out <= 16'h5115;
             14'hd22 	:	val_out <= 16'h511b;
             14'hd23 	:	val_out <= 16'h5121;
             14'hd24 	:	val_out <= 16'h5127;
             14'hd25 	:	val_out <= 16'h512d;
             14'hd26 	:	val_out <= 16'h5132;
             14'hd27 	:	val_out <= 16'h5138;
             14'hd28 	:	val_out <= 16'h513e;
             14'hd29 	:	val_out <= 16'h5144;
             14'hd2a 	:	val_out <= 16'h514a;
             14'hd2b 	:	val_out <= 16'h5150;
             14'hd2c 	:	val_out <= 16'h5156;
             14'hd2d 	:	val_out <= 16'h515c;
             14'hd2e 	:	val_out <= 16'h5162;
             14'hd2f 	:	val_out <= 16'h5168;
             14'hd30 	:	val_out <= 16'h516e;
             14'hd31 	:	val_out <= 16'h5174;
             14'hd32 	:	val_out <= 16'h517a;
             14'hd33 	:	val_out <= 16'h5180;
             14'hd34 	:	val_out <= 16'h5186;
             14'hd35 	:	val_out <= 16'h518c;
             14'hd36 	:	val_out <= 16'h5192;
             14'hd37 	:	val_out <= 16'h5198;
             14'hd38 	:	val_out <= 16'h519e;
             14'hd39 	:	val_out <= 16'h51a4;
             14'hd3a 	:	val_out <= 16'h51aa;
             14'hd3b 	:	val_out <= 16'h51b0;
             14'hd3c 	:	val_out <= 16'h51b6;
             14'hd3d 	:	val_out <= 16'h51bb;
             14'hd3e 	:	val_out <= 16'h51c1;
             14'hd3f 	:	val_out <= 16'h51c7;
             14'hd40 	:	val_out <= 16'h51cd;
             14'hd41 	:	val_out <= 16'h51d3;
             14'hd42 	:	val_out <= 16'h51d9;
             14'hd43 	:	val_out <= 16'h51df;
             14'hd44 	:	val_out <= 16'h51e5;
             14'hd45 	:	val_out <= 16'h51eb;
             14'hd46 	:	val_out <= 16'h51f1;
             14'hd47 	:	val_out <= 16'h51f7;
             14'hd48 	:	val_out <= 16'h51fd;
             14'hd49 	:	val_out <= 16'h5203;
             14'hd4a 	:	val_out <= 16'h5209;
             14'hd4b 	:	val_out <= 16'h520f;
             14'hd4c 	:	val_out <= 16'h5215;
             14'hd4d 	:	val_out <= 16'h521b;
             14'hd4e 	:	val_out <= 16'h5221;
             14'hd4f 	:	val_out <= 16'h5227;
             14'hd50 	:	val_out <= 16'h522d;
             14'hd51 	:	val_out <= 16'h5233;
             14'hd52 	:	val_out <= 16'h5238;
             14'hd53 	:	val_out <= 16'h523e;
             14'hd54 	:	val_out <= 16'h5244;
             14'hd55 	:	val_out <= 16'h524a;
             14'hd56 	:	val_out <= 16'h5250;
             14'hd57 	:	val_out <= 16'h5256;
             14'hd58 	:	val_out <= 16'h525c;
             14'hd59 	:	val_out <= 16'h5262;
             14'hd5a 	:	val_out <= 16'h5268;
             14'hd5b 	:	val_out <= 16'h526e;
             14'hd5c 	:	val_out <= 16'h5274;
             14'hd5d 	:	val_out <= 16'h527a;
             14'hd5e 	:	val_out <= 16'h5280;
             14'hd5f 	:	val_out <= 16'h5286;
             14'hd60 	:	val_out <= 16'h528c;
             14'hd61 	:	val_out <= 16'h5292;
             14'hd62 	:	val_out <= 16'h5298;
             14'hd63 	:	val_out <= 16'h529e;
             14'hd64 	:	val_out <= 16'h52a4;
             14'hd65 	:	val_out <= 16'h52aa;
             14'hd66 	:	val_out <= 16'h52af;
             14'hd67 	:	val_out <= 16'h52b5;
             14'hd68 	:	val_out <= 16'h52bb;
             14'hd69 	:	val_out <= 16'h52c1;
             14'hd6a 	:	val_out <= 16'h52c7;
             14'hd6b 	:	val_out <= 16'h52cd;
             14'hd6c 	:	val_out <= 16'h52d3;
             14'hd6d 	:	val_out <= 16'h52d9;
             14'hd6e 	:	val_out <= 16'h52df;
             14'hd6f 	:	val_out <= 16'h52e5;
             14'hd70 	:	val_out <= 16'h52eb;
             14'hd71 	:	val_out <= 16'h52f1;
             14'hd72 	:	val_out <= 16'h52f7;
             14'hd73 	:	val_out <= 16'h52fd;
             14'hd74 	:	val_out <= 16'h5303;
             14'hd75 	:	val_out <= 16'h5309;
             14'hd76 	:	val_out <= 16'h530f;
             14'hd77 	:	val_out <= 16'h5315;
             14'hd78 	:	val_out <= 16'h531a;
             14'hd79 	:	val_out <= 16'h5320;
             14'hd7a 	:	val_out <= 16'h5326;
             14'hd7b 	:	val_out <= 16'h532c;
             14'hd7c 	:	val_out <= 16'h5332;
             14'hd7d 	:	val_out <= 16'h5338;
             14'hd7e 	:	val_out <= 16'h533e;
             14'hd7f 	:	val_out <= 16'h5344;
             14'hd80 	:	val_out <= 16'h534a;
             14'hd81 	:	val_out <= 16'h5350;
             14'hd82 	:	val_out <= 16'h5356;
             14'hd83 	:	val_out <= 16'h535c;
             14'hd84 	:	val_out <= 16'h5362;
             14'hd85 	:	val_out <= 16'h5368;
             14'hd86 	:	val_out <= 16'h536e;
             14'hd87 	:	val_out <= 16'h5374;
             14'hd88 	:	val_out <= 16'h537a;
             14'hd89 	:	val_out <= 16'h537f;
             14'hd8a 	:	val_out <= 16'h5385;
             14'hd8b 	:	val_out <= 16'h538b;
             14'hd8c 	:	val_out <= 16'h5391;
             14'hd8d 	:	val_out <= 16'h5397;
             14'hd8e 	:	val_out <= 16'h539d;
             14'hd8f 	:	val_out <= 16'h53a3;
             14'hd90 	:	val_out <= 16'h53a9;
             14'hd91 	:	val_out <= 16'h53af;
             14'hd92 	:	val_out <= 16'h53b5;
             14'hd93 	:	val_out <= 16'h53bb;
             14'hd94 	:	val_out <= 16'h53c1;
             14'hd95 	:	val_out <= 16'h53c7;
             14'hd96 	:	val_out <= 16'h53cd;
             14'hd97 	:	val_out <= 16'h53d3;
             14'hd98 	:	val_out <= 16'h53d9;
             14'hd99 	:	val_out <= 16'h53de;
             14'hd9a 	:	val_out <= 16'h53e4;
             14'hd9b 	:	val_out <= 16'h53ea;
             14'hd9c 	:	val_out <= 16'h53f0;
             14'hd9d 	:	val_out <= 16'h53f6;
             14'hd9e 	:	val_out <= 16'h53fc;
             14'hd9f 	:	val_out <= 16'h5402;
             14'hda0 	:	val_out <= 16'h5408;
             14'hda1 	:	val_out <= 16'h540e;
             14'hda2 	:	val_out <= 16'h5414;
             14'hda3 	:	val_out <= 16'h541a;
             14'hda4 	:	val_out <= 16'h5420;
             14'hda5 	:	val_out <= 16'h5426;
             14'hda6 	:	val_out <= 16'h542c;
             14'hda7 	:	val_out <= 16'h5432;
             14'hda8 	:	val_out <= 16'h5438;
             14'hda9 	:	val_out <= 16'h543d;
             14'hdaa 	:	val_out <= 16'h5443;
             14'hdab 	:	val_out <= 16'h5449;
             14'hdac 	:	val_out <= 16'h544f;
             14'hdad 	:	val_out <= 16'h5455;
             14'hdae 	:	val_out <= 16'h545b;
             14'hdaf 	:	val_out <= 16'h5461;
             14'hdb0 	:	val_out <= 16'h5467;
             14'hdb1 	:	val_out <= 16'h546d;
             14'hdb2 	:	val_out <= 16'h5473;
             14'hdb3 	:	val_out <= 16'h5479;
             14'hdb4 	:	val_out <= 16'h547f;
             14'hdb5 	:	val_out <= 16'h5485;
             14'hdb6 	:	val_out <= 16'h548b;
             14'hdb7 	:	val_out <= 16'h5490;
             14'hdb8 	:	val_out <= 16'h5496;
             14'hdb9 	:	val_out <= 16'h549c;
             14'hdba 	:	val_out <= 16'h54a2;
             14'hdbb 	:	val_out <= 16'h54a8;
             14'hdbc 	:	val_out <= 16'h54ae;
             14'hdbd 	:	val_out <= 16'h54b4;
             14'hdbe 	:	val_out <= 16'h54ba;
             14'hdbf 	:	val_out <= 16'h54c0;
             14'hdc0 	:	val_out <= 16'h54c6;
             14'hdc1 	:	val_out <= 16'h54cc;
             14'hdc2 	:	val_out <= 16'h54d2;
             14'hdc3 	:	val_out <= 16'h54d8;
             14'hdc4 	:	val_out <= 16'h54de;
             14'hdc5 	:	val_out <= 16'h54e3;
             14'hdc6 	:	val_out <= 16'h54e9;
             14'hdc7 	:	val_out <= 16'h54ef;
             14'hdc8 	:	val_out <= 16'h54f5;
             14'hdc9 	:	val_out <= 16'h54fb;
             14'hdca 	:	val_out <= 16'h5501;
             14'hdcb 	:	val_out <= 16'h5507;
             14'hdcc 	:	val_out <= 16'h550d;
             14'hdcd 	:	val_out <= 16'h5513;
             14'hdce 	:	val_out <= 16'h5519;
             14'hdcf 	:	val_out <= 16'h551f;
             14'hdd0 	:	val_out <= 16'h5525;
             14'hdd1 	:	val_out <= 16'h552b;
             14'hdd2 	:	val_out <= 16'h5531;
             14'hdd3 	:	val_out <= 16'h5536;
             14'hdd4 	:	val_out <= 16'h553c;
             14'hdd5 	:	val_out <= 16'h5542;
             14'hdd6 	:	val_out <= 16'h5548;
             14'hdd7 	:	val_out <= 16'h554e;
             14'hdd8 	:	val_out <= 16'h5554;
             14'hdd9 	:	val_out <= 16'h555a;
             14'hdda 	:	val_out <= 16'h5560;
             14'hddb 	:	val_out <= 16'h5566;
             14'hddc 	:	val_out <= 16'h556c;
             14'hddd 	:	val_out <= 16'h5572;
             14'hdde 	:	val_out <= 16'h5578;
             14'hddf 	:	val_out <= 16'h557e;
             14'hde0 	:	val_out <= 16'h5583;
             14'hde1 	:	val_out <= 16'h5589;
             14'hde2 	:	val_out <= 16'h558f;
             14'hde3 	:	val_out <= 16'h5595;
             14'hde4 	:	val_out <= 16'h559b;
             14'hde5 	:	val_out <= 16'h55a1;
             14'hde6 	:	val_out <= 16'h55a7;
             14'hde7 	:	val_out <= 16'h55ad;
             14'hde8 	:	val_out <= 16'h55b3;
             14'hde9 	:	val_out <= 16'h55b9;
             14'hdea 	:	val_out <= 16'h55bf;
             14'hdeb 	:	val_out <= 16'h55c5;
             14'hdec 	:	val_out <= 16'h55cb;
             14'hded 	:	val_out <= 16'h55d0;
             14'hdee 	:	val_out <= 16'h55d6;
             14'hdef 	:	val_out <= 16'h55dc;
             14'hdf0 	:	val_out <= 16'h55e2;
             14'hdf1 	:	val_out <= 16'h55e8;
             14'hdf2 	:	val_out <= 16'h55ee;
             14'hdf3 	:	val_out <= 16'h55f4;
             14'hdf4 	:	val_out <= 16'h55fa;
             14'hdf5 	:	val_out <= 16'h5600;
             14'hdf6 	:	val_out <= 16'h5606;
             14'hdf7 	:	val_out <= 16'h560c;
             14'hdf8 	:	val_out <= 16'h5612;
             14'hdf9 	:	val_out <= 16'h5617;
             14'hdfa 	:	val_out <= 16'h561d;
             14'hdfb 	:	val_out <= 16'h5623;
             14'hdfc 	:	val_out <= 16'h5629;
             14'hdfd 	:	val_out <= 16'h562f;
             14'hdfe 	:	val_out <= 16'h5635;
             14'hdff 	:	val_out <= 16'h563b;
             14'he00 	:	val_out <= 16'h5641;
             14'he01 	:	val_out <= 16'h5647;
             14'he02 	:	val_out <= 16'h564d;
             14'he03 	:	val_out <= 16'h5653;
             14'he04 	:	val_out <= 16'h5659;
             14'he05 	:	val_out <= 16'h565e;
             14'he06 	:	val_out <= 16'h5664;
             14'he07 	:	val_out <= 16'h566a;
             14'he08 	:	val_out <= 16'h5670;
             14'he09 	:	val_out <= 16'h5676;
             14'he0a 	:	val_out <= 16'h567c;
             14'he0b 	:	val_out <= 16'h5682;
             14'he0c 	:	val_out <= 16'h5688;
             14'he0d 	:	val_out <= 16'h568e;
             14'he0e 	:	val_out <= 16'h5694;
             14'he0f 	:	val_out <= 16'h569a;
             14'he10 	:	val_out <= 16'h569f;
             14'he11 	:	val_out <= 16'h56a5;
             14'he12 	:	val_out <= 16'h56ab;
             14'he13 	:	val_out <= 16'h56b1;
             14'he14 	:	val_out <= 16'h56b7;
             14'he15 	:	val_out <= 16'h56bd;
             14'he16 	:	val_out <= 16'h56c3;
             14'he17 	:	val_out <= 16'h56c9;
             14'he18 	:	val_out <= 16'h56cf;
             14'he19 	:	val_out <= 16'h56d5;
             14'he1a 	:	val_out <= 16'h56db;
             14'he1b 	:	val_out <= 16'h56e1;
             14'he1c 	:	val_out <= 16'h56e6;
             14'he1d 	:	val_out <= 16'h56ec;
             14'he1e 	:	val_out <= 16'h56f2;
             14'he1f 	:	val_out <= 16'h56f8;
             14'he20 	:	val_out <= 16'h56fe;
             14'he21 	:	val_out <= 16'h5704;
             14'he22 	:	val_out <= 16'h570a;
             14'he23 	:	val_out <= 16'h5710;
             14'he24 	:	val_out <= 16'h5716;
             14'he25 	:	val_out <= 16'h571c;
             14'he26 	:	val_out <= 16'h5722;
             14'he27 	:	val_out <= 16'h5727;
             14'he28 	:	val_out <= 16'h572d;
             14'he29 	:	val_out <= 16'h5733;
             14'he2a 	:	val_out <= 16'h5739;
             14'he2b 	:	val_out <= 16'h573f;
             14'he2c 	:	val_out <= 16'h5745;
             14'he2d 	:	val_out <= 16'h574b;
             14'he2e 	:	val_out <= 16'h5751;
             14'he2f 	:	val_out <= 16'h5757;
             14'he30 	:	val_out <= 16'h575d;
             14'he31 	:	val_out <= 16'h5763;
             14'he32 	:	val_out <= 16'h5768;
             14'he33 	:	val_out <= 16'h576e;
             14'he34 	:	val_out <= 16'h5774;
             14'he35 	:	val_out <= 16'h577a;
             14'he36 	:	val_out <= 16'h5780;
             14'he37 	:	val_out <= 16'h5786;
             14'he38 	:	val_out <= 16'h578c;
             14'he39 	:	val_out <= 16'h5792;
             14'he3a 	:	val_out <= 16'h5798;
             14'he3b 	:	val_out <= 16'h579e;
             14'he3c 	:	val_out <= 16'h57a3;
             14'he3d 	:	val_out <= 16'h57a9;
             14'he3e 	:	val_out <= 16'h57af;
             14'he3f 	:	val_out <= 16'h57b5;
             14'he40 	:	val_out <= 16'h57bb;
             14'he41 	:	val_out <= 16'h57c1;
             14'he42 	:	val_out <= 16'h57c7;
             14'he43 	:	val_out <= 16'h57cd;
             14'he44 	:	val_out <= 16'h57d3;
             14'he45 	:	val_out <= 16'h57d9;
             14'he46 	:	val_out <= 16'h57de;
             14'he47 	:	val_out <= 16'h57e4;
             14'he48 	:	val_out <= 16'h57ea;
             14'he49 	:	val_out <= 16'h57f0;
             14'he4a 	:	val_out <= 16'h57f6;
             14'he4b 	:	val_out <= 16'h57fc;
             14'he4c 	:	val_out <= 16'h5802;
             14'he4d 	:	val_out <= 16'h5808;
             14'he4e 	:	val_out <= 16'h580e;
             14'he4f 	:	val_out <= 16'h5814;
             14'he50 	:	val_out <= 16'h5819;
             14'he51 	:	val_out <= 16'h581f;
             14'he52 	:	val_out <= 16'h5825;
             14'he53 	:	val_out <= 16'h582b;
             14'he54 	:	val_out <= 16'h5831;
             14'he55 	:	val_out <= 16'h5837;
             14'he56 	:	val_out <= 16'h583d;
             14'he57 	:	val_out <= 16'h5843;
             14'he58 	:	val_out <= 16'h5849;
             14'he59 	:	val_out <= 16'h584f;
             14'he5a 	:	val_out <= 16'h5854;
             14'he5b 	:	val_out <= 16'h585a;
             14'he5c 	:	val_out <= 16'h5860;
             14'he5d 	:	val_out <= 16'h5866;
             14'he5e 	:	val_out <= 16'h586c;
             14'he5f 	:	val_out <= 16'h5872;
             14'he60 	:	val_out <= 16'h5878;
             14'he61 	:	val_out <= 16'h587e;
             14'he62 	:	val_out <= 16'h5884;
             14'he63 	:	val_out <= 16'h588a;
             14'he64 	:	val_out <= 16'h588f;
             14'he65 	:	val_out <= 16'h5895;
             14'he66 	:	val_out <= 16'h589b;
             14'he67 	:	val_out <= 16'h58a1;
             14'he68 	:	val_out <= 16'h58a7;
             14'he69 	:	val_out <= 16'h58ad;
             14'he6a 	:	val_out <= 16'h58b3;
             14'he6b 	:	val_out <= 16'h58b9;
             14'he6c 	:	val_out <= 16'h58bf;
             14'he6d 	:	val_out <= 16'h58c4;
             14'he6e 	:	val_out <= 16'h58ca;
             14'he6f 	:	val_out <= 16'h58d0;
             14'he70 	:	val_out <= 16'h58d6;
             14'he71 	:	val_out <= 16'h58dc;
             14'he72 	:	val_out <= 16'h58e2;
             14'he73 	:	val_out <= 16'h58e8;
             14'he74 	:	val_out <= 16'h58ee;
             14'he75 	:	val_out <= 16'h58f4;
             14'he76 	:	val_out <= 16'h58fa;
             14'he77 	:	val_out <= 16'h58ff;
             14'he78 	:	val_out <= 16'h5905;
             14'he79 	:	val_out <= 16'h590b;
             14'he7a 	:	val_out <= 16'h5911;
             14'he7b 	:	val_out <= 16'h5917;
             14'he7c 	:	val_out <= 16'h591d;
             14'he7d 	:	val_out <= 16'h5923;
             14'he7e 	:	val_out <= 16'h5929;
             14'he7f 	:	val_out <= 16'h592f;
             14'he80 	:	val_out <= 16'h5934;
             14'he81 	:	val_out <= 16'h593a;
             14'he82 	:	val_out <= 16'h5940;
             14'he83 	:	val_out <= 16'h5946;
             14'he84 	:	val_out <= 16'h594c;
             14'he85 	:	val_out <= 16'h5952;
             14'he86 	:	val_out <= 16'h5958;
             14'he87 	:	val_out <= 16'h595e;
             14'he88 	:	val_out <= 16'h5964;
             14'he89 	:	val_out <= 16'h5969;
             14'he8a 	:	val_out <= 16'h596f;
             14'he8b 	:	val_out <= 16'h5975;
             14'he8c 	:	val_out <= 16'h597b;
             14'he8d 	:	val_out <= 16'h5981;
             14'he8e 	:	val_out <= 16'h5987;
             14'he8f 	:	val_out <= 16'h598d;
             14'he90 	:	val_out <= 16'h5993;
             14'he91 	:	val_out <= 16'h5999;
             14'he92 	:	val_out <= 16'h599e;
             14'he93 	:	val_out <= 16'h59a4;
             14'he94 	:	val_out <= 16'h59aa;
             14'he95 	:	val_out <= 16'h59b0;
             14'he96 	:	val_out <= 16'h59b6;
             14'he97 	:	val_out <= 16'h59bc;
             14'he98 	:	val_out <= 16'h59c2;
             14'he99 	:	val_out <= 16'h59c8;
             14'he9a 	:	val_out <= 16'h59cd;
             14'he9b 	:	val_out <= 16'h59d3;
             14'he9c 	:	val_out <= 16'h59d9;
             14'he9d 	:	val_out <= 16'h59df;
             14'he9e 	:	val_out <= 16'h59e5;
             14'he9f 	:	val_out <= 16'h59eb;
             14'hea0 	:	val_out <= 16'h59f1;
             14'hea1 	:	val_out <= 16'h59f7;
             14'hea2 	:	val_out <= 16'h59fd;
             14'hea3 	:	val_out <= 16'h5a02;
             14'hea4 	:	val_out <= 16'h5a08;
             14'hea5 	:	val_out <= 16'h5a0e;
             14'hea6 	:	val_out <= 16'h5a14;
             14'hea7 	:	val_out <= 16'h5a1a;
             14'hea8 	:	val_out <= 16'h5a20;
             14'hea9 	:	val_out <= 16'h5a26;
             14'heaa 	:	val_out <= 16'h5a2c;
             14'heab 	:	val_out <= 16'h5a31;
             14'heac 	:	val_out <= 16'h5a37;
             14'head 	:	val_out <= 16'h5a3d;
             14'heae 	:	val_out <= 16'h5a43;
             14'heaf 	:	val_out <= 16'h5a49;
             14'heb0 	:	val_out <= 16'h5a4f;
             14'heb1 	:	val_out <= 16'h5a55;
             14'heb2 	:	val_out <= 16'h5a5b;
             14'heb3 	:	val_out <= 16'h5a60;
             14'heb4 	:	val_out <= 16'h5a66;
             14'heb5 	:	val_out <= 16'h5a6c;
             14'heb6 	:	val_out <= 16'h5a72;
             14'heb7 	:	val_out <= 16'h5a78;
             14'heb8 	:	val_out <= 16'h5a7e;
             14'heb9 	:	val_out <= 16'h5a84;
             14'heba 	:	val_out <= 16'h5a8a;
             14'hebb 	:	val_out <= 16'h5a90;
             14'hebc 	:	val_out <= 16'h5a95;
             14'hebd 	:	val_out <= 16'h5a9b;
             14'hebe 	:	val_out <= 16'h5aa1;
             14'hebf 	:	val_out <= 16'h5aa7;
             14'hec0 	:	val_out <= 16'h5aad;
             14'hec1 	:	val_out <= 16'h5ab3;
             14'hec2 	:	val_out <= 16'h5ab9;
             14'hec3 	:	val_out <= 16'h5abf;
             14'hec4 	:	val_out <= 16'h5ac4;
             14'hec5 	:	val_out <= 16'h5aca;
             14'hec6 	:	val_out <= 16'h5ad0;
             14'hec7 	:	val_out <= 16'h5ad6;
             14'hec8 	:	val_out <= 16'h5adc;
             14'hec9 	:	val_out <= 16'h5ae2;
             14'heca 	:	val_out <= 16'h5ae8;
             14'hecb 	:	val_out <= 16'h5aee;
             14'hecc 	:	val_out <= 16'h5af3;
             14'hecd 	:	val_out <= 16'h5af9;
             14'hece 	:	val_out <= 16'h5aff;
             14'hecf 	:	val_out <= 16'h5b05;
             14'hed0 	:	val_out <= 16'h5b0b;
             14'hed1 	:	val_out <= 16'h5b11;
             14'hed2 	:	val_out <= 16'h5b17;
             14'hed3 	:	val_out <= 16'h5b1d;
             14'hed4 	:	val_out <= 16'h5b22;
             14'hed5 	:	val_out <= 16'h5b28;
             14'hed6 	:	val_out <= 16'h5b2e;
             14'hed7 	:	val_out <= 16'h5b34;
             14'hed8 	:	val_out <= 16'h5b3a;
             14'hed9 	:	val_out <= 16'h5b40;
             14'heda 	:	val_out <= 16'h5b46;
             14'hedb 	:	val_out <= 16'h5b4b;
             14'hedc 	:	val_out <= 16'h5b51;
             14'hedd 	:	val_out <= 16'h5b57;
             14'hede 	:	val_out <= 16'h5b5d;
             14'hedf 	:	val_out <= 16'h5b63;
             14'hee0 	:	val_out <= 16'h5b69;
             14'hee1 	:	val_out <= 16'h5b6f;
             14'hee2 	:	val_out <= 16'h5b75;
             14'hee3 	:	val_out <= 16'h5b7a;
             14'hee4 	:	val_out <= 16'h5b80;
             14'hee5 	:	val_out <= 16'h5b86;
             14'hee6 	:	val_out <= 16'h5b8c;
             14'hee7 	:	val_out <= 16'h5b92;
             14'hee8 	:	val_out <= 16'h5b98;
             14'hee9 	:	val_out <= 16'h5b9e;
             14'heea 	:	val_out <= 16'h5ba3;
             14'heeb 	:	val_out <= 16'h5ba9;
             14'heec 	:	val_out <= 16'h5baf;
             14'heed 	:	val_out <= 16'h5bb5;
             14'heee 	:	val_out <= 16'h5bbb;
             14'heef 	:	val_out <= 16'h5bc1;
             14'hef0 	:	val_out <= 16'h5bc7;
             14'hef1 	:	val_out <= 16'h5bcd;
             14'hef2 	:	val_out <= 16'h5bd2;
             14'hef3 	:	val_out <= 16'h5bd8;
             14'hef4 	:	val_out <= 16'h5bde;
             14'hef5 	:	val_out <= 16'h5be4;
             14'hef6 	:	val_out <= 16'h5bea;
             14'hef7 	:	val_out <= 16'h5bf0;
             14'hef8 	:	val_out <= 16'h5bf6;
             14'hef9 	:	val_out <= 16'h5bfb;
             14'hefa 	:	val_out <= 16'h5c01;
             14'hefb 	:	val_out <= 16'h5c07;
             14'hefc 	:	val_out <= 16'h5c0d;
             14'hefd 	:	val_out <= 16'h5c13;
             14'hefe 	:	val_out <= 16'h5c19;
             14'heff 	:	val_out <= 16'h5c1f;
             14'hf00 	:	val_out <= 16'h5c25;
             14'hf01 	:	val_out <= 16'h5c2a;
             14'hf02 	:	val_out <= 16'h5c30;
             14'hf03 	:	val_out <= 16'h5c36;
             14'hf04 	:	val_out <= 16'h5c3c;
             14'hf05 	:	val_out <= 16'h5c42;
             14'hf06 	:	val_out <= 16'h5c48;
             14'hf07 	:	val_out <= 16'h5c4e;
             14'hf08 	:	val_out <= 16'h5c53;
             14'hf09 	:	val_out <= 16'h5c59;
             14'hf0a 	:	val_out <= 16'h5c5f;
             14'hf0b 	:	val_out <= 16'h5c65;
             14'hf0c 	:	val_out <= 16'h5c6b;
             14'hf0d 	:	val_out <= 16'h5c71;
             14'hf0e 	:	val_out <= 16'h5c77;
             14'hf0f 	:	val_out <= 16'h5c7c;
             14'hf10 	:	val_out <= 16'h5c82;
             14'hf11 	:	val_out <= 16'h5c88;
             14'hf12 	:	val_out <= 16'h5c8e;
             14'hf13 	:	val_out <= 16'h5c94;
             14'hf14 	:	val_out <= 16'h5c9a;
             14'hf15 	:	val_out <= 16'h5ca0;
             14'hf16 	:	val_out <= 16'h5ca5;
             14'hf17 	:	val_out <= 16'h5cab;
             14'hf18 	:	val_out <= 16'h5cb1;
             14'hf19 	:	val_out <= 16'h5cb7;
             14'hf1a 	:	val_out <= 16'h5cbd;
             14'hf1b 	:	val_out <= 16'h5cc3;
             14'hf1c 	:	val_out <= 16'h5cc9;
             14'hf1d 	:	val_out <= 16'h5cce;
             14'hf1e 	:	val_out <= 16'h5cd4;
             14'hf1f 	:	val_out <= 16'h5cda;
             14'hf20 	:	val_out <= 16'h5ce0;
             14'hf21 	:	val_out <= 16'h5ce6;
             14'hf22 	:	val_out <= 16'h5cec;
             14'hf23 	:	val_out <= 16'h5cf2;
             14'hf24 	:	val_out <= 16'h5cf7;
             14'hf25 	:	val_out <= 16'h5cfd;
             14'hf26 	:	val_out <= 16'h5d03;
             14'hf27 	:	val_out <= 16'h5d09;
             14'hf28 	:	val_out <= 16'h5d0f;
             14'hf29 	:	val_out <= 16'h5d15;
             14'hf2a 	:	val_out <= 16'h5d1b;
             14'hf2b 	:	val_out <= 16'h5d20;
             14'hf2c 	:	val_out <= 16'h5d26;
             14'hf2d 	:	val_out <= 16'h5d2c;
             14'hf2e 	:	val_out <= 16'h5d32;
             14'hf2f 	:	val_out <= 16'h5d38;
             14'hf30 	:	val_out <= 16'h5d3e;
             14'hf31 	:	val_out <= 16'h5d43;
             14'hf32 	:	val_out <= 16'h5d49;
             14'hf33 	:	val_out <= 16'h5d4f;
             14'hf34 	:	val_out <= 16'h5d55;
             14'hf35 	:	val_out <= 16'h5d5b;
             14'hf36 	:	val_out <= 16'h5d61;
             14'hf37 	:	val_out <= 16'h5d67;
             14'hf38 	:	val_out <= 16'h5d6c;
             14'hf39 	:	val_out <= 16'h5d72;
             14'hf3a 	:	val_out <= 16'h5d78;
             14'hf3b 	:	val_out <= 16'h5d7e;
             14'hf3c 	:	val_out <= 16'h5d84;
             14'hf3d 	:	val_out <= 16'h5d8a;
             14'hf3e 	:	val_out <= 16'h5d90;
             14'hf3f 	:	val_out <= 16'h5d95;
             14'hf40 	:	val_out <= 16'h5d9b;
             14'hf41 	:	val_out <= 16'h5da1;
             14'hf42 	:	val_out <= 16'h5da7;
             14'hf43 	:	val_out <= 16'h5dad;
             14'hf44 	:	val_out <= 16'h5db3;
             14'hf45 	:	val_out <= 16'h5db8;
             14'hf46 	:	val_out <= 16'h5dbe;
             14'hf47 	:	val_out <= 16'h5dc4;
             14'hf48 	:	val_out <= 16'h5dca;
             14'hf49 	:	val_out <= 16'h5dd0;
             14'hf4a 	:	val_out <= 16'h5dd6;
             14'hf4b 	:	val_out <= 16'h5ddc;
             14'hf4c 	:	val_out <= 16'h5de1;
             14'hf4d 	:	val_out <= 16'h5de7;
             14'hf4e 	:	val_out <= 16'h5ded;
             14'hf4f 	:	val_out <= 16'h5df3;
             14'hf50 	:	val_out <= 16'h5df9;
             14'hf51 	:	val_out <= 16'h5dff;
             14'hf52 	:	val_out <= 16'h5e04;
             14'hf53 	:	val_out <= 16'h5e0a;
             14'hf54 	:	val_out <= 16'h5e10;
             14'hf55 	:	val_out <= 16'h5e16;
             14'hf56 	:	val_out <= 16'h5e1c;
             14'hf57 	:	val_out <= 16'h5e22;
             14'hf58 	:	val_out <= 16'h5e28;
             14'hf59 	:	val_out <= 16'h5e2d;
             14'hf5a 	:	val_out <= 16'h5e33;
             14'hf5b 	:	val_out <= 16'h5e39;
             14'hf5c 	:	val_out <= 16'h5e3f;
             14'hf5d 	:	val_out <= 16'h5e45;
             14'hf5e 	:	val_out <= 16'h5e4b;
             14'hf5f 	:	val_out <= 16'h5e50;
             14'hf60 	:	val_out <= 16'h5e56;
             14'hf61 	:	val_out <= 16'h5e5c;
             14'hf62 	:	val_out <= 16'h5e62;
             14'hf63 	:	val_out <= 16'h5e68;
             14'hf64 	:	val_out <= 16'h5e6e;
             14'hf65 	:	val_out <= 16'h5e73;
             14'hf66 	:	val_out <= 16'h5e79;
             14'hf67 	:	val_out <= 16'h5e7f;
             14'hf68 	:	val_out <= 16'h5e85;
             14'hf69 	:	val_out <= 16'h5e8b;
             14'hf6a 	:	val_out <= 16'h5e91;
             14'hf6b 	:	val_out <= 16'h5e97;
             14'hf6c 	:	val_out <= 16'h5e9c;
             14'hf6d 	:	val_out <= 16'h5ea2;
             14'hf6e 	:	val_out <= 16'h5ea8;
             14'hf6f 	:	val_out <= 16'h5eae;
             14'hf70 	:	val_out <= 16'h5eb4;
             14'hf71 	:	val_out <= 16'h5eba;
             14'hf72 	:	val_out <= 16'h5ebf;
             14'hf73 	:	val_out <= 16'h5ec5;
             14'hf74 	:	val_out <= 16'h5ecb;
             14'hf75 	:	val_out <= 16'h5ed1;
             14'hf76 	:	val_out <= 16'h5ed7;
             14'hf77 	:	val_out <= 16'h5edd;
             14'hf78 	:	val_out <= 16'h5ee2;
             14'hf79 	:	val_out <= 16'h5ee8;
             14'hf7a 	:	val_out <= 16'h5eee;
             14'hf7b 	:	val_out <= 16'h5ef4;
             14'hf7c 	:	val_out <= 16'h5efa;
             14'hf7d 	:	val_out <= 16'h5f00;
             14'hf7e 	:	val_out <= 16'h5f05;
             14'hf7f 	:	val_out <= 16'h5f0b;
             14'hf80 	:	val_out <= 16'h5f11;
             14'hf81 	:	val_out <= 16'h5f17;
             14'hf82 	:	val_out <= 16'h5f1d;
             14'hf83 	:	val_out <= 16'h5f23;
             14'hf84 	:	val_out <= 16'h5f28;
             14'hf85 	:	val_out <= 16'h5f2e;
             14'hf86 	:	val_out <= 16'h5f34;
             14'hf87 	:	val_out <= 16'h5f3a;
             14'hf88 	:	val_out <= 16'h5f40;
             14'hf89 	:	val_out <= 16'h5f46;
             14'hf8a 	:	val_out <= 16'h5f4b;
             14'hf8b 	:	val_out <= 16'h5f51;
             14'hf8c 	:	val_out <= 16'h5f57;
             14'hf8d 	:	val_out <= 16'h5f5d;
             14'hf8e 	:	val_out <= 16'h5f63;
             14'hf8f 	:	val_out <= 16'h5f69;
             14'hf90 	:	val_out <= 16'h5f6e;
             14'hf91 	:	val_out <= 16'h5f74;
             14'hf92 	:	val_out <= 16'h5f7a;
             14'hf93 	:	val_out <= 16'h5f80;
             14'hf94 	:	val_out <= 16'h5f86;
             14'hf95 	:	val_out <= 16'h5f8c;
             14'hf96 	:	val_out <= 16'h5f91;
             14'hf97 	:	val_out <= 16'h5f97;
             14'hf98 	:	val_out <= 16'h5f9d;
             14'hf99 	:	val_out <= 16'h5fa3;
             14'hf9a 	:	val_out <= 16'h5fa9;
             14'hf9b 	:	val_out <= 16'h5fae;
             14'hf9c 	:	val_out <= 16'h5fb4;
             14'hf9d 	:	val_out <= 16'h5fba;
             14'hf9e 	:	val_out <= 16'h5fc0;
             14'hf9f 	:	val_out <= 16'h5fc6;
             14'hfa0 	:	val_out <= 16'h5fcc;
             14'hfa1 	:	val_out <= 16'h5fd1;
             14'hfa2 	:	val_out <= 16'h5fd7;
             14'hfa3 	:	val_out <= 16'h5fdd;
             14'hfa4 	:	val_out <= 16'h5fe3;
             14'hfa5 	:	val_out <= 16'h5fe9;
             14'hfa6 	:	val_out <= 16'h5fef;
             14'hfa7 	:	val_out <= 16'h5ff4;
             14'hfa8 	:	val_out <= 16'h5ffa;
             14'hfa9 	:	val_out <= 16'h6000;
             14'hfaa 	:	val_out <= 16'h6006;
             14'hfab 	:	val_out <= 16'h600c;
             14'hfac 	:	val_out <= 16'h6012;
             14'hfad 	:	val_out <= 16'h6017;
             14'hfae 	:	val_out <= 16'h601d;
             14'hfaf 	:	val_out <= 16'h6023;
             14'hfb0 	:	val_out <= 16'h6029;
             14'hfb1 	:	val_out <= 16'h602f;
             14'hfb2 	:	val_out <= 16'h6034;
             14'hfb3 	:	val_out <= 16'h603a;
             14'hfb4 	:	val_out <= 16'h6040;
             14'hfb5 	:	val_out <= 16'h6046;
             14'hfb6 	:	val_out <= 16'h604c;
             14'hfb7 	:	val_out <= 16'h6052;
             14'hfb8 	:	val_out <= 16'h6057;
             14'hfb9 	:	val_out <= 16'h605d;
             14'hfba 	:	val_out <= 16'h6063;
             14'hfbb 	:	val_out <= 16'h6069;
             14'hfbc 	:	val_out <= 16'h606f;
             14'hfbd 	:	val_out <= 16'h6075;
             14'hfbe 	:	val_out <= 16'h607a;
             14'hfbf 	:	val_out <= 16'h6080;
             14'hfc0 	:	val_out <= 16'h6086;
             14'hfc1 	:	val_out <= 16'h608c;
             14'hfc2 	:	val_out <= 16'h6092;
             14'hfc3 	:	val_out <= 16'h6097;
             14'hfc4 	:	val_out <= 16'h609d;
             14'hfc5 	:	val_out <= 16'h60a3;
             14'hfc6 	:	val_out <= 16'h60a9;
             14'hfc7 	:	val_out <= 16'h60af;
             14'hfc8 	:	val_out <= 16'h60b5;
             14'hfc9 	:	val_out <= 16'h60ba;
             14'hfca 	:	val_out <= 16'h60c0;
             14'hfcb 	:	val_out <= 16'h60c6;
             14'hfcc 	:	val_out <= 16'h60cc;
             14'hfcd 	:	val_out <= 16'h60d2;
             14'hfce 	:	val_out <= 16'h60d7;
             14'hfcf 	:	val_out <= 16'h60dd;
             14'hfd0 	:	val_out <= 16'h60e3;
             14'hfd1 	:	val_out <= 16'h60e9;
             14'hfd2 	:	val_out <= 16'h60ef;
             14'hfd3 	:	val_out <= 16'h60f4;
             14'hfd4 	:	val_out <= 16'h60fa;
             14'hfd5 	:	val_out <= 16'h6100;
             14'hfd6 	:	val_out <= 16'h6106;
             14'hfd7 	:	val_out <= 16'h610c;
             14'hfd8 	:	val_out <= 16'h6112;
             14'hfd9 	:	val_out <= 16'h6117;
             14'hfda 	:	val_out <= 16'h611d;
             14'hfdb 	:	val_out <= 16'h6123;
             14'hfdc 	:	val_out <= 16'h6129;
             14'hfdd 	:	val_out <= 16'h612f;
             14'hfde 	:	val_out <= 16'h6134;
             14'hfdf 	:	val_out <= 16'h613a;
             14'hfe0 	:	val_out <= 16'h6140;
             14'hfe1 	:	val_out <= 16'h6146;
             14'hfe2 	:	val_out <= 16'h614c;
             14'hfe3 	:	val_out <= 16'h6152;
             14'hfe4 	:	val_out <= 16'h6157;
             14'hfe5 	:	val_out <= 16'h615d;
             14'hfe6 	:	val_out <= 16'h6163;
             14'hfe7 	:	val_out <= 16'h6169;
             14'hfe8 	:	val_out <= 16'h616f;
             14'hfe9 	:	val_out <= 16'h6174;
             14'hfea 	:	val_out <= 16'h617a;
             14'hfeb 	:	val_out <= 16'h6180;
             14'hfec 	:	val_out <= 16'h6186;
             14'hfed 	:	val_out <= 16'h618c;
             14'hfee 	:	val_out <= 16'h6191;
             14'hfef 	:	val_out <= 16'h6197;
             14'hff0 	:	val_out <= 16'h619d;
             14'hff1 	:	val_out <= 16'h61a3;
             14'hff2 	:	val_out <= 16'h61a9;
             14'hff3 	:	val_out <= 16'h61ae;
             14'hff4 	:	val_out <= 16'h61b4;
             14'hff5 	:	val_out <= 16'h61ba;
             14'hff6 	:	val_out <= 16'h61c0;
             14'hff7 	:	val_out <= 16'h61c6;
             14'hff8 	:	val_out <= 16'h61cb;
             14'hff9 	:	val_out <= 16'h61d1;
             14'hffa 	:	val_out <= 16'h61d7;
             14'hffb 	:	val_out <= 16'h61dd;
             14'hffc 	:	val_out <= 16'h61e3;
             14'hffd 	:	val_out <= 16'h61e9;
             14'hffe 	:	val_out <= 16'h61ee;
             14'hfff 	:	val_out <= 16'h61f4;
             14'h1000 	:	val_out <= 16'h61fa;
             14'h1001 	:	val_out <= 16'h6200;
             14'h1002 	:	val_out <= 16'h6206;
             14'h1003 	:	val_out <= 16'h620b;
             14'h1004 	:	val_out <= 16'h6211;
             14'h1005 	:	val_out <= 16'h6217;
             14'h1006 	:	val_out <= 16'h621d;
             14'h1007 	:	val_out <= 16'h6223;
             14'h1008 	:	val_out <= 16'h6228;
             14'h1009 	:	val_out <= 16'h622e;
             14'h100a 	:	val_out <= 16'h6234;
             14'h100b 	:	val_out <= 16'h623a;
             14'h100c 	:	val_out <= 16'h6240;
             14'h100d 	:	val_out <= 16'h6245;
             14'h100e 	:	val_out <= 16'h624b;
             14'h100f 	:	val_out <= 16'h6251;
             14'h1010 	:	val_out <= 16'h6257;
             14'h1011 	:	val_out <= 16'h625d;
             14'h1012 	:	val_out <= 16'h6262;
             14'h1013 	:	val_out <= 16'h6268;
             14'h1014 	:	val_out <= 16'h626e;
             14'h1015 	:	val_out <= 16'h6274;
             14'h1016 	:	val_out <= 16'h627a;
             14'h1017 	:	val_out <= 16'h627f;
             14'h1018 	:	val_out <= 16'h6285;
             14'h1019 	:	val_out <= 16'h628b;
             14'h101a 	:	val_out <= 16'h6291;
             14'h101b 	:	val_out <= 16'h6297;
             14'h101c 	:	val_out <= 16'h629c;
             14'h101d 	:	val_out <= 16'h62a2;
             14'h101e 	:	val_out <= 16'h62a8;
             14'h101f 	:	val_out <= 16'h62ae;
             14'h1020 	:	val_out <= 16'h62b4;
             14'h1021 	:	val_out <= 16'h62b9;
             14'h1022 	:	val_out <= 16'h62bf;
             14'h1023 	:	val_out <= 16'h62c5;
             14'h1024 	:	val_out <= 16'h62cb;
             14'h1025 	:	val_out <= 16'h62d1;
             14'h1026 	:	val_out <= 16'h62d6;
             14'h1027 	:	val_out <= 16'h62dc;
             14'h1028 	:	val_out <= 16'h62e2;
             14'h1029 	:	val_out <= 16'h62e8;
             14'h102a 	:	val_out <= 16'h62ee;
             14'h102b 	:	val_out <= 16'h62f3;
             14'h102c 	:	val_out <= 16'h62f9;
             14'h102d 	:	val_out <= 16'h62ff;
             14'h102e 	:	val_out <= 16'h6305;
             14'h102f 	:	val_out <= 16'h630b;
             14'h1030 	:	val_out <= 16'h6310;
             14'h1031 	:	val_out <= 16'h6316;
             14'h1032 	:	val_out <= 16'h631c;
             14'h1033 	:	val_out <= 16'h6322;
             14'h1034 	:	val_out <= 16'h6327;
             14'h1035 	:	val_out <= 16'h632d;
             14'h1036 	:	val_out <= 16'h6333;
             14'h1037 	:	val_out <= 16'h6339;
             14'h1038 	:	val_out <= 16'h633f;
             14'h1039 	:	val_out <= 16'h6344;
             14'h103a 	:	val_out <= 16'h634a;
             14'h103b 	:	val_out <= 16'h6350;
             14'h103c 	:	val_out <= 16'h6356;
             14'h103d 	:	val_out <= 16'h635c;
             14'h103e 	:	val_out <= 16'h6361;
             14'h103f 	:	val_out <= 16'h6367;
             14'h1040 	:	val_out <= 16'h636d;
             14'h1041 	:	val_out <= 16'h6373;
             14'h1042 	:	val_out <= 16'h6379;
             14'h1043 	:	val_out <= 16'h637e;
             14'h1044 	:	val_out <= 16'h6384;
             14'h1045 	:	val_out <= 16'h638a;
             14'h1046 	:	val_out <= 16'h6390;
             14'h1047 	:	val_out <= 16'h6395;
             14'h1048 	:	val_out <= 16'h639b;
             14'h1049 	:	val_out <= 16'h63a1;
             14'h104a 	:	val_out <= 16'h63a7;
             14'h104b 	:	val_out <= 16'h63ad;
             14'h104c 	:	val_out <= 16'h63b2;
             14'h104d 	:	val_out <= 16'h63b8;
             14'h104e 	:	val_out <= 16'h63be;
             14'h104f 	:	val_out <= 16'h63c4;
             14'h1050 	:	val_out <= 16'h63ca;
             14'h1051 	:	val_out <= 16'h63cf;
             14'h1052 	:	val_out <= 16'h63d5;
             14'h1053 	:	val_out <= 16'h63db;
             14'h1054 	:	val_out <= 16'h63e1;
             14'h1055 	:	val_out <= 16'h63e7;
             14'h1056 	:	val_out <= 16'h63ec;
             14'h1057 	:	val_out <= 16'h63f2;
             14'h1058 	:	val_out <= 16'h63f8;
             14'h1059 	:	val_out <= 16'h63fe;
             14'h105a 	:	val_out <= 16'h6403;
             14'h105b 	:	val_out <= 16'h6409;
             14'h105c 	:	val_out <= 16'h640f;
             14'h105d 	:	val_out <= 16'h6415;
             14'h105e 	:	val_out <= 16'h641b;
             14'h105f 	:	val_out <= 16'h6420;
             14'h1060 	:	val_out <= 16'h6426;
             14'h1061 	:	val_out <= 16'h642c;
             14'h1062 	:	val_out <= 16'h6432;
             14'h1063 	:	val_out <= 16'h6437;
             14'h1064 	:	val_out <= 16'h643d;
             14'h1065 	:	val_out <= 16'h6443;
             14'h1066 	:	val_out <= 16'h6449;
             14'h1067 	:	val_out <= 16'h644f;
             14'h1068 	:	val_out <= 16'h6454;
             14'h1069 	:	val_out <= 16'h645a;
             14'h106a 	:	val_out <= 16'h6460;
             14'h106b 	:	val_out <= 16'h6466;
             14'h106c 	:	val_out <= 16'h646c;
             14'h106d 	:	val_out <= 16'h6471;
             14'h106e 	:	val_out <= 16'h6477;
             14'h106f 	:	val_out <= 16'h647d;
             14'h1070 	:	val_out <= 16'h6483;
             14'h1071 	:	val_out <= 16'h6488;
             14'h1072 	:	val_out <= 16'h648e;
             14'h1073 	:	val_out <= 16'h6494;
             14'h1074 	:	val_out <= 16'h649a;
             14'h1075 	:	val_out <= 16'h64a0;
             14'h1076 	:	val_out <= 16'h64a5;
             14'h1077 	:	val_out <= 16'h64ab;
             14'h1078 	:	val_out <= 16'h64b1;
             14'h1079 	:	val_out <= 16'h64b7;
             14'h107a 	:	val_out <= 16'h64bc;
             14'h107b 	:	val_out <= 16'h64c2;
             14'h107c 	:	val_out <= 16'h64c8;
             14'h107d 	:	val_out <= 16'h64ce;
             14'h107e 	:	val_out <= 16'h64d3;
             14'h107f 	:	val_out <= 16'h64d9;
             14'h1080 	:	val_out <= 16'h64df;
             14'h1081 	:	val_out <= 16'h64e5;
             14'h1082 	:	val_out <= 16'h64eb;
             14'h1083 	:	val_out <= 16'h64f0;
             14'h1084 	:	val_out <= 16'h64f6;
             14'h1085 	:	val_out <= 16'h64fc;
             14'h1086 	:	val_out <= 16'h6502;
             14'h1087 	:	val_out <= 16'h6507;
             14'h1088 	:	val_out <= 16'h650d;
             14'h1089 	:	val_out <= 16'h6513;
             14'h108a 	:	val_out <= 16'h6519;
             14'h108b 	:	val_out <= 16'h651f;
             14'h108c 	:	val_out <= 16'h6524;
             14'h108d 	:	val_out <= 16'h652a;
             14'h108e 	:	val_out <= 16'h6530;
             14'h108f 	:	val_out <= 16'h6536;
             14'h1090 	:	val_out <= 16'h653b;
             14'h1091 	:	val_out <= 16'h6541;
             14'h1092 	:	val_out <= 16'h6547;
             14'h1093 	:	val_out <= 16'h654d;
             14'h1094 	:	val_out <= 16'h6552;
             14'h1095 	:	val_out <= 16'h6558;
             14'h1096 	:	val_out <= 16'h655e;
             14'h1097 	:	val_out <= 16'h6564;
             14'h1098 	:	val_out <= 16'h656a;
             14'h1099 	:	val_out <= 16'h656f;
             14'h109a 	:	val_out <= 16'h6575;
             14'h109b 	:	val_out <= 16'h657b;
             14'h109c 	:	val_out <= 16'h6581;
             14'h109d 	:	val_out <= 16'h6586;
             14'h109e 	:	val_out <= 16'h658c;
             14'h109f 	:	val_out <= 16'h6592;
             14'h10a0 	:	val_out <= 16'h6598;
             14'h10a1 	:	val_out <= 16'h659d;
             14'h10a2 	:	val_out <= 16'h65a3;
             14'h10a3 	:	val_out <= 16'h65a9;
             14'h10a4 	:	val_out <= 16'h65af;
             14'h10a5 	:	val_out <= 16'h65b5;
             14'h10a6 	:	val_out <= 16'h65ba;
             14'h10a7 	:	val_out <= 16'h65c0;
             14'h10a8 	:	val_out <= 16'h65c6;
             14'h10a9 	:	val_out <= 16'h65cc;
             14'h10aa 	:	val_out <= 16'h65d1;
             14'h10ab 	:	val_out <= 16'h65d7;
             14'h10ac 	:	val_out <= 16'h65dd;
             14'h10ad 	:	val_out <= 16'h65e3;
             14'h10ae 	:	val_out <= 16'h65e8;
             14'h10af 	:	val_out <= 16'h65ee;
             14'h10b0 	:	val_out <= 16'h65f4;
             14'h10b1 	:	val_out <= 16'h65fa;
             14'h10b2 	:	val_out <= 16'h65ff;
             14'h10b3 	:	val_out <= 16'h6605;
             14'h10b4 	:	val_out <= 16'h660b;
             14'h10b5 	:	val_out <= 16'h6611;
             14'h10b6 	:	val_out <= 16'h6617;
             14'h10b7 	:	val_out <= 16'h661c;
             14'h10b8 	:	val_out <= 16'h6622;
             14'h10b9 	:	val_out <= 16'h6628;
             14'h10ba 	:	val_out <= 16'h662e;
             14'h10bb 	:	val_out <= 16'h6633;
             14'h10bc 	:	val_out <= 16'h6639;
             14'h10bd 	:	val_out <= 16'h663f;
             14'h10be 	:	val_out <= 16'h6645;
             14'h10bf 	:	val_out <= 16'h664a;
             14'h10c0 	:	val_out <= 16'h6650;
             14'h10c1 	:	val_out <= 16'h6656;
             14'h10c2 	:	val_out <= 16'h665c;
             14'h10c3 	:	val_out <= 16'h6661;
             14'h10c4 	:	val_out <= 16'h6667;
             14'h10c5 	:	val_out <= 16'h666d;
             14'h10c6 	:	val_out <= 16'h6673;
             14'h10c7 	:	val_out <= 16'h6678;
             14'h10c8 	:	val_out <= 16'h667e;
             14'h10c9 	:	val_out <= 16'h6684;
             14'h10ca 	:	val_out <= 16'h668a;
             14'h10cb 	:	val_out <= 16'h668f;
             14'h10cc 	:	val_out <= 16'h6695;
             14'h10cd 	:	val_out <= 16'h669b;
             14'h10ce 	:	val_out <= 16'h66a1;
             14'h10cf 	:	val_out <= 16'h66a7;
             14'h10d0 	:	val_out <= 16'h66ac;
             14'h10d1 	:	val_out <= 16'h66b2;
             14'h10d2 	:	val_out <= 16'h66b8;
             14'h10d3 	:	val_out <= 16'h66be;
             14'h10d4 	:	val_out <= 16'h66c3;
             14'h10d5 	:	val_out <= 16'h66c9;
             14'h10d6 	:	val_out <= 16'h66cf;
             14'h10d7 	:	val_out <= 16'h66d5;
             14'h10d8 	:	val_out <= 16'h66da;
             14'h10d9 	:	val_out <= 16'h66e0;
             14'h10da 	:	val_out <= 16'h66e6;
             14'h10db 	:	val_out <= 16'h66ec;
             14'h10dc 	:	val_out <= 16'h66f1;
             14'h10dd 	:	val_out <= 16'h66f7;
             14'h10de 	:	val_out <= 16'h66fd;
             14'h10df 	:	val_out <= 16'h6703;
             14'h10e0 	:	val_out <= 16'h6708;
             14'h10e1 	:	val_out <= 16'h670e;
             14'h10e2 	:	val_out <= 16'h6714;
             14'h10e3 	:	val_out <= 16'h671a;
             14'h10e4 	:	val_out <= 16'h671f;
             14'h10e5 	:	val_out <= 16'h6725;
             14'h10e6 	:	val_out <= 16'h672b;
             14'h10e7 	:	val_out <= 16'h6731;
             14'h10e8 	:	val_out <= 16'h6736;
             14'h10e9 	:	val_out <= 16'h673c;
             14'h10ea 	:	val_out <= 16'h6742;
             14'h10eb 	:	val_out <= 16'h6748;
             14'h10ec 	:	val_out <= 16'h674d;
             14'h10ed 	:	val_out <= 16'h6753;
             14'h10ee 	:	val_out <= 16'h6759;
             14'h10ef 	:	val_out <= 16'h675f;
             14'h10f0 	:	val_out <= 16'h6764;
             14'h10f1 	:	val_out <= 16'h676a;
             14'h10f2 	:	val_out <= 16'h6770;
             14'h10f3 	:	val_out <= 16'h6776;
             14'h10f4 	:	val_out <= 16'h677b;
             14'h10f5 	:	val_out <= 16'h6781;
             14'h10f6 	:	val_out <= 16'h6787;
             14'h10f7 	:	val_out <= 16'h678d;
             14'h10f8 	:	val_out <= 16'h6792;
             14'h10f9 	:	val_out <= 16'h6798;
             14'h10fa 	:	val_out <= 16'h679e;
             14'h10fb 	:	val_out <= 16'h67a4;
             14'h10fc 	:	val_out <= 16'h67a9;
             14'h10fd 	:	val_out <= 16'h67af;
             14'h10fe 	:	val_out <= 16'h67b5;
             14'h10ff 	:	val_out <= 16'h67bb;
             14'h1100 	:	val_out <= 16'h67c0;
             14'h1101 	:	val_out <= 16'h67c6;
             14'h1102 	:	val_out <= 16'h67cc;
             14'h1103 	:	val_out <= 16'h67d1;
             14'h1104 	:	val_out <= 16'h67d7;
             14'h1105 	:	val_out <= 16'h67dd;
             14'h1106 	:	val_out <= 16'h67e3;
             14'h1107 	:	val_out <= 16'h67e8;
             14'h1108 	:	val_out <= 16'h67ee;
             14'h1109 	:	val_out <= 16'h67f4;
             14'h110a 	:	val_out <= 16'h67fa;
             14'h110b 	:	val_out <= 16'h67ff;
             14'h110c 	:	val_out <= 16'h6805;
             14'h110d 	:	val_out <= 16'h680b;
             14'h110e 	:	val_out <= 16'h6811;
             14'h110f 	:	val_out <= 16'h6816;
             14'h1110 	:	val_out <= 16'h681c;
             14'h1111 	:	val_out <= 16'h6822;
             14'h1112 	:	val_out <= 16'h6828;
             14'h1113 	:	val_out <= 16'h682d;
             14'h1114 	:	val_out <= 16'h6833;
             14'h1115 	:	val_out <= 16'h6839;
             14'h1116 	:	val_out <= 16'h683f;
             14'h1117 	:	val_out <= 16'h6844;
             14'h1118 	:	val_out <= 16'h684a;
             14'h1119 	:	val_out <= 16'h6850;
             14'h111a 	:	val_out <= 16'h6856;
             14'h111b 	:	val_out <= 16'h685b;
             14'h111c 	:	val_out <= 16'h6861;
             14'h111d 	:	val_out <= 16'h6867;
             14'h111e 	:	val_out <= 16'h686c;
             14'h111f 	:	val_out <= 16'h6872;
             14'h1120 	:	val_out <= 16'h6878;
             14'h1121 	:	val_out <= 16'h687e;
             14'h1122 	:	val_out <= 16'h6883;
             14'h1123 	:	val_out <= 16'h6889;
             14'h1124 	:	val_out <= 16'h688f;
             14'h1125 	:	val_out <= 16'h6895;
             14'h1126 	:	val_out <= 16'h689a;
             14'h1127 	:	val_out <= 16'h68a0;
             14'h1128 	:	val_out <= 16'h68a6;
             14'h1129 	:	val_out <= 16'h68ac;
             14'h112a 	:	val_out <= 16'h68b1;
             14'h112b 	:	val_out <= 16'h68b7;
             14'h112c 	:	val_out <= 16'h68bd;
             14'h112d 	:	val_out <= 16'h68c3;
             14'h112e 	:	val_out <= 16'h68c8;
             14'h112f 	:	val_out <= 16'h68ce;
             14'h1130 	:	val_out <= 16'h68d4;
             14'h1131 	:	val_out <= 16'h68d9;
             14'h1132 	:	val_out <= 16'h68df;
             14'h1133 	:	val_out <= 16'h68e5;
             14'h1134 	:	val_out <= 16'h68eb;
             14'h1135 	:	val_out <= 16'h68f0;
             14'h1136 	:	val_out <= 16'h68f6;
             14'h1137 	:	val_out <= 16'h68fc;
             14'h1138 	:	val_out <= 16'h6902;
             14'h1139 	:	val_out <= 16'h6907;
             14'h113a 	:	val_out <= 16'h690d;
             14'h113b 	:	val_out <= 16'h6913;
             14'h113c 	:	val_out <= 16'h6918;
             14'h113d 	:	val_out <= 16'h691e;
             14'h113e 	:	val_out <= 16'h6924;
             14'h113f 	:	val_out <= 16'h692a;
             14'h1140 	:	val_out <= 16'h692f;
             14'h1141 	:	val_out <= 16'h6935;
             14'h1142 	:	val_out <= 16'h693b;
             14'h1143 	:	val_out <= 16'h6941;
             14'h1144 	:	val_out <= 16'h6946;
             14'h1145 	:	val_out <= 16'h694c;
             14'h1146 	:	val_out <= 16'h6952;
             14'h1147 	:	val_out <= 16'h6957;
             14'h1148 	:	val_out <= 16'h695d;
             14'h1149 	:	val_out <= 16'h6963;
             14'h114a 	:	val_out <= 16'h6969;
             14'h114b 	:	val_out <= 16'h696e;
             14'h114c 	:	val_out <= 16'h6974;
             14'h114d 	:	val_out <= 16'h697a;
             14'h114e 	:	val_out <= 16'h6980;
             14'h114f 	:	val_out <= 16'h6985;
             14'h1150 	:	val_out <= 16'h698b;
             14'h1151 	:	val_out <= 16'h6991;
             14'h1152 	:	val_out <= 16'h6996;
             14'h1153 	:	val_out <= 16'h699c;
             14'h1154 	:	val_out <= 16'h69a2;
             14'h1155 	:	val_out <= 16'h69a8;
             14'h1156 	:	val_out <= 16'h69ad;
             14'h1157 	:	val_out <= 16'h69b3;
             14'h1158 	:	val_out <= 16'h69b9;
             14'h1159 	:	val_out <= 16'h69bf;
             14'h115a 	:	val_out <= 16'h69c4;
             14'h115b 	:	val_out <= 16'h69ca;
             14'h115c 	:	val_out <= 16'h69d0;
             14'h115d 	:	val_out <= 16'h69d5;
             14'h115e 	:	val_out <= 16'h69db;
             14'h115f 	:	val_out <= 16'h69e1;
             14'h1160 	:	val_out <= 16'h69e7;
             14'h1161 	:	val_out <= 16'h69ec;
             14'h1162 	:	val_out <= 16'h69f2;
             14'h1163 	:	val_out <= 16'h69f8;
             14'h1164 	:	val_out <= 16'h69fd;
             14'h1165 	:	val_out <= 16'h6a03;
             14'h1166 	:	val_out <= 16'h6a09;
             14'h1167 	:	val_out <= 16'h6a0f;
             14'h1168 	:	val_out <= 16'h6a14;
             14'h1169 	:	val_out <= 16'h6a1a;
             14'h116a 	:	val_out <= 16'h6a20;
             14'h116b 	:	val_out <= 16'h6a25;
             14'h116c 	:	val_out <= 16'h6a2b;
             14'h116d 	:	val_out <= 16'h6a31;
             14'h116e 	:	val_out <= 16'h6a37;
             14'h116f 	:	val_out <= 16'h6a3c;
             14'h1170 	:	val_out <= 16'h6a42;
             14'h1171 	:	val_out <= 16'h6a48;
             14'h1172 	:	val_out <= 16'h6a4d;
             14'h1173 	:	val_out <= 16'h6a53;
             14'h1174 	:	val_out <= 16'h6a59;
             14'h1175 	:	val_out <= 16'h6a5f;
             14'h1176 	:	val_out <= 16'h6a64;
             14'h1177 	:	val_out <= 16'h6a6a;
             14'h1178 	:	val_out <= 16'h6a70;
             14'h1179 	:	val_out <= 16'h6a75;
             14'h117a 	:	val_out <= 16'h6a7b;
             14'h117b 	:	val_out <= 16'h6a81;
             14'h117c 	:	val_out <= 16'h6a87;
             14'h117d 	:	val_out <= 16'h6a8c;
             14'h117e 	:	val_out <= 16'h6a92;
             14'h117f 	:	val_out <= 16'h6a98;
             14'h1180 	:	val_out <= 16'h6a9d;
             14'h1181 	:	val_out <= 16'h6aa3;
             14'h1182 	:	val_out <= 16'h6aa9;
             14'h1183 	:	val_out <= 16'h6aaf;
             14'h1184 	:	val_out <= 16'h6ab4;
             14'h1185 	:	val_out <= 16'h6aba;
             14'h1186 	:	val_out <= 16'h6ac0;
             14'h1187 	:	val_out <= 16'h6ac5;
             14'h1188 	:	val_out <= 16'h6acb;
             14'h1189 	:	val_out <= 16'h6ad1;
             14'h118a 	:	val_out <= 16'h6ad7;
             14'h118b 	:	val_out <= 16'h6adc;
             14'h118c 	:	val_out <= 16'h6ae2;
             14'h118d 	:	val_out <= 16'h6ae8;
             14'h118e 	:	val_out <= 16'h6aed;
             14'h118f 	:	val_out <= 16'h6af3;
             14'h1190 	:	val_out <= 16'h6af9;
             14'h1191 	:	val_out <= 16'h6aff;
             14'h1192 	:	val_out <= 16'h6b04;
             14'h1193 	:	val_out <= 16'h6b0a;
             14'h1194 	:	val_out <= 16'h6b10;
             14'h1195 	:	val_out <= 16'h6b15;
             14'h1196 	:	val_out <= 16'h6b1b;
             14'h1197 	:	val_out <= 16'h6b21;
             14'h1198 	:	val_out <= 16'h6b27;
             14'h1199 	:	val_out <= 16'h6b2c;
             14'h119a 	:	val_out <= 16'h6b32;
             14'h119b 	:	val_out <= 16'h6b38;
             14'h119c 	:	val_out <= 16'h6b3d;
             14'h119d 	:	val_out <= 16'h6b43;
             14'h119e 	:	val_out <= 16'h6b49;
             14'h119f 	:	val_out <= 16'h6b4e;
             14'h11a0 	:	val_out <= 16'h6b54;
             14'h11a1 	:	val_out <= 16'h6b5a;
             14'h11a2 	:	val_out <= 16'h6b60;
             14'h11a3 	:	val_out <= 16'h6b65;
             14'h11a4 	:	val_out <= 16'h6b6b;
             14'h11a5 	:	val_out <= 16'h6b71;
             14'h11a6 	:	val_out <= 16'h6b76;
             14'h11a7 	:	val_out <= 16'h6b7c;
             14'h11a8 	:	val_out <= 16'h6b82;
             14'h11a9 	:	val_out <= 16'h6b87;
             14'h11aa 	:	val_out <= 16'h6b8d;
             14'h11ab 	:	val_out <= 16'h6b93;
             14'h11ac 	:	val_out <= 16'h6b99;
             14'h11ad 	:	val_out <= 16'h6b9e;
             14'h11ae 	:	val_out <= 16'h6ba4;
             14'h11af 	:	val_out <= 16'h6baa;
             14'h11b0 	:	val_out <= 16'h6baf;
             14'h11b1 	:	val_out <= 16'h6bb5;
             14'h11b2 	:	val_out <= 16'h6bbb;
             14'h11b3 	:	val_out <= 16'h6bc0;
             14'h11b4 	:	val_out <= 16'h6bc6;
             14'h11b5 	:	val_out <= 16'h6bcc;
             14'h11b6 	:	val_out <= 16'h6bd2;
             14'h11b7 	:	val_out <= 16'h6bd7;
             14'h11b8 	:	val_out <= 16'h6bdd;
             14'h11b9 	:	val_out <= 16'h6be3;
             14'h11ba 	:	val_out <= 16'h6be8;
             14'h11bb 	:	val_out <= 16'h6bee;
             14'h11bc 	:	val_out <= 16'h6bf4;
             14'h11bd 	:	val_out <= 16'h6bf9;
             14'h11be 	:	val_out <= 16'h6bff;
             14'h11bf 	:	val_out <= 16'h6c05;
             14'h11c0 	:	val_out <= 16'h6c0b;
             14'h11c1 	:	val_out <= 16'h6c10;
             14'h11c2 	:	val_out <= 16'h6c16;
             14'h11c3 	:	val_out <= 16'h6c1c;
             14'h11c4 	:	val_out <= 16'h6c21;
             14'h11c5 	:	val_out <= 16'h6c27;
             14'h11c6 	:	val_out <= 16'h6c2d;
             14'h11c7 	:	val_out <= 16'h6c32;
             14'h11c8 	:	val_out <= 16'h6c38;
             14'h11c9 	:	val_out <= 16'h6c3e;
             14'h11ca 	:	val_out <= 16'h6c44;
             14'h11cb 	:	val_out <= 16'h6c49;
             14'h11cc 	:	val_out <= 16'h6c4f;
             14'h11cd 	:	val_out <= 16'h6c55;
             14'h11ce 	:	val_out <= 16'h6c5a;
             14'h11cf 	:	val_out <= 16'h6c60;
             14'h11d0 	:	val_out <= 16'h6c66;
             14'h11d1 	:	val_out <= 16'h6c6b;
             14'h11d2 	:	val_out <= 16'h6c71;
             14'h11d3 	:	val_out <= 16'h6c77;
             14'h11d4 	:	val_out <= 16'h6c7c;
             14'h11d5 	:	val_out <= 16'h6c82;
             14'h11d6 	:	val_out <= 16'h6c88;
             14'h11d7 	:	val_out <= 16'h6c8e;
             14'h11d8 	:	val_out <= 16'h6c93;
             14'h11d9 	:	val_out <= 16'h6c99;
             14'h11da 	:	val_out <= 16'h6c9f;
             14'h11db 	:	val_out <= 16'h6ca4;
             14'h11dc 	:	val_out <= 16'h6caa;
             14'h11dd 	:	val_out <= 16'h6cb0;
             14'h11de 	:	val_out <= 16'h6cb5;
             14'h11df 	:	val_out <= 16'h6cbb;
             14'h11e0 	:	val_out <= 16'h6cc1;
             14'h11e1 	:	val_out <= 16'h6cc6;
             14'h11e2 	:	val_out <= 16'h6ccc;
             14'h11e3 	:	val_out <= 16'h6cd2;
             14'h11e4 	:	val_out <= 16'h6cd7;
             14'h11e5 	:	val_out <= 16'h6cdd;
             14'h11e6 	:	val_out <= 16'h6ce3;
             14'h11e7 	:	val_out <= 16'h6ce9;
             14'h11e8 	:	val_out <= 16'h6cee;
             14'h11e9 	:	val_out <= 16'h6cf4;
             14'h11ea 	:	val_out <= 16'h6cfa;
             14'h11eb 	:	val_out <= 16'h6cff;
             14'h11ec 	:	val_out <= 16'h6d05;
             14'h11ed 	:	val_out <= 16'h6d0b;
             14'h11ee 	:	val_out <= 16'h6d10;
             14'h11ef 	:	val_out <= 16'h6d16;
             14'h11f0 	:	val_out <= 16'h6d1c;
             14'h11f1 	:	val_out <= 16'h6d21;
             14'h11f2 	:	val_out <= 16'h6d27;
             14'h11f3 	:	val_out <= 16'h6d2d;
             14'h11f4 	:	val_out <= 16'h6d32;
             14'h11f5 	:	val_out <= 16'h6d38;
             14'h11f6 	:	val_out <= 16'h6d3e;
             14'h11f7 	:	val_out <= 16'h6d43;
             14'h11f8 	:	val_out <= 16'h6d49;
             14'h11f9 	:	val_out <= 16'h6d4f;
             14'h11fa 	:	val_out <= 16'h6d55;
             14'h11fb 	:	val_out <= 16'h6d5a;
             14'h11fc 	:	val_out <= 16'h6d60;
             14'h11fd 	:	val_out <= 16'h6d66;
             14'h11fe 	:	val_out <= 16'h6d6b;
             14'h11ff 	:	val_out <= 16'h6d71;
             14'h1200 	:	val_out <= 16'h6d77;
             14'h1201 	:	val_out <= 16'h6d7c;
             14'h1202 	:	val_out <= 16'h6d82;
             14'h1203 	:	val_out <= 16'h6d88;
             14'h1204 	:	val_out <= 16'h6d8d;
             14'h1205 	:	val_out <= 16'h6d93;
             14'h1206 	:	val_out <= 16'h6d99;
             14'h1207 	:	val_out <= 16'h6d9e;
             14'h1208 	:	val_out <= 16'h6da4;
             14'h1209 	:	val_out <= 16'h6daa;
             14'h120a 	:	val_out <= 16'h6daf;
             14'h120b 	:	val_out <= 16'h6db5;
             14'h120c 	:	val_out <= 16'h6dbb;
             14'h120d 	:	val_out <= 16'h6dc0;
             14'h120e 	:	val_out <= 16'h6dc6;
             14'h120f 	:	val_out <= 16'h6dcc;
             14'h1210 	:	val_out <= 16'h6dd1;
             14'h1211 	:	val_out <= 16'h6dd7;
             14'h1212 	:	val_out <= 16'h6ddd;
             14'h1213 	:	val_out <= 16'h6de2;
             14'h1214 	:	val_out <= 16'h6de8;
             14'h1215 	:	val_out <= 16'h6dee;
             14'h1216 	:	val_out <= 16'h6df3;
             14'h1217 	:	val_out <= 16'h6df9;
             14'h1218 	:	val_out <= 16'h6dff;
             14'h1219 	:	val_out <= 16'h6e05;
             14'h121a 	:	val_out <= 16'h6e0a;
             14'h121b 	:	val_out <= 16'h6e10;
             14'h121c 	:	val_out <= 16'h6e16;
             14'h121d 	:	val_out <= 16'h6e1b;
             14'h121e 	:	val_out <= 16'h6e21;
             14'h121f 	:	val_out <= 16'h6e27;
             14'h1220 	:	val_out <= 16'h6e2c;
             14'h1221 	:	val_out <= 16'h6e32;
             14'h1222 	:	val_out <= 16'h6e38;
             14'h1223 	:	val_out <= 16'h6e3d;
             14'h1224 	:	val_out <= 16'h6e43;
             14'h1225 	:	val_out <= 16'h6e49;
             14'h1226 	:	val_out <= 16'h6e4e;
             14'h1227 	:	val_out <= 16'h6e54;
             14'h1228 	:	val_out <= 16'h6e5a;
             14'h1229 	:	val_out <= 16'h6e5f;
             14'h122a 	:	val_out <= 16'h6e65;
             14'h122b 	:	val_out <= 16'h6e6b;
             14'h122c 	:	val_out <= 16'h6e70;
             14'h122d 	:	val_out <= 16'h6e76;
             14'h122e 	:	val_out <= 16'h6e7c;
             14'h122f 	:	val_out <= 16'h6e81;
             14'h1230 	:	val_out <= 16'h6e87;
             14'h1231 	:	val_out <= 16'h6e8d;
             14'h1232 	:	val_out <= 16'h6e92;
             14'h1233 	:	val_out <= 16'h6e98;
             14'h1234 	:	val_out <= 16'h6e9e;
             14'h1235 	:	val_out <= 16'h6ea3;
             14'h1236 	:	val_out <= 16'h6ea9;
             14'h1237 	:	val_out <= 16'h6eaf;
             14'h1238 	:	val_out <= 16'h6eb4;
             14'h1239 	:	val_out <= 16'h6eba;
             14'h123a 	:	val_out <= 16'h6ec0;
             14'h123b 	:	val_out <= 16'h6ec5;
             14'h123c 	:	val_out <= 16'h6ecb;
             14'h123d 	:	val_out <= 16'h6ed1;
             14'h123e 	:	val_out <= 16'h6ed6;
             14'h123f 	:	val_out <= 16'h6edc;
             14'h1240 	:	val_out <= 16'h6ee2;
             14'h1241 	:	val_out <= 16'h6ee7;
             14'h1242 	:	val_out <= 16'h6eed;
             14'h1243 	:	val_out <= 16'h6ef3;
             14'h1244 	:	val_out <= 16'h6ef8;
             14'h1245 	:	val_out <= 16'h6efe;
             14'h1246 	:	val_out <= 16'h6f04;
             14'h1247 	:	val_out <= 16'h6f09;
             14'h1248 	:	val_out <= 16'h6f0f;
             14'h1249 	:	val_out <= 16'h6f15;
             14'h124a 	:	val_out <= 16'h6f1a;
             14'h124b 	:	val_out <= 16'h6f20;
             14'h124c 	:	val_out <= 16'h6f26;
             14'h124d 	:	val_out <= 16'h6f2b;
             14'h124e 	:	val_out <= 16'h6f31;
             14'h124f 	:	val_out <= 16'h6f36;
             14'h1250 	:	val_out <= 16'h6f3c;
             14'h1251 	:	val_out <= 16'h6f42;
             14'h1252 	:	val_out <= 16'h6f47;
             14'h1253 	:	val_out <= 16'h6f4d;
             14'h1254 	:	val_out <= 16'h6f53;
             14'h1255 	:	val_out <= 16'h6f58;
             14'h1256 	:	val_out <= 16'h6f5e;
             14'h1257 	:	val_out <= 16'h6f64;
             14'h1258 	:	val_out <= 16'h6f69;
             14'h1259 	:	val_out <= 16'h6f6f;
             14'h125a 	:	val_out <= 16'h6f75;
             14'h125b 	:	val_out <= 16'h6f7a;
             14'h125c 	:	val_out <= 16'h6f80;
             14'h125d 	:	val_out <= 16'h6f86;
             14'h125e 	:	val_out <= 16'h6f8b;
             14'h125f 	:	val_out <= 16'h6f91;
             14'h1260 	:	val_out <= 16'h6f97;
             14'h1261 	:	val_out <= 16'h6f9c;
             14'h1262 	:	val_out <= 16'h6fa2;
             14'h1263 	:	val_out <= 16'h6fa8;
             14'h1264 	:	val_out <= 16'h6fad;
             14'h1265 	:	val_out <= 16'h6fb3;
             14'h1266 	:	val_out <= 16'h6fb9;
             14'h1267 	:	val_out <= 16'h6fbe;
             14'h1268 	:	val_out <= 16'h6fc4;
             14'h1269 	:	val_out <= 16'h6fca;
             14'h126a 	:	val_out <= 16'h6fcf;
             14'h126b 	:	val_out <= 16'h6fd5;
             14'h126c 	:	val_out <= 16'h6fda;
             14'h126d 	:	val_out <= 16'h6fe0;
             14'h126e 	:	val_out <= 16'h6fe6;
             14'h126f 	:	val_out <= 16'h6feb;
             14'h1270 	:	val_out <= 16'h6ff1;
             14'h1271 	:	val_out <= 16'h6ff7;
             14'h1272 	:	val_out <= 16'h6ffc;
             14'h1273 	:	val_out <= 16'h7002;
             14'h1274 	:	val_out <= 16'h7008;
             14'h1275 	:	val_out <= 16'h700d;
             14'h1276 	:	val_out <= 16'h7013;
             14'h1277 	:	val_out <= 16'h7019;
             14'h1278 	:	val_out <= 16'h701e;
             14'h1279 	:	val_out <= 16'h7024;
             14'h127a 	:	val_out <= 16'h702a;
             14'h127b 	:	val_out <= 16'h702f;
             14'h127c 	:	val_out <= 16'h7035;
             14'h127d 	:	val_out <= 16'h703b;
             14'h127e 	:	val_out <= 16'h7040;
             14'h127f 	:	val_out <= 16'h7046;
             14'h1280 	:	val_out <= 16'h704b;
             14'h1281 	:	val_out <= 16'h7051;
             14'h1282 	:	val_out <= 16'h7057;
             14'h1283 	:	val_out <= 16'h705c;
             14'h1284 	:	val_out <= 16'h7062;
             14'h1285 	:	val_out <= 16'h7068;
             14'h1286 	:	val_out <= 16'h706d;
             14'h1287 	:	val_out <= 16'h7073;
             14'h1288 	:	val_out <= 16'h7079;
             14'h1289 	:	val_out <= 16'h707e;
             14'h128a 	:	val_out <= 16'h7084;
             14'h128b 	:	val_out <= 16'h708a;
             14'h128c 	:	val_out <= 16'h708f;
             14'h128d 	:	val_out <= 16'h7095;
             14'h128e 	:	val_out <= 16'h709b;
             14'h128f 	:	val_out <= 16'h70a0;
             14'h1290 	:	val_out <= 16'h70a6;
             14'h1291 	:	val_out <= 16'h70ab;
             14'h1292 	:	val_out <= 16'h70b1;
             14'h1293 	:	val_out <= 16'h70b7;
             14'h1294 	:	val_out <= 16'h70bc;
             14'h1295 	:	val_out <= 16'h70c2;
             14'h1296 	:	val_out <= 16'h70c8;
             14'h1297 	:	val_out <= 16'h70cd;
             14'h1298 	:	val_out <= 16'h70d3;
             14'h1299 	:	val_out <= 16'h70d9;
             14'h129a 	:	val_out <= 16'h70de;
             14'h129b 	:	val_out <= 16'h70e4;
             14'h129c 	:	val_out <= 16'h70e9;
             14'h129d 	:	val_out <= 16'h70ef;
             14'h129e 	:	val_out <= 16'h70f5;
             14'h129f 	:	val_out <= 16'h70fa;
             14'h12a0 	:	val_out <= 16'h7100;
             14'h12a1 	:	val_out <= 16'h7106;
             14'h12a2 	:	val_out <= 16'h710b;
             14'h12a3 	:	val_out <= 16'h7111;
             14'h12a4 	:	val_out <= 16'h7117;
             14'h12a5 	:	val_out <= 16'h711c;
             14'h12a6 	:	val_out <= 16'h7122;
             14'h12a7 	:	val_out <= 16'h7127;
             14'h12a8 	:	val_out <= 16'h712d;
             14'h12a9 	:	val_out <= 16'h7133;
             14'h12aa 	:	val_out <= 16'h7138;
             14'h12ab 	:	val_out <= 16'h713e;
             14'h12ac 	:	val_out <= 16'h7144;
             14'h12ad 	:	val_out <= 16'h7149;
             14'h12ae 	:	val_out <= 16'h714f;
             14'h12af 	:	val_out <= 16'h7155;
             14'h12b0 	:	val_out <= 16'h715a;
             14'h12b1 	:	val_out <= 16'h7160;
             14'h12b2 	:	val_out <= 16'h7165;
             14'h12b3 	:	val_out <= 16'h716b;
             14'h12b4 	:	val_out <= 16'h7171;
             14'h12b5 	:	val_out <= 16'h7176;
             14'h12b6 	:	val_out <= 16'h717c;
             14'h12b7 	:	val_out <= 16'h7182;
             14'h12b8 	:	val_out <= 16'h7187;
             14'h12b9 	:	val_out <= 16'h718d;
             14'h12ba 	:	val_out <= 16'h7193;
             14'h12bb 	:	val_out <= 16'h7198;
             14'h12bc 	:	val_out <= 16'h719e;
             14'h12bd 	:	val_out <= 16'h71a3;
             14'h12be 	:	val_out <= 16'h71a9;
             14'h12bf 	:	val_out <= 16'h71af;
             14'h12c0 	:	val_out <= 16'h71b4;
             14'h12c1 	:	val_out <= 16'h71ba;
             14'h12c2 	:	val_out <= 16'h71c0;
             14'h12c3 	:	val_out <= 16'h71c5;
             14'h12c4 	:	val_out <= 16'h71cb;
             14'h12c5 	:	val_out <= 16'h71d0;
             14'h12c6 	:	val_out <= 16'h71d6;
             14'h12c7 	:	val_out <= 16'h71dc;
             14'h12c8 	:	val_out <= 16'h71e1;
             14'h12c9 	:	val_out <= 16'h71e7;
             14'h12ca 	:	val_out <= 16'h71ed;
             14'h12cb 	:	val_out <= 16'h71f2;
             14'h12cc 	:	val_out <= 16'h71f8;
             14'h12cd 	:	val_out <= 16'h71fd;
             14'h12ce 	:	val_out <= 16'h7203;
             14'h12cf 	:	val_out <= 16'h7209;
             14'h12d0 	:	val_out <= 16'h720e;
             14'h12d1 	:	val_out <= 16'h7214;
             14'h12d2 	:	val_out <= 16'h721a;
             14'h12d3 	:	val_out <= 16'h721f;
             14'h12d4 	:	val_out <= 16'h7225;
             14'h12d5 	:	val_out <= 16'h722a;
             14'h12d6 	:	val_out <= 16'h7230;
             14'h12d7 	:	val_out <= 16'h7236;
             14'h12d8 	:	val_out <= 16'h723b;
             14'h12d9 	:	val_out <= 16'h7241;
             14'h12da 	:	val_out <= 16'h7247;
             14'h12db 	:	val_out <= 16'h724c;
             14'h12dc 	:	val_out <= 16'h7252;
             14'h12dd 	:	val_out <= 16'h7257;
             14'h12de 	:	val_out <= 16'h725d;
             14'h12df 	:	val_out <= 16'h7263;
             14'h12e0 	:	val_out <= 16'h7268;
             14'h12e1 	:	val_out <= 16'h726e;
             14'h12e2 	:	val_out <= 16'h7274;
             14'h12e3 	:	val_out <= 16'h7279;
             14'h12e4 	:	val_out <= 16'h727f;
             14'h12e5 	:	val_out <= 16'h7284;
             14'h12e6 	:	val_out <= 16'h728a;
             14'h12e7 	:	val_out <= 16'h7290;
             14'h12e8 	:	val_out <= 16'h7295;
             14'h12e9 	:	val_out <= 16'h729b;
             14'h12ea 	:	val_out <= 16'h72a1;
             14'h12eb 	:	val_out <= 16'h72a6;
             14'h12ec 	:	val_out <= 16'h72ac;
             14'h12ed 	:	val_out <= 16'h72b1;
             14'h12ee 	:	val_out <= 16'h72b7;
             14'h12ef 	:	val_out <= 16'h72bd;
             14'h12f0 	:	val_out <= 16'h72c2;
             14'h12f1 	:	val_out <= 16'h72c8;
             14'h12f2 	:	val_out <= 16'h72cd;
             14'h12f3 	:	val_out <= 16'h72d3;
             14'h12f4 	:	val_out <= 16'h72d9;
             14'h12f5 	:	val_out <= 16'h72de;
             14'h12f6 	:	val_out <= 16'h72e4;
             14'h12f7 	:	val_out <= 16'h72ea;
             14'h12f8 	:	val_out <= 16'h72ef;
             14'h12f9 	:	val_out <= 16'h72f5;
             14'h12fa 	:	val_out <= 16'h72fa;
             14'h12fb 	:	val_out <= 16'h7300;
             14'h12fc 	:	val_out <= 16'h7306;
             14'h12fd 	:	val_out <= 16'h730b;
             14'h12fe 	:	val_out <= 16'h7311;
             14'h12ff 	:	val_out <= 16'h7316;
             14'h1300 	:	val_out <= 16'h731c;
             14'h1301 	:	val_out <= 16'h7322;
             14'h1302 	:	val_out <= 16'h7327;
             14'h1303 	:	val_out <= 16'h732d;
             14'h1304 	:	val_out <= 16'h7332;
             14'h1305 	:	val_out <= 16'h7338;
             14'h1306 	:	val_out <= 16'h733e;
             14'h1307 	:	val_out <= 16'h7343;
             14'h1308 	:	val_out <= 16'h7349;
             14'h1309 	:	val_out <= 16'h734f;
             14'h130a 	:	val_out <= 16'h7354;
             14'h130b 	:	val_out <= 16'h735a;
             14'h130c 	:	val_out <= 16'h735f;
             14'h130d 	:	val_out <= 16'h7365;
             14'h130e 	:	val_out <= 16'h736b;
             14'h130f 	:	val_out <= 16'h7370;
             14'h1310 	:	val_out <= 16'h7376;
             14'h1311 	:	val_out <= 16'h737b;
             14'h1312 	:	val_out <= 16'h7381;
             14'h1313 	:	val_out <= 16'h7387;
             14'h1314 	:	val_out <= 16'h738c;
             14'h1315 	:	val_out <= 16'h7392;
             14'h1316 	:	val_out <= 16'h7397;
             14'h1317 	:	val_out <= 16'h739d;
             14'h1318 	:	val_out <= 16'h73a3;
             14'h1319 	:	val_out <= 16'h73a8;
             14'h131a 	:	val_out <= 16'h73ae;
             14'h131b 	:	val_out <= 16'h73b3;
             14'h131c 	:	val_out <= 16'h73b9;
             14'h131d 	:	val_out <= 16'h73bf;
             14'h131e 	:	val_out <= 16'h73c4;
             14'h131f 	:	val_out <= 16'h73ca;
             14'h1320 	:	val_out <= 16'h73cf;
             14'h1321 	:	val_out <= 16'h73d5;
             14'h1322 	:	val_out <= 16'h73db;
             14'h1323 	:	val_out <= 16'h73e0;
             14'h1324 	:	val_out <= 16'h73e6;
             14'h1325 	:	val_out <= 16'h73eb;
             14'h1326 	:	val_out <= 16'h73f1;
             14'h1327 	:	val_out <= 16'h73f7;
             14'h1328 	:	val_out <= 16'h73fc;
             14'h1329 	:	val_out <= 16'h7402;
             14'h132a 	:	val_out <= 16'h7408;
             14'h132b 	:	val_out <= 16'h740d;
             14'h132c 	:	val_out <= 16'h7413;
             14'h132d 	:	val_out <= 16'h7418;
             14'h132e 	:	val_out <= 16'h741e;
             14'h132f 	:	val_out <= 16'h7424;
             14'h1330 	:	val_out <= 16'h7429;
             14'h1331 	:	val_out <= 16'h742f;
             14'h1332 	:	val_out <= 16'h7434;
             14'h1333 	:	val_out <= 16'h743a;
             14'h1334 	:	val_out <= 16'h743f;
             14'h1335 	:	val_out <= 16'h7445;
             14'h1336 	:	val_out <= 16'h744b;
             14'h1337 	:	val_out <= 16'h7450;
             14'h1338 	:	val_out <= 16'h7456;
             14'h1339 	:	val_out <= 16'h745b;
             14'h133a 	:	val_out <= 16'h7461;
             14'h133b 	:	val_out <= 16'h7467;
             14'h133c 	:	val_out <= 16'h746c;
             14'h133d 	:	val_out <= 16'h7472;
             14'h133e 	:	val_out <= 16'h7477;
             14'h133f 	:	val_out <= 16'h747d;
             14'h1340 	:	val_out <= 16'h7483;
             14'h1341 	:	val_out <= 16'h7488;
             14'h1342 	:	val_out <= 16'h748e;
             14'h1343 	:	val_out <= 16'h7493;
             14'h1344 	:	val_out <= 16'h7499;
             14'h1345 	:	val_out <= 16'h749f;
             14'h1346 	:	val_out <= 16'h74a4;
             14'h1347 	:	val_out <= 16'h74aa;
             14'h1348 	:	val_out <= 16'h74af;
             14'h1349 	:	val_out <= 16'h74b5;
             14'h134a 	:	val_out <= 16'h74bb;
             14'h134b 	:	val_out <= 16'h74c0;
             14'h134c 	:	val_out <= 16'h74c6;
             14'h134d 	:	val_out <= 16'h74cb;
             14'h134e 	:	val_out <= 16'h74d1;
             14'h134f 	:	val_out <= 16'h74d7;
             14'h1350 	:	val_out <= 16'h74dc;
             14'h1351 	:	val_out <= 16'h74e2;
             14'h1352 	:	val_out <= 16'h74e7;
             14'h1353 	:	val_out <= 16'h74ed;
             14'h1354 	:	val_out <= 16'h74f2;
             14'h1355 	:	val_out <= 16'h74f8;
             14'h1356 	:	val_out <= 16'h74fe;
             14'h1357 	:	val_out <= 16'h7503;
             14'h1358 	:	val_out <= 16'h7509;
             14'h1359 	:	val_out <= 16'h750e;
             14'h135a 	:	val_out <= 16'h7514;
             14'h135b 	:	val_out <= 16'h751a;
             14'h135c 	:	val_out <= 16'h751f;
             14'h135d 	:	val_out <= 16'h7525;
             14'h135e 	:	val_out <= 16'h752a;
             14'h135f 	:	val_out <= 16'h7530;
             14'h1360 	:	val_out <= 16'h7536;
             14'h1361 	:	val_out <= 16'h753b;
             14'h1362 	:	val_out <= 16'h7541;
             14'h1363 	:	val_out <= 16'h7546;
             14'h1364 	:	val_out <= 16'h754c;
             14'h1365 	:	val_out <= 16'h7551;
             14'h1366 	:	val_out <= 16'h7557;
             14'h1367 	:	val_out <= 16'h755d;
             14'h1368 	:	val_out <= 16'h7562;
             14'h1369 	:	val_out <= 16'h7568;
             14'h136a 	:	val_out <= 16'h756d;
             14'h136b 	:	val_out <= 16'h7573;
             14'h136c 	:	val_out <= 16'h7579;
             14'h136d 	:	val_out <= 16'h757e;
             14'h136e 	:	val_out <= 16'h7584;
             14'h136f 	:	val_out <= 16'h7589;
             14'h1370 	:	val_out <= 16'h758f;
             14'h1371 	:	val_out <= 16'h7594;
             14'h1372 	:	val_out <= 16'h759a;
             14'h1373 	:	val_out <= 16'h75a0;
             14'h1374 	:	val_out <= 16'h75a5;
             14'h1375 	:	val_out <= 16'h75ab;
             14'h1376 	:	val_out <= 16'h75b0;
             14'h1377 	:	val_out <= 16'h75b6;
             14'h1378 	:	val_out <= 16'h75bc;
             14'h1379 	:	val_out <= 16'h75c1;
             14'h137a 	:	val_out <= 16'h75c7;
             14'h137b 	:	val_out <= 16'h75cc;
             14'h137c 	:	val_out <= 16'h75d2;
             14'h137d 	:	val_out <= 16'h75d7;
             14'h137e 	:	val_out <= 16'h75dd;
             14'h137f 	:	val_out <= 16'h75e3;
             14'h1380 	:	val_out <= 16'h75e8;
             14'h1381 	:	val_out <= 16'h75ee;
             14'h1382 	:	val_out <= 16'h75f3;
             14'h1383 	:	val_out <= 16'h75f9;
             14'h1384 	:	val_out <= 16'h75fe;
             14'h1385 	:	val_out <= 16'h7604;
             14'h1386 	:	val_out <= 16'h760a;
             14'h1387 	:	val_out <= 16'h760f;
             14'h1388 	:	val_out <= 16'h7615;
             14'h1389 	:	val_out <= 16'h761a;
             14'h138a 	:	val_out <= 16'h7620;
             14'h138b 	:	val_out <= 16'h7625;
             14'h138c 	:	val_out <= 16'h762b;
             14'h138d 	:	val_out <= 16'h7631;
             14'h138e 	:	val_out <= 16'h7636;
             14'h138f 	:	val_out <= 16'h763c;
             14'h1390 	:	val_out <= 16'h7641;
             14'h1391 	:	val_out <= 16'h7647;
             14'h1392 	:	val_out <= 16'h764c;
             14'h1393 	:	val_out <= 16'h7652;
             14'h1394 	:	val_out <= 16'h7658;
             14'h1395 	:	val_out <= 16'h765d;
             14'h1396 	:	val_out <= 16'h7663;
             14'h1397 	:	val_out <= 16'h7668;
             14'h1398 	:	val_out <= 16'h766e;
             14'h1399 	:	val_out <= 16'h7673;
             14'h139a 	:	val_out <= 16'h7679;
             14'h139b 	:	val_out <= 16'h767f;
             14'h139c 	:	val_out <= 16'h7684;
             14'h139d 	:	val_out <= 16'h768a;
             14'h139e 	:	val_out <= 16'h768f;
             14'h139f 	:	val_out <= 16'h7695;
             14'h13a0 	:	val_out <= 16'h769a;
             14'h13a1 	:	val_out <= 16'h76a0;
             14'h13a2 	:	val_out <= 16'h76a6;
             14'h13a3 	:	val_out <= 16'h76ab;
             14'h13a4 	:	val_out <= 16'h76b1;
             14'h13a5 	:	val_out <= 16'h76b6;
             14'h13a6 	:	val_out <= 16'h76bc;
             14'h13a7 	:	val_out <= 16'h76c1;
             14'h13a8 	:	val_out <= 16'h76c7;
             14'h13a9 	:	val_out <= 16'h76cd;
             14'h13aa 	:	val_out <= 16'h76d2;
             14'h13ab 	:	val_out <= 16'h76d8;
             14'h13ac 	:	val_out <= 16'h76dd;
             14'h13ad 	:	val_out <= 16'h76e3;
             14'h13ae 	:	val_out <= 16'h76e8;
             14'h13af 	:	val_out <= 16'h76ee;
             14'h13b0 	:	val_out <= 16'h76f4;
             14'h13b1 	:	val_out <= 16'h76f9;
             14'h13b2 	:	val_out <= 16'h76ff;
             14'h13b3 	:	val_out <= 16'h7704;
             14'h13b4 	:	val_out <= 16'h770a;
             14'h13b5 	:	val_out <= 16'h770f;
             14'h13b6 	:	val_out <= 16'h7715;
             14'h13b7 	:	val_out <= 16'h771a;
             14'h13b8 	:	val_out <= 16'h7720;
             14'h13b9 	:	val_out <= 16'h7726;
             14'h13ba 	:	val_out <= 16'h772b;
             14'h13bb 	:	val_out <= 16'h7731;
             14'h13bc 	:	val_out <= 16'h7736;
             14'h13bd 	:	val_out <= 16'h773c;
             14'h13be 	:	val_out <= 16'h7741;
             14'h13bf 	:	val_out <= 16'h7747;
             14'h13c0 	:	val_out <= 16'h774d;
             14'h13c1 	:	val_out <= 16'h7752;
             14'h13c2 	:	val_out <= 16'h7758;
             14'h13c3 	:	val_out <= 16'h775d;
             14'h13c4 	:	val_out <= 16'h7763;
             14'h13c5 	:	val_out <= 16'h7768;
             14'h13c6 	:	val_out <= 16'h776e;
             14'h13c7 	:	val_out <= 16'h7773;
             14'h13c8 	:	val_out <= 16'h7779;
             14'h13c9 	:	val_out <= 16'h777f;
             14'h13ca 	:	val_out <= 16'h7784;
             14'h13cb 	:	val_out <= 16'h778a;
             14'h13cc 	:	val_out <= 16'h778f;
             14'h13cd 	:	val_out <= 16'h7795;
             14'h13ce 	:	val_out <= 16'h779a;
             14'h13cf 	:	val_out <= 16'h77a0;
             14'h13d0 	:	val_out <= 16'h77a5;
             14'h13d1 	:	val_out <= 16'h77ab;
             14'h13d2 	:	val_out <= 16'h77b1;
             14'h13d3 	:	val_out <= 16'h77b6;
             14'h13d4 	:	val_out <= 16'h77bc;
             14'h13d5 	:	val_out <= 16'h77c1;
             14'h13d6 	:	val_out <= 16'h77c7;
             14'h13d7 	:	val_out <= 16'h77cc;
             14'h13d8 	:	val_out <= 16'h77d2;
             14'h13d9 	:	val_out <= 16'h77d7;
             14'h13da 	:	val_out <= 16'h77dd;
             14'h13db 	:	val_out <= 16'h77e3;
             14'h13dc 	:	val_out <= 16'h77e8;
             14'h13dd 	:	val_out <= 16'h77ee;
             14'h13de 	:	val_out <= 16'h77f3;
             14'h13df 	:	val_out <= 16'h77f9;
             14'h13e0 	:	val_out <= 16'h77fe;
             14'h13e1 	:	val_out <= 16'h7804;
             14'h13e2 	:	val_out <= 16'h7809;
             14'h13e3 	:	val_out <= 16'h780f;
             14'h13e4 	:	val_out <= 16'h7814;
             14'h13e5 	:	val_out <= 16'h781a;
             14'h13e6 	:	val_out <= 16'h7820;
             14'h13e7 	:	val_out <= 16'h7825;
             14'h13e8 	:	val_out <= 16'h782b;
             14'h13e9 	:	val_out <= 16'h7830;
             14'h13ea 	:	val_out <= 16'h7836;
             14'h13eb 	:	val_out <= 16'h783b;
             14'h13ec 	:	val_out <= 16'h7841;
             14'h13ed 	:	val_out <= 16'h7846;
             14'h13ee 	:	val_out <= 16'h784c;
             14'h13ef 	:	val_out <= 16'h7851;
             14'h13f0 	:	val_out <= 16'h7857;
             14'h13f1 	:	val_out <= 16'h785d;
             14'h13f2 	:	val_out <= 16'h7862;
             14'h13f3 	:	val_out <= 16'h7868;
             14'h13f4 	:	val_out <= 16'h786d;
             14'h13f5 	:	val_out <= 16'h7873;
             14'h13f6 	:	val_out <= 16'h7878;
             14'h13f7 	:	val_out <= 16'h787e;
             14'h13f8 	:	val_out <= 16'h7883;
             14'h13f9 	:	val_out <= 16'h7889;
             14'h13fa 	:	val_out <= 16'h788e;
             14'h13fb 	:	val_out <= 16'h7894;
             14'h13fc 	:	val_out <= 16'h789a;
             14'h13fd 	:	val_out <= 16'h789f;
             14'h13fe 	:	val_out <= 16'h78a5;
             14'h13ff 	:	val_out <= 16'h78aa;
             14'h1400 	:	val_out <= 16'h78b0;
             14'h1401 	:	val_out <= 16'h78b5;
             14'h1402 	:	val_out <= 16'h78bb;
             14'h1403 	:	val_out <= 16'h78c0;
             14'h1404 	:	val_out <= 16'h78c6;
             14'h1405 	:	val_out <= 16'h78cb;
             14'h1406 	:	val_out <= 16'h78d1;
             14'h1407 	:	val_out <= 16'h78d7;
             14'h1408 	:	val_out <= 16'h78dc;
             14'h1409 	:	val_out <= 16'h78e2;
             14'h140a 	:	val_out <= 16'h78e7;
             14'h140b 	:	val_out <= 16'h78ed;
             14'h140c 	:	val_out <= 16'h78f2;
             14'h140d 	:	val_out <= 16'h78f8;
             14'h140e 	:	val_out <= 16'h78fd;
             14'h140f 	:	val_out <= 16'h7903;
             14'h1410 	:	val_out <= 16'h7908;
             14'h1411 	:	val_out <= 16'h790e;
             14'h1412 	:	val_out <= 16'h7913;
             14'h1413 	:	val_out <= 16'h7919;
             14'h1414 	:	val_out <= 16'h791e;
             14'h1415 	:	val_out <= 16'h7924;
             14'h1416 	:	val_out <= 16'h792a;
             14'h1417 	:	val_out <= 16'h792f;
             14'h1418 	:	val_out <= 16'h7935;
             14'h1419 	:	val_out <= 16'h793a;
             14'h141a 	:	val_out <= 16'h7940;
             14'h141b 	:	val_out <= 16'h7945;
             14'h141c 	:	val_out <= 16'h794b;
             14'h141d 	:	val_out <= 16'h7950;
             14'h141e 	:	val_out <= 16'h7956;
             14'h141f 	:	val_out <= 16'h795b;
             14'h1420 	:	val_out <= 16'h7961;
             14'h1421 	:	val_out <= 16'h7966;
             14'h1422 	:	val_out <= 16'h796c;
             14'h1423 	:	val_out <= 16'h7971;
             14'h1424 	:	val_out <= 16'h7977;
             14'h1425 	:	val_out <= 16'h797d;
             14'h1426 	:	val_out <= 16'h7982;
             14'h1427 	:	val_out <= 16'h7988;
             14'h1428 	:	val_out <= 16'h798d;
             14'h1429 	:	val_out <= 16'h7993;
             14'h142a 	:	val_out <= 16'h7998;
             14'h142b 	:	val_out <= 16'h799e;
             14'h142c 	:	val_out <= 16'h79a3;
             14'h142d 	:	val_out <= 16'h79a9;
             14'h142e 	:	val_out <= 16'h79ae;
             14'h142f 	:	val_out <= 16'h79b4;
             14'h1430 	:	val_out <= 16'h79b9;
             14'h1431 	:	val_out <= 16'h79bf;
             14'h1432 	:	val_out <= 16'h79c4;
             14'h1433 	:	val_out <= 16'h79ca;
             14'h1434 	:	val_out <= 16'h79cf;
             14'h1435 	:	val_out <= 16'h79d5;
             14'h1436 	:	val_out <= 16'h79db;
             14'h1437 	:	val_out <= 16'h79e0;
             14'h1438 	:	val_out <= 16'h79e6;
             14'h1439 	:	val_out <= 16'h79eb;
             14'h143a 	:	val_out <= 16'h79f1;
             14'h143b 	:	val_out <= 16'h79f6;
             14'h143c 	:	val_out <= 16'h79fc;
             14'h143d 	:	val_out <= 16'h7a01;
             14'h143e 	:	val_out <= 16'h7a07;
             14'h143f 	:	val_out <= 16'h7a0c;
             14'h1440 	:	val_out <= 16'h7a12;
             14'h1441 	:	val_out <= 16'h7a17;
             14'h1442 	:	val_out <= 16'h7a1d;
             14'h1443 	:	val_out <= 16'h7a22;
             14'h1444 	:	val_out <= 16'h7a28;
             14'h1445 	:	val_out <= 16'h7a2d;
             14'h1446 	:	val_out <= 16'h7a33;
             14'h1447 	:	val_out <= 16'h7a38;
             14'h1448 	:	val_out <= 16'h7a3e;
             14'h1449 	:	val_out <= 16'h7a43;
             14'h144a 	:	val_out <= 16'h7a49;
             14'h144b 	:	val_out <= 16'h7a4f;
             14'h144c 	:	val_out <= 16'h7a54;
             14'h144d 	:	val_out <= 16'h7a5a;
             14'h144e 	:	val_out <= 16'h7a5f;
             14'h144f 	:	val_out <= 16'h7a65;
             14'h1450 	:	val_out <= 16'h7a6a;
             14'h1451 	:	val_out <= 16'h7a70;
             14'h1452 	:	val_out <= 16'h7a75;
             14'h1453 	:	val_out <= 16'h7a7b;
             14'h1454 	:	val_out <= 16'h7a80;
             14'h1455 	:	val_out <= 16'h7a86;
             14'h1456 	:	val_out <= 16'h7a8b;
             14'h1457 	:	val_out <= 16'h7a91;
             14'h1458 	:	val_out <= 16'h7a96;
             14'h1459 	:	val_out <= 16'h7a9c;
             14'h145a 	:	val_out <= 16'h7aa1;
             14'h145b 	:	val_out <= 16'h7aa7;
             14'h145c 	:	val_out <= 16'h7aac;
             14'h145d 	:	val_out <= 16'h7ab2;
             14'h145e 	:	val_out <= 16'h7ab7;
             14'h145f 	:	val_out <= 16'h7abd;
             14'h1460 	:	val_out <= 16'h7ac2;
             14'h1461 	:	val_out <= 16'h7ac8;
             14'h1462 	:	val_out <= 16'h7acd;
             14'h1463 	:	val_out <= 16'h7ad3;
             14'h1464 	:	val_out <= 16'h7ad8;
             14'h1465 	:	val_out <= 16'h7ade;
             14'h1466 	:	val_out <= 16'h7ae3;
             14'h1467 	:	val_out <= 16'h7ae9;
             14'h1468 	:	val_out <= 16'h7aee;
             14'h1469 	:	val_out <= 16'h7af4;
             14'h146a 	:	val_out <= 16'h7af9;
             14'h146b 	:	val_out <= 16'h7aff;
             14'h146c 	:	val_out <= 16'h7b05;
             14'h146d 	:	val_out <= 16'h7b0a;
             14'h146e 	:	val_out <= 16'h7b10;
             14'h146f 	:	val_out <= 16'h7b15;
             14'h1470 	:	val_out <= 16'h7b1b;
             14'h1471 	:	val_out <= 16'h7b20;
             14'h1472 	:	val_out <= 16'h7b26;
             14'h1473 	:	val_out <= 16'h7b2b;
             14'h1474 	:	val_out <= 16'h7b31;
             14'h1475 	:	val_out <= 16'h7b36;
             14'h1476 	:	val_out <= 16'h7b3c;
             14'h1477 	:	val_out <= 16'h7b41;
             14'h1478 	:	val_out <= 16'h7b47;
             14'h1479 	:	val_out <= 16'h7b4c;
             14'h147a 	:	val_out <= 16'h7b52;
             14'h147b 	:	val_out <= 16'h7b57;
             14'h147c 	:	val_out <= 16'h7b5d;
             14'h147d 	:	val_out <= 16'h7b62;
             14'h147e 	:	val_out <= 16'h7b68;
             14'h147f 	:	val_out <= 16'h7b6d;
             14'h1480 	:	val_out <= 16'h7b73;
             14'h1481 	:	val_out <= 16'h7b78;
             14'h1482 	:	val_out <= 16'h7b7e;
             14'h1483 	:	val_out <= 16'h7b83;
             14'h1484 	:	val_out <= 16'h7b89;
             14'h1485 	:	val_out <= 16'h7b8e;
             14'h1486 	:	val_out <= 16'h7b94;
             14'h1487 	:	val_out <= 16'h7b99;
             14'h1488 	:	val_out <= 16'h7b9f;
             14'h1489 	:	val_out <= 16'h7ba4;
             14'h148a 	:	val_out <= 16'h7baa;
             14'h148b 	:	val_out <= 16'h7baf;
             14'h148c 	:	val_out <= 16'h7bb5;
             14'h148d 	:	val_out <= 16'h7bba;
             14'h148e 	:	val_out <= 16'h7bc0;
             14'h148f 	:	val_out <= 16'h7bc5;
             14'h1490 	:	val_out <= 16'h7bcb;
             14'h1491 	:	val_out <= 16'h7bd0;
             14'h1492 	:	val_out <= 16'h7bd6;
             14'h1493 	:	val_out <= 16'h7bdb;
             14'h1494 	:	val_out <= 16'h7be1;
             14'h1495 	:	val_out <= 16'h7be6;
             14'h1496 	:	val_out <= 16'h7bec;
             14'h1497 	:	val_out <= 16'h7bf1;
             14'h1498 	:	val_out <= 16'h7bf7;
             14'h1499 	:	val_out <= 16'h7bfc;
             14'h149a 	:	val_out <= 16'h7c02;
             14'h149b 	:	val_out <= 16'h7c07;
             14'h149c 	:	val_out <= 16'h7c0d;
             14'h149d 	:	val_out <= 16'h7c12;
             14'h149e 	:	val_out <= 16'h7c18;
             14'h149f 	:	val_out <= 16'h7c1d;
             14'h14a0 	:	val_out <= 16'h7c23;
             14'h14a1 	:	val_out <= 16'h7c28;
             14'h14a2 	:	val_out <= 16'h7c2e;
             14'h14a3 	:	val_out <= 16'h7c33;
             14'h14a4 	:	val_out <= 16'h7c39;
             14'h14a5 	:	val_out <= 16'h7c3e;
             14'h14a6 	:	val_out <= 16'h7c44;
             14'h14a7 	:	val_out <= 16'h7c49;
             14'h14a8 	:	val_out <= 16'h7c4f;
             14'h14a9 	:	val_out <= 16'h7c54;
             14'h14aa 	:	val_out <= 16'h7c5a;
             14'h14ab 	:	val_out <= 16'h7c5f;
             14'h14ac 	:	val_out <= 16'h7c65;
             14'h14ad 	:	val_out <= 16'h7c6a;
             14'h14ae 	:	val_out <= 16'h7c70;
             14'h14af 	:	val_out <= 16'h7c75;
             14'h14b0 	:	val_out <= 16'h7c7b;
             14'h14b1 	:	val_out <= 16'h7c80;
             14'h14b2 	:	val_out <= 16'h7c86;
             14'h14b3 	:	val_out <= 16'h7c8b;
             14'h14b4 	:	val_out <= 16'h7c90;
             14'h14b5 	:	val_out <= 16'h7c96;
             14'h14b6 	:	val_out <= 16'h7c9b;
             14'h14b7 	:	val_out <= 16'h7ca1;
             14'h14b8 	:	val_out <= 16'h7ca6;
             14'h14b9 	:	val_out <= 16'h7cac;
             14'h14ba 	:	val_out <= 16'h7cb1;
             14'h14bb 	:	val_out <= 16'h7cb7;
             14'h14bc 	:	val_out <= 16'h7cbc;
             14'h14bd 	:	val_out <= 16'h7cc2;
             14'h14be 	:	val_out <= 16'h7cc7;
             14'h14bf 	:	val_out <= 16'h7ccd;
             14'h14c0 	:	val_out <= 16'h7cd2;
             14'h14c1 	:	val_out <= 16'h7cd8;
             14'h14c2 	:	val_out <= 16'h7cdd;
             14'h14c3 	:	val_out <= 16'h7ce3;
             14'h14c4 	:	val_out <= 16'h7ce8;
             14'h14c5 	:	val_out <= 16'h7cee;
             14'h14c6 	:	val_out <= 16'h7cf3;
             14'h14c7 	:	val_out <= 16'h7cf9;
             14'h14c8 	:	val_out <= 16'h7cfe;
             14'h14c9 	:	val_out <= 16'h7d04;
             14'h14ca 	:	val_out <= 16'h7d09;
             14'h14cb 	:	val_out <= 16'h7d0f;
             14'h14cc 	:	val_out <= 16'h7d14;
             14'h14cd 	:	val_out <= 16'h7d1a;
             14'h14ce 	:	val_out <= 16'h7d1f;
             14'h14cf 	:	val_out <= 16'h7d25;
             14'h14d0 	:	val_out <= 16'h7d2a;
             14'h14d1 	:	val_out <= 16'h7d30;
             14'h14d2 	:	val_out <= 16'h7d35;
             14'h14d3 	:	val_out <= 16'h7d3b;
             14'h14d4 	:	val_out <= 16'h7d40;
             14'h14d5 	:	val_out <= 16'h7d45;
             14'h14d6 	:	val_out <= 16'h7d4b;
             14'h14d7 	:	val_out <= 16'h7d50;
             14'h14d8 	:	val_out <= 16'h7d56;
             14'h14d9 	:	val_out <= 16'h7d5b;
             14'h14da 	:	val_out <= 16'h7d61;
             14'h14db 	:	val_out <= 16'h7d66;
             14'h14dc 	:	val_out <= 16'h7d6c;
             14'h14dd 	:	val_out <= 16'h7d71;
             14'h14de 	:	val_out <= 16'h7d77;
             14'h14df 	:	val_out <= 16'h7d7c;
             14'h14e0 	:	val_out <= 16'h7d82;
             14'h14e1 	:	val_out <= 16'h7d87;
             14'h14e2 	:	val_out <= 16'h7d8d;
             14'h14e3 	:	val_out <= 16'h7d92;
             14'h14e4 	:	val_out <= 16'h7d98;
             14'h14e5 	:	val_out <= 16'h7d9d;
             14'h14e6 	:	val_out <= 16'h7da3;
             14'h14e7 	:	val_out <= 16'h7da8;
             14'h14e8 	:	val_out <= 16'h7dae;
             14'h14e9 	:	val_out <= 16'h7db3;
             14'h14ea 	:	val_out <= 16'h7db8;
             14'h14eb 	:	val_out <= 16'h7dbe;
             14'h14ec 	:	val_out <= 16'h7dc3;
             14'h14ed 	:	val_out <= 16'h7dc9;
             14'h14ee 	:	val_out <= 16'h7dce;
             14'h14ef 	:	val_out <= 16'h7dd4;
             14'h14f0 	:	val_out <= 16'h7dd9;
             14'h14f1 	:	val_out <= 16'h7ddf;
             14'h14f2 	:	val_out <= 16'h7de4;
             14'h14f3 	:	val_out <= 16'h7dea;
             14'h14f4 	:	val_out <= 16'h7def;
             14'h14f5 	:	val_out <= 16'h7df5;
             14'h14f6 	:	val_out <= 16'h7dfa;
             14'h14f7 	:	val_out <= 16'h7e00;
             14'h14f8 	:	val_out <= 16'h7e05;
             14'h14f9 	:	val_out <= 16'h7e0b;
             14'h14fa 	:	val_out <= 16'h7e10;
             14'h14fb 	:	val_out <= 16'h7e15;
             14'h14fc 	:	val_out <= 16'h7e1b;
             14'h14fd 	:	val_out <= 16'h7e20;
             14'h14fe 	:	val_out <= 16'h7e26;
             14'h14ff 	:	val_out <= 16'h7e2b;
             14'h1500 	:	val_out <= 16'h7e31;
             14'h1501 	:	val_out <= 16'h7e36;
             14'h1502 	:	val_out <= 16'h7e3c;
             14'h1503 	:	val_out <= 16'h7e41;
             14'h1504 	:	val_out <= 16'h7e47;
             14'h1505 	:	val_out <= 16'h7e4c;
             14'h1506 	:	val_out <= 16'h7e52;
             14'h1507 	:	val_out <= 16'h7e57;
             14'h1508 	:	val_out <= 16'h7e5d;
             14'h1509 	:	val_out <= 16'h7e62;
             14'h150a 	:	val_out <= 16'h7e67;
             14'h150b 	:	val_out <= 16'h7e6d;
             14'h150c 	:	val_out <= 16'h7e72;
             14'h150d 	:	val_out <= 16'h7e78;
             14'h150e 	:	val_out <= 16'h7e7d;
             14'h150f 	:	val_out <= 16'h7e83;
             14'h1510 	:	val_out <= 16'h7e88;
             14'h1511 	:	val_out <= 16'h7e8e;
             14'h1512 	:	val_out <= 16'h7e93;
             14'h1513 	:	val_out <= 16'h7e99;
             14'h1514 	:	val_out <= 16'h7e9e;
             14'h1515 	:	val_out <= 16'h7ea4;
             14'h1516 	:	val_out <= 16'h7ea9;
             14'h1517 	:	val_out <= 16'h7eae;
             14'h1518 	:	val_out <= 16'h7eb4;
             14'h1519 	:	val_out <= 16'h7eb9;
             14'h151a 	:	val_out <= 16'h7ebf;
             14'h151b 	:	val_out <= 16'h7ec4;
             14'h151c 	:	val_out <= 16'h7eca;
             14'h151d 	:	val_out <= 16'h7ecf;
             14'h151e 	:	val_out <= 16'h7ed5;
             14'h151f 	:	val_out <= 16'h7eda;
             14'h1520 	:	val_out <= 16'h7ee0;
             14'h1521 	:	val_out <= 16'h7ee5;
             14'h1522 	:	val_out <= 16'h7eeb;
             14'h1523 	:	val_out <= 16'h7ef0;
             14'h1524 	:	val_out <= 16'h7ef5;
             14'h1525 	:	val_out <= 16'h7efb;
             14'h1526 	:	val_out <= 16'h7f00;
             14'h1527 	:	val_out <= 16'h7f06;
             14'h1528 	:	val_out <= 16'h7f0b;
             14'h1529 	:	val_out <= 16'h7f11;
             14'h152a 	:	val_out <= 16'h7f16;
             14'h152b 	:	val_out <= 16'h7f1c;
             14'h152c 	:	val_out <= 16'h7f21;
             14'h152d 	:	val_out <= 16'h7f27;
             14'h152e 	:	val_out <= 16'h7f2c;
             14'h152f 	:	val_out <= 16'h7f31;
             14'h1530 	:	val_out <= 16'h7f37;
             14'h1531 	:	val_out <= 16'h7f3c;
             14'h1532 	:	val_out <= 16'h7f42;
             14'h1533 	:	val_out <= 16'h7f47;
             14'h1534 	:	val_out <= 16'h7f4d;
             14'h1535 	:	val_out <= 16'h7f52;
             14'h1536 	:	val_out <= 16'h7f58;
             14'h1537 	:	val_out <= 16'h7f5d;
             14'h1538 	:	val_out <= 16'h7f62;
             14'h1539 	:	val_out <= 16'h7f68;
             14'h153a 	:	val_out <= 16'h7f6d;
             14'h153b 	:	val_out <= 16'h7f73;
             14'h153c 	:	val_out <= 16'h7f78;
             14'h153d 	:	val_out <= 16'h7f7e;
             14'h153e 	:	val_out <= 16'h7f83;
             14'h153f 	:	val_out <= 16'h7f89;
             14'h1540 	:	val_out <= 16'h7f8e;
             14'h1541 	:	val_out <= 16'h7f94;
             14'h1542 	:	val_out <= 16'h7f99;
             14'h1543 	:	val_out <= 16'h7f9e;
             14'h1544 	:	val_out <= 16'h7fa4;
             14'h1545 	:	val_out <= 16'h7fa9;
             14'h1546 	:	val_out <= 16'h7faf;
             14'h1547 	:	val_out <= 16'h7fb4;
             14'h1548 	:	val_out <= 16'h7fba;
             14'h1549 	:	val_out <= 16'h7fbf;
             14'h154a 	:	val_out <= 16'h7fc5;
             14'h154b 	:	val_out <= 16'h7fca;
             14'h154c 	:	val_out <= 16'h7fcf;
             14'h154d 	:	val_out <= 16'h7fd5;
             14'h154e 	:	val_out <= 16'h7fda;
             14'h154f 	:	val_out <= 16'h7fe0;
             14'h1550 	:	val_out <= 16'h7fe5;
             14'h1551 	:	val_out <= 16'h7feb;
             14'h1552 	:	val_out <= 16'h7ff0;
             14'h1553 	:	val_out <= 16'h7ff6;
             14'h1554 	:	val_out <= 16'h7ffb;
             14'h1555 	:	val_out <= 16'h8000;
             14'h1556 	:	val_out <= 16'h8006;
             14'h1557 	:	val_out <= 16'h800b;
             14'h1558 	:	val_out <= 16'h8011;
             14'h1559 	:	val_out <= 16'h8016;
             14'h155a 	:	val_out <= 16'h801c;
             14'h155b 	:	val_out <= 16'h8021;
             14'h155c 	:	val_out <= 16'h8026;
             14'h155d 	:	val_out <= 16'h802c;
             14'h155e 	:	val_out <= 16'h8031;
             14'h155f 	:	val_out <= 16'h8037;
             14'h1560 	:	val_out <= 16'h803c;
             14'h1561 	:	val_out <= 16'h8042;
             14'h1562 	:	val_out <= 16'h8047;
             14'h1563 	:	val_out <= 16'h804d;
             14'h1564 	:	val_out <= 16'h8052;
             14'h1565 	:	val_out <= 16'h8057;
             14'h1566 	:	val_out <= 16'h805d;
             14'h1567 	:	val_out <= 16'h8062;
             14'h1568 	:	val_out <= 16'h8068;
             14'h1569 	:	val_out <= 16'h806d;
             14'h156a 	:	val_out <= 16'h8073;
             14'h156b 	:	val_out <= 16'h8078;
             14'h156c 	:	val_out <= 16'h807d;
             14'h156d 	:	val_out <= 16'h8083;
             14'h156e 	:	val_out <= 16'h8088;
             14'h156f 	:	val_out <= 16'h808e;
             14'h1570 	:	val_out <= 16'h8093;
             14'h1571 	:	val_out <= 16'h8099;
             14'h1572 	:	val_out <= 16'h809e;
             14'h1573 	:	val_out <= 16'h80a4;
             14'h1574 	:	val_out <= 16'h80a9;
             14'h1575 	:	val_out <= 16'h80ae;
             14'h1576 	:	val_out <= 16'h80b4;
             14'h1577 	:	val_out <= 16'h80b9;
             14'h1578 	:	val_out <= 16'h80bf;
             14'h1579 	:	val_out <= 16'h80c4;
             14'h157a 	:	val_out <= 16'h80ca;
             14'h157b 	:	val_out <= 16'h80cf;
             14'h157c 	:	val_out <= 16'h80d4;
             14'h157d 	:	val_out <= 16'h80da;
             14'h157e 	:	val_out <= 16'h80df;
             14'h157f 	:	val_out <= 16'h80e5;
             14'h1580 	:	val_out <= 16'h80ea;
             14'h1581 	:	val_out <= 16'h80f0;
             14'h1582 	:	val_out <= 16'h80f5;
             14'h1583 	:	val_out <= 16'h80fa;
             14'h1584 	:	val_out <= 16'h8100;
             14'h1585 	:	val_out <= 16'h8105;
             14'h1586 	:	val_out <= 16'h810b;
             14'h1587 	:	val_out <= 16'h8110;
             14'h1588 	:	val_out <= 16'h8116;
             14'h1589 	:	val_out <= 16'h811b;
             14'h158a 	:	val_out <= 16'h8120;
             14'h158b 	:	val_out <= 16'h8126;
             14'h158c 	:	val_out <= 16'h812b;
             14'h158d 	:	val_out <= 16'h8131;
             14'h158e 	:	val_out <= 16'h8136;
             14'h158f 	:	val_out <= 16'h813b;
             14'h1590 	:	val_out <= 16'h8141;
             14'h1591 	:	val_out <= 16'h8146;
             14'h1592 	:	val_out <= 16'h814c;
             14'h1593 	:	val_out <= 16'h8151;
             14'h1594 	:	val_out <= 16'h8157;
             14'h1595 	:	val_out <= 16'h815c;
             14'h1596 	:	val_out <= 16'h8161;
             14'h1597 	:	val_out <= 16'h8167;
             14'h1598 	:	val_out <= 16'h816c;
             14'h1599 	:	val_out <= 16'h8172;
             14'h159a 	:	val_out <= 16'h8177;
             14'h159b 	:	val_out <= 16'h817d;
             14'h159c 	:	val_out <= 16'h8182;
             14'h159d 	:	val_out <= 16'h8187;
             14'h159e 	:	val_out <= 16'h818d;
             14'h159f 	:	val_out <= 16'h8192;
             14'h15a0 	:	val_out <= 16'h8198;
             14'h15a1 	:	val_out <= 16'h819d;
             14'h15a2 	:	val_out <= 16'h81a2;
             14'h15a3 	:	val_out <= 16'h81a8;
             14'h15a4 	:	val_out <= 16'h81ad;
             14'h15a5 	:	val_out <= 16'h81b3;
             14'h15a6 	:	val_out <= 16'h81b8;
             14'h15a7 	:	val_out <= 16'h81be;
             14'h15a8 	:	val_out <= 16'h81c3;
             14'h15a9 	:	val_out <= 16'h81c8;
             14'h15aa 	:	val_out <= 16'h81ce;
             14'h15ab 	:	val_out <= 16'h81d3;
             14'h15ac 	:	val_out <= 16'h81d9;
             14'h15ad 	:	val_out <= 16'h81de;
             14'h15ae 	:	val_out <= 16'h81e3;
             14'h15af 	:	val_out <= 16'h81e9;
             14'h15b0 	:	val_out <= 16'h81ee;
             14'h15b1 	:	val_out <= 16'h81f4;
             14'h15b2 	:	val_out <= 16'h81f9;
             14'h15b3 	:	val_out <= 16'h81ff;
             14'h15b4 	:	val_out <= 16'h8204;
             14'h15b5 	:	val_out <= 16'h8209;
             14'h15b6 	:	val_out <= 16'h820f;
             14'h15b7 	:	val_out <= 16'h8214;
             14'h15b8 	:	val_out <= 16'h821a;
             14'h15b9 	:	val_out <= 16'h821f;
             14'h15ba 	:	val_out <= 16'h8224;
             14'h15bb 	:	val_out <= 16'h822a;
             14'h15bc 	:	val_out <= 16'h822f;
             14'h15bd 	:	val_out <= 16'h8235;
             14'h15be 	:	val_out <= 16'h823a;
             14'h15bf 	:	val_out <= 16'h823f;
             14'h15c0 	:	val_out <= 16'h8245;
             14'h15c1 	:	val_out <= 16'h824a;
             14'h15c2 	:	val_out <= 16'h8250;
             14'h15c3 	:	val_out <= 16'h8255;
             14'h15c4 	:	val_out <= 16'h825b;
             14'h15c5 	:	val_out <= 16'h8260;
             14'h15c6 	:	val_out <= 16'h8265;
             14'h15c7 	:	val_out <= 16'h826b;
             14'h15c8 	:	val_out <= 16'h8270;
             14'h15c9 	:	val_out <= 16'h8276;
             14'h15ca 	:	val_out <= 16'h827b;
             14'h15cb 	:	val_out <= 16'h8280;
             14'h15cc 	:	val_out <= 16'h8286;
             14'h15cd 	:	val_out <= 16'h828b;
             14'h15ce 	:	val_out <= 16'h8291;
             14'h15cf 	:	val_out <= 16'h8296;
             14'h15d0 	:	val_out <= 16'h829b;
             14'h15d1 	:	val_out <= 16'h82a1;
             14'h15d2 	:	val_out <= 16'h82a6;
             14'h15d3 	:	val_out <= 16'h82ac;
             14'h15d4 	:	val_out <= 16'h82b1;
             14'h15d5 	:	val_out <= 16'h82b6;
             14'h15d6 	:	val_out <= 16'h82bc;
             14'h15d7 	:	val_out <= 16'h82c1;
             14'h15d8 	:	val_out <= 16'h82c7;
             14'h15d9 	:	val_out <= 16'h82cc;
             14'h15da 	:	val_out <= 16'h82d1;
             14'h15db 	:	val_out <= 16'h82d7;
             14'h15dc 	:	val_out <= 16'h82dc;
             14'h15dd 	:	val_out <= 16'h82e2;
             14'h15de 	:	val_out <= 16'h82e7;
             14'h15df 	:	val_out <= 16'h82ec;
             14'h15e0 	:	val_out <= 16'h82f2;
             14'h15e1 	:	val_out <= 16'h82f7;
             14'h15e2 	:	val_out <= 16'h82fd;
             14'h15e3 	:	val_out <= 16'h8302;
             14'h15e4 	:	val_out <= 16'h8307;
             14'h15e5 	:	val_out <= 16'h830d;
             14'h15e6 	:	val_out <= 16'h8312;
             14'h15e7 	:	val_out <= 16'h8318;
             14'h15e8 	:	val_out <= 16'h831d;
             14'h15e9 	:	val_out <= 16'h8322;
             14'h15ea 	:	val_out <= 16'h8328;
             14'h15eb 	:	val_out <= 16'h832d;
             14'h15ec 	:	val_out <= 16'h8333;
             14'h15ed 	:	val_out <= 16'h8338;
             14'h15ee 	:	val_out <= 16'h833d;
             14'h15ef 	:	val_out <= 16'h8343;
             14'h15f0 	:	val_out <= 16'h8348;
             14'h15f1 	:	val_out <= 16'h834e;
             14'h15f2 	:	val_out <= 16'h8353;
             14'h15f3 	:	val_out <= 16'h8358;
             14'h15f4 	:	val_out <= 16'h835e;
             14'h15f5 	:	val_out <= 16'h8363;
             14'h15f6 	:	val_out <= 16'h8369;
             14'h15f7 	:	val_out <= 16'h836e;
             14'h15f8 	:	val_out <= 16'h8373;
             14'h15f9 	:	val_out <= 16'h8379;
             14'h15fa 	:	val_out <= 16'h837e;
             14'h15fb 	:	val_out <= 16'h8383;
             14'h15fc 	:	val_out <= 16'h8389;
             14'h15fd 	:	val_out <= 16'h838e;
             14'h15fe 	:	val_out <= 16'h8394;
             14'h15ff 	:	val_out <= 16'h8399;
             14'h1600 	:	val_out <= 16'h839e;
             14'h1601 	:	val_out <= 16'h83a4;
             14'h1602 	:	val_out <= 16'h83a9;
             14'h1603 	:	val_out <= 16'h83af;
             14'h1604 	:	val_out <= 16'h83b4;
             14'h1605 	:	val_out <= 16'h83b9;
             14'h1606 	:	val_out <= 16'h83bf;
             14'h1607 	:	val_out <= 16'h83c4;
             14'h1608 	:	val_out <= 16'h83ca;
             14'h1609 	:	val_out <= 16'h83cf;
             14'h160a 	:	val_out <= 16'h83d4;
             14'h160b 	:	val_out <= 16'h83da;
             14'h160c 	:	val_out <= 16'h83df;
             14'h160d 	:	val_out <= 16'h83e4;
             14'h160e 	:	val_out <= 16'h83ea;
             14'h160f 	:	val_out <= 16'h83ef;
             14'h1610 	:	val_out <= 16'h83f5;
             14'h1611 	:	val_out <= 16'h83fa;
             14'h1612 	:	val_out <= 16'h83ff;
             14'h1613 	:	val_out <= 16'h8405;
             14'h1614 	:	val_out <= 16'h840a;
             14'h1615 	:	val_out <= 16'h8410;
             14'h1616 	:	val_out <= 16'h8415;
             14'h1617 	:	val_out <= 16'h841a;
             14'h1618 	:	val_out <= 16'h8420;
             14'h1619 	:	val_out <= 16'h8425;
             14'h161a 	:	val_out <= 16'h842a;
             14'h161b 	:	val_out <= 16'h8430;
             14'h161c 	:	val_out <= 16'h8435;
             14'h161d 	:	val_out <= 16'h843b;
             14'h161e 	:	val_out <= 16'h8440;
             14'h161f 	:	val_out <= 16'h8445;
             14'h1620 	:	val_out <= 16'h844b;
             14'h1621 	:	val_out <= 16'h8450;
             14'h1622 	:	val_out <= 16'h8455;
             14'h1623 	:	val_out <= 16'h845b;
             14'h1624 	:	val_out <= 16'h8460;
             14'h1625 	:	val_out <= 16'h8466;
             14'h1626 	:	val_out <= 16'h846b;
             14'h1627 	:	val_out <= 16'h8470;
             14'h1628 	:	val_out <= 16'h8476;
             14'h1629 	:	val_out <= 16'h847b;
             14'h162a 	:	val_out <= 16'h8481;
             14'h162b 	:	val_out <= 16'h8486;
             14'h162c 	:	val_out <= 16'h848b;
             14'h162d 	:	val_out <= 16'h8491;
             14'h162e 	:	val_out <= 16'h8496;
             14'h162f 	:	val_out <= 16'h849b;
             14'h1630 	:	val_out <= 16'h84a1;
             14'h1631 	:	val_out <= 16'h84a6;
             14'h1632 	:	val_out <= 16'h84ab;
             14'h1633 	:	val_out <= 16'h84b1;
             14'h1634 	:	val_out <= 16'h84b6;
             14'h1635 	:	val_out <= 16'h84bc;
             14'h1636 	:	val_out <= 16'h84c1;
             14'h1637 	:	val_out <= 16'h84c6;
             14'h1638 	:	val_out <= 16'h84cc;
             14'h1639 	:	val_out <= 16'h84d1;
             14'h163a 	:	val_out <= 16'h84d6;
             14'h163b 	:	val_out <= 16'h84dc;
             14'h163c 	:	val_out <= 16'h84e1;
             14'h163d 	:	val_out <= 16'h84e7;
             14'h163e 	:	val_out <= 16'h84ec;
             14'h163f 	:	val_out <= 16'h84f1;
             14'h1640 	:	val_out <= 16'h84f7;
             14'h1641 	:	val_out <= 16'h84fc;
             14'h1642 	:	val_out <= 16'h8501;
             14'h1643 	:	val_out <= 16'h8507;
             14'h1644 	:	val_out <= 16'h850c;
             14'h1645 	:	val_out <= 16'h8512;
             14'h1646 	:	val_out <= 16'h8517;
             14'h1647 	:	val_out <= 16'h851c;
             14'h1648 	:	val_out <= 16'h8522;
             14'h1649 	:	val_out <= 16'h8527;
             14'h164a 	:	val_out <= 16'h852c;
             14'h164b 	:	val_out <= 16'h8532;
             14'h164c 	:	val_out <= 16'h8537;
             14'h164d 	:	val_out <= 16'h853c;
             14'h164e 	:	val_out <= 16'h8542;
             14'h164f 	:	val_out <= 16'h8547;
             14'h1650 	:	val_out <= 16'h854d;
             14'h1651 	:	val_out <= 16'h8552;
             14'h1652 	:	val_out <= 16'h8557;
             14'h1653 	:	val_out <= 16'h855d;
             14'h1654 	:	val_out <= 16'h8562;
             14'h1655 	:	val_out <= 16'h8567;
             14'h1656 	:	val_out <= 16'h856d;
             14'h1657 	:	val_out <= 16'h8572;
             14'h1658 	:	val_out <= 16'h8577;
             14'h1659 	:	val_out <= 16'h857d;
             14'h165a 	:	val_out <= 16'h8582;
             14'h165b 	:	val_out <= 16'h8588;
             14'h165c 	:	val_out <= 16'h858d;
             14'h165d 	:	val_out <= 16'h8592;
             14'h165e 	:	val_out <= 16'h8598;
             14'h165f 	:	val_out <= 16'h859d;
             14'h1660 	:	val_out <= 16'h85a2;
             14'h1661 	:	val_out <= 16'h85a8;
             14'h1662 	:	val_out <= 16'h85ad;
             14'h1663 	:	val_out <= 16'h85b2;
             14'h1664 	:	val_out <= 16'h85b8;
             14'h1665 	:	val_out <= 16'h85bd;
             14'h1666 	:	val_out <= 16'h85c3;
             14'h1667 	:	val_out <= 16'h85c8;
             14'h1668 	:	val_out <= 16'h85cd;
             14'h1669 	:	val_out <= 16'h85d3;
             14'h166a 	:	val_out <= 16'h85d8;
             14'h166b 	:	val_out <= 16'h85dd;
             14'h166c 	:	val_out <= 16'h85e3;
             14'h166d 	:	val_out <= 16'h85e8;
             14'h166e 	:	val_out <= 16'h85ed;
             14'h166f 	:	val_out <= 16'h85f3;
             14'h1670 	:	val_out <= 16'h85f8;
             14'h1671 	:	val_out <= 16'h85fd;
             14'h1672 	:	val_out <= 16'h8603;
             14'h1673 	:	val_out <= 16'h8608;
             14'h1674 	:	val_out <= 16'h860d;
             14'h1675 	:	val_out <= 16'h8613;
             14'h1676 	:	val_out <= 16'h8618;
             14'h1677 	:	val_out <= 16'h861e;
             14'h1678 	:	val_out <= 16'h8623;
             14'h1679 	:	val_out <= 16'h8628;
             14'h167a 	:	val_out <= 16'h862e;
             14'h167b 	:	val_out <= 16'h8633;
             14'h167c 	:	val_out <= 16'h8638;
             14'h167d 	:	val_out <= 16'h863e;
             14'h167e 	:	val_out <= 16'h8643;
             14'h167f 	:	val_out <= 16'h8648;
             14'h1680 	:	val_out <= 16'h864e;
             14'h1681 	:	val_out <= 16'h8653;
             14'h1682 	:	val_out <= 16'h8658;
             14'h1683 	:	val_out <= 16'h865e;
             14'h1684 	:	val_out <= 16'h8663;
             14'h1685 	:	val_out <= 16'h8668;
             14'h1686 	:	val_out <= 16'h866e;
             14'h1687 	:	val_out <= 16'h8673;
             14'h1688 	:	val_out <= 16'h8678;
             14'h1689 	:	val_out <= 16'h867e;
             14'h168a 	:	val_out <= 16'h8683;
             14'h168b 	:	val_out <= 16'h8689;
             14'h168c 	:	val_out <= 16'h868e;
             14'h168d 	:	val_out <= 16'h8693;
             14'h168e 	:	val_out <= 16'h8699;
             14'h168f 	:	val_out <= 16'h869e;
             14'h1690 	:	val_out <= 16'h86a3;
             14'h1691 	:	val_out <= 16'h86a9;
             14'h1692 	:	val_out <= 16'h86ae;
             14'h1693 	:	val_out <= 16'h86b3;
             14'h1694 	:	val_out <= 16'h86b9;
             14'h1695 	:	val_out <= 16'h86be;
             14'h1696 	:	val_out <= 16'h86c3;
             14'h1697 	:	val_out <= 16'h86c9;
             14'h1698 	:	val_out <= 16'h86ce;
             14'h1699 	:	val_out <= 16'h86d3;
             14'h169a 	:	val_out <= 16'h86d9;
             14'h169b 	:	val_out <= 16'h86de;
             14'h169c 	:	val_out <= 16'h86e3;
             14'h169d 	:	val_out <= 16'h86e9;
             14'h169e 	:	val_out <= 16'h86ee;
             14'h169f 	:	val_out <= 16'h86f3;
             14'h16a0 	:	val_out <= 16'h86f9;
             14'h16a1 	:	val_out <= 16'h86fe;
             14'h16a2 	:	val_out <= 16'h8703;
             14'h16a3 	:	val_out <= 16'h8709;
             14'h16a4 	:	val_out <= 16'h870e;
             14'h16a5 	:	val_out <= 16'h8713;
             14'h16a6 	:	val_out <= 16'h8719;
             14'h16a7 	:	val_out <= 16'h871e;
             14'h16a8 	:	val_out <= 16'h8723;
             14'h16a9 	:	val_out <= 16'h8729;
             14'h16aa 	:	val_out <= 16'h872e;
             14'h16ab 	:	val_out <= 16'h8733;
             14'h16ac 	:	val_out <= 16'h8739;
             14'h16ad 	:	val_out <= 16'h873e;
             14'h16ae 	:	val_out <= 16'h8743;
             14'h16af 	:	val_out <= 16'h8749;
             14'h16b0 	:	val_out <= 16'h874e;
             14'h16b1 	:	val_out <= 16'h8753;
             14'h16b2 	:	val_out <= 16'h8759;
             14'h16b3 	:	val_out <= 16'h875e;
             14'h16b4 	:	val_out <= 16'h8763;
             14'h16b5 	:	val_out <= 16'h8769;
             14'h16b6 	:	val_out <= 16'h876e;
             14'h16b7 	:	val_out <= 16'h8773;
             14'h16b8 	:	val_out <= 16'h8779;
             14'h16b9 	:	val_out <= 16'h877e;
             14'h16ba 	:	val_out <= 16'h8783;
             14'h16bb 	:	val_out <= 16'h8789;
             14'h16bc 	:	val_out <= 16'h878e;
             14'h16bd 	:	val_out <= 16'h8793;
             14'h16be 	:	val_out <= 16'h8799;
             14'h16bf 	:	val_out <= 16'h879e;
             14'h16c0 	:	val_out <= 16'h87a3;
             14'h16c1 	:	val_out <= 16'h87a9;
             14'h16c2 	:	val_out <= 16'h87ae;
             14'h16c3 	:	val_out <= 16'h87b3;
             14'h16c4 	:	val_out <= 16'h87b9;
             14'h16c5 	:	val_out <= 16'h87be;
             14'h16c6 	:	val_out <= 16'h87c3;
             14'h16c7 	:	val_out <= 16'h87c9;
             14'h16c8 	:	val_out <= 16'h87ce;
             14'h16c9 	:	val_out <= 16'h87d3;
             14'h16ca 	:	val_out <= 16'h87d9;
             14'h16cb 	:	val_out <= 16'h87de;
             14'h16cc 	:	val_out <= 16'h87e3;
             14'h16cd 	:	val_out <= 16'h87e9;
             14'h16ce 	:	val_out <= 16'h87ee;
             14'h16cf 	:	val_out <= 16'h87f3;
             14'h16d0 	:	val_out <= 16'h87f9;
             14'h16d1 	:	val_out <= 16'h87fe;
             14'h16d2 	:	val_out <= 16'h8803;
             14'h16d3 	:	val_out <= 16'h8809;
             14'h16d4 	:	val_out <= 16'h880e;
             14'h16d5 	:	val_out <= 16'h8813;
             14'h16d6 	:	val_out <= 16'h8819;
             14'h16d7 	:	val_out <= 16'h881e;
             14'h16d8 	:	val_out <= 16'h8823;
             14'h16d9 	:	val_out <= 16'h8828;
             14'h16da 	:	val_out <= 16'h882e;
             14'h16db 	:	val_out <= 16'h8833;
             14'h16dc 	:	val_out <= 16'h8838;
             14'h16dd 	:	val_out <= 16'h883e;
             14'h16de 	:	val_out <= 16'h8843;
             14'h16df 	:	val_out <= 16'h8848;
             14'h16e0 	:	val_out <= 16'h884e;
             14'h16e1 	:	val_out <= 16'h8853;
             14'h16e2 	:	val_out <= 16'h8858;
             14'h16e3 	:	val_out <= 16'h885e;
             14'h16e4 	:	val_out <= 16'h8863;
             14'h16e5 	:	val_out <= 16'h8868;
             14'h16e6 	:	val_out <= 16'h886e;
             14'h16e7 	:	val_out <= 16'h8873;
             14'h16e8 	:	val_out <= 16'h8878;
             14'h16e9 	:	val_out <= 16'h887e;
             14'h16ea 	:	val_out <= 16'h8883;
             14'h16eb 	:	val_out <= 16'h8888;
             14'h16ec 	:	val_out <= 16'h888e;
             14'h16ed 	:	val_out <= 16'h8893;
             14'h16ee 	:	val_out <= 16'h8898;
             14'h16ef 	:	val_out <= 16'h889d;
             14'h16f0 	:	val_out <= 16'h88a3;
             14'h16f1 	:	val_out <= 16'h88a8;
             14'h16f2 	:	val_out <= 16'h88ad;
             14'h16f3 	:	val_out <= 16'h88b3;
             14'h16f4 	:	val_out <= 16'h88b8;
             14'h16f5 	:	val_out <= 16'h88bd;
             14'h16f6 	:	val_out <= 16'h88c3;
             14'h16f7 	:	val_out <= 16'h88c8;
             14'h16f8 	:	val_out <= 16'h88cd;
             14'h16f9 	:	val_out <= 16'h88d3;
             14'h16fa 	:	val_out <= 16'h88d8;
             14'h16fb 	:	val_out <= 16'h88dd;
             14'h16fc 	:	val_out <= 16'h88e3;
             14'h16fd 	:	val_out <= 16'h88e8;
             14'h16fe 	:	val_out <= 16'h88ed;
             14'h16ff 	:	val_out <= 16'h88f2;
             14'h1700 	:	val_out <= 16'h88f8;
             14'h1701 	:	val_out <= 16'h88fd;
             14'h1702 	:	val_out <= 16'h8902;
             14'h1703 	:	val_out <= 16'h8908;
             14'h1704 	:	val_out <= 16'h890d;
             14'h1705 	:	val_out <= 16'h8912;
             14'h1706 	:	val_out <= 16'h8918;
             14'h1707 	:	val_out <= 16'h891d;
             14'h1708 	:	val_out <= 16'h8922;
             14'h1709 	:	val_out <= 16'h8928;
             14'h170a 	:	val_out <= 16'h892d;
             14'h170b 	:	val_out <= 16'h8932;
             14'h170c 	:	val_out <= 16'h8937;
             14'h170d 	:	val_out <= 16'h893d;
             14'h170e 	:	val_out <= 16'h8942;
             14'h170f 	:	val_out <= 16'h8947;
             14'h1710 	:	val_out <= 16'h894d;
             14'h1711 	:	val_out <= 16'h8952;
             14'h1712 	:	val_out <= 16'h8957;
             14'h1713 	:	val_out <= 16'h895d;
             14'h1714 	:	val_out <= 16'h8962;
             14'h1715 	:	val_out <= 16'h8967;
             14'h1716 	:	val_out <= 16'h896c;
             14'h1717 	:	val_out <= 16'h8972;
             14'h1718 	:	val_out <= 16'h8977;
             14'h1719 	:	val_out <= 16'h897c;
             14'h171a 	:	val_out <= 16'h8982;
             14'h171b 	:	val_out <= 16'h8987;
             14'h171c 	:	val_out <= 16'h898c;
             14'h171d 	:	val_out <= 16'h8992;
             14'h171e 	:	val_out <= 16'h8997;
             14'h171f 	:	val_out <= 16'h899c;
             14'h1720 	:	val_out <= 16'h89a1;
             14'h1721 	:	val_out <= 16'h89a7;
             14'h1722 	:	val_out <= 16'h89ac;
             14'h1723 	:	val_out <= 16'h89b1;
             14'h1724 	:	val_out <= 16'h89b7;
             14'h1725 	:	val_out <= 16'h89bc;
             14'h1726 	:	val_out <= 16'h89c1;
             14'h1727 	:	val_out <= 16'h89c7;
             14'h1728 	:	val_out <= 16'h89cc;
             14'h1729 	:	val_out <= 16'h89d1;
             14'h172a 	:	val_out <= 16'h89d6;
             14'h172b 	:	val_out <= 16'h89dc;
             14'h172c 	:	val_out <= 16'h89e1;
             14'h172d 	:	val_out <= 16'h89e6;
             14'h172e 	:	val_out <= 16'h89ec;
             14'h172f 	:	val_out <= 16'h89f1;
             14'h1730 	:	val_out <= 16'h89f6;
             14'h1731 	:	val_out <= 16'h89fb;
             14'h1732 	:	val_out <= 16'h8a01;
             14'h1733 	:	val_out <= 16'h8a06;
             14'h1734 	:	val_out <= 16'h8a0b;
             14'h1735 	:	val_out <= 16'h8a11;
             14'h1736 	:	val_out <= 16'h8a16;
             14'h1737 	:	val_out <= 16'h8a1b;
             14'h1738 	:	val_out <= 16'h8a21;
             14'h1739 	:	val_out <= 16'h8a26;
             14'h173a 	:	val_out <= 16'h8a2b;
             14'h173b 	:	val_out <= 16'h8a30;
             14'h173c 	:	val_out <= 16'h8a36;
             14'h173d 	:	val_out <= 16'h8a3b;
             14'h173e 	:	val_out <= 16'h8a40;
             14'h173f 	:	val_out <= 16'h8a46;
             14'h1740 	:	val_out <= 16'h8a4b;
             14'h1741 	:	val_out <= 16'h8a50;
             14'h1742 	:	val_out <= 16'h8a55;
             14'h1743 	:	val_out <= 16'h8a5b;
             14'h1744 	:	val_out <= 16'h8a60;
             14'h1745 	:	val_out <= 16'h8a65;
             14'h1746 	:	val_out <= 16'h8a6b;
             14'h1747 	:	val_out <= 16'h8a70;
             14'h1748 	:	val_out <= 16'h8a75;
             14'h1749 	:	val_out <= 16'h8a7a;
             14'h174a 	:	val_out <= 16'h8a80;
             14'h174b 	:	val_out <= 16'h8a85;
             14'h174c 	:	val_out <= 16'h8a8a;
             14'h174d 	:	val_out <= 16'h8a90;
             14'h174e 	:	val_out <= 16'h8a95;
             14'h174f 	:	val_out <= 16'h8a9a;
             14'h1750 	:	val_out <= 16'h8a9f;
             14'h1751 	:	val_out <= 16'h8aa5;
             14'h1752 	:	val_out <= 16'h8aaa;
             14'h1753 	:	val_out <= 16'h8aaf;
             14'h1754 	:	val_out <= 16'h8ab5;
             14'h1755 	:	val_out <= 16'h8aba;
             14'h1756 	:	val_out <= 16'h8abf;
             14'h1757 	:	val_out <= 16'h8ac4;
             14'h1758 	:	val_out <= 16'h8aca;
             14'h1759 	:	val_out <= 16'h8acf;
             14'h175a 	:	val_out <= 16'h8ad4;
             14'h175b 	:	val_out <= 16'h8ad9;
             14'h175c 	:	val_out <= 16'h8adf;
             14'h175d 	:	val_out <= 16'h8ae4;
             14'h175e 	:	val_out <= 16'h8ae9;
             14'h175f 	:	val_out <= 16'h8aef;
             14'h1760 	:	val_out <= 16'h8af4;
             14'h1761 	:	val_out <= 16'h8af9;
             14'h1762 	:	val_out <= 16'h8afe;
             14'h1763 	:	val_out <= 16'h8b04;
             14'h1764 	:	val_out <= 16'h8b09;
             14'h1765 	:	val_out <= 16'h8b0e;
             14'h1766 	:	val_out <= 16'h8b14;
             14'h1767 	:	val_out <= 16'h8b19;
             14'h1768 	:	val_out <= 16'h8b1e;
             14'h1769 	:	val_out <= 16'h8b23;
             14'h176a 	:	val_out <= 16'h8b29;
             14'h176b 	:	val_out <= 16'h8b2e;
             14'h176c 	:	val_out <= 16'h8b33;
             14'h176d 	:	val_out <= 16'h8b38;
             14'h176e 	:	val_out <= 16'h8b3e;
             14'h176f 	:	val_out <= 16'h8b43;
             14'h1770 	:	val_out <= 16'h8b48;
             14'h1771 	:	val_out <= 16'h8b4e;
             14'h1772 	:	val_out <= 16'h8b53;
             14'h1773 	:	val_out <= 16'h8b58;
             14'h1774 	:	val_out <= 16'h8b5d;
             14'h1775 	:	val_out <= 16'h8b63;
             14'h1776 	:	val_out <= 16'h8b68;
             14'h1777 	:	val_out <= 16'h8b6d;
             14'h1778 	:	val_out <= 16'h8b72;
             14'h1779 	:	val_out <= 16'h8b78;
             14'h177a 	:	val_out <= 16'h8b7d;
             14'h177b 	:	val_out <= 16'h8b82;
             14'h177c 	:	val_out <= 16'h8b87;
             14'h177d 	:	val_out <= 16'h8b8d;
             14'h177e 	:	val_out <= 16'h8b92;
             14'h177f 	:	val_out <= 16'h8b97;
             14'h1780 	:	val_out <= 16'h8b9d;
             14'h1781 	:	val_out <= 16'h8ba2;
             14'h1782 	:	val_out <= 16'h8ba7;
             14'h1783 	:	val_out <= 16'h8bac;
             14'h1784 	:	val_out <= 16'h8bb2;
             14'h1785 	:	val_out <= 16'h8bb7;
             14'h1786 	:	val_out <= 16'h8bbc;
             14'h1787 	:	val_out <= 16'h8bc1;
             14'h1788 	:	val_out <= 16'h8bc7;
             14'h1789 	:	val_out <= 16'h8bcc;
             14'h178a 	:	val_out <= 16'h8bd1;
             14'h178b 	:	val_out <= 16'h8bd6;
             14'h178c 	:	val_out <= 16'h8bdc;
             14'h178d 	:	val_out <= 16'h8be1;
             14'h178e 	:	val_out <= 16'h8be6;
             14'h178f 	:	val_out <= 16'h8bec;
             14'h1790 	:	val_out <= 16'h8bf1;
             14'h1791 	:	val_out <= 16'h8bf6;
             14'h1792 	:	val_out <= 16'h8bfb;
             14'h1793 	:	val_out <= 16'h8c01;
             14'h1794 	:	val_out <= 16'h8c06;
             14'h1795 	:	val_out <= 16'h8c0b;
             14'h1796 	:	val_out <= 16'h8c10;
             14'h1797 	:	val_out <= 16'h8c16;
             14'h1798 	:	val_out <= 16'h8c1b;
             14'h1799 	:	val_out <= 16'h8c20;
             14'h179a 	:	val_out <= 16'h8c25;
             14'h179b 	:	val_out <= 16'h8c2b;
             14'h179c 	:	val_out <= 16'h8c30;
             14'h179d 	:	val_out <= 16'h8c35;
             14'h179e 	:	val_out <= 16'h8c3a;
             14'h179f 	:	val_out <= 16'h8c40;
             14'h17a0 	:	val_out <= 16'h8c45;
             14'h17a1 	:	val_out <= 16'h8c4a;
             14'h17a2 	:	val_out <= 16'h8c4f;
             14'h17a3 	:	val_out <= 16'h8c55;
             14'h17a4 	:	val_out <= 16'h8c5a;
             14'h17a5 	:	val_out <= 16'h8c5f;
             14'h17a6 	:	val_out <= 16'h8c64;
             14'h17a7 	:	val_out <= 16'h8c6a;
             14'h17a8 	:	val_out <= 16'h8c6f;
             14'h17a9 	:	val_out <= 16'h8c74;
             14'h17aa 	:	val_out <= 16'h8c79;
             14'h17ab 	:	val_out <= 16'h8c7f;
             14'h17ac 	:	val_out <= 16'h8c84;
             14'h17ad 	:	val_out <= 16'h8c89;
             14'h17ae 	:	val_out <= 16'h8c8e;
             14'h17af 	:	val_out <= 16'h8c94;
             14'h17b0 	:	val_out <= 16'h8c99;
             14'h17b1 	:	val_out <= 16'h8c9e;
             14'h17b2 	:	val_out <= 16'h8ca3;
             14'h17b3 	:	val_out <= 16'h8ca9;
             14'h17b4 	:	val_out <= 16'h8cae;
             14'h17b5 	:	val_out <= 16'h8cb3;
             14'h17b6 	:	val_out <= 16'h8cb8;
             14'h17b7 	:	val_out <= 16'h8cbe;
             14'h17b8 	:	val_out <= 16'h8cc3;
             14'h17b9 	:	val_out <= 16'h8cc8;
             14'h17ba 	:	val_out <= 16'h8ccd;
             14'h17bb 	:	val_out <= 16'h8cd3;
             14'h17bc 	:	val_out <= 16'h8cd8;
             14'h17bd 	:	val_out <= 16'h8cdd;
             14'h17be 	:	val_out <= 16'h8ce2;
             14'h17bf 	:	val_out <= 16'h8ce8;
             14'h17c0 	:	val_out <= 16'h8ced;
             14'h17c1 	:	val_out <= 16'h8cf2;
             14'h17c2 	:	val_out <= 16'h8cf7;
             14'h17c3 	:	val_out <= 16'h8cfd;
             14'h17c4 	:	val_out <= 16'h8d02;
             14'h17c5 	:	val_out <= 16'h8d07;
             14'h17c6 	:	val_out <= 16'h8d0c;
             14'h17c7 	:	val_out <= 16'h8d12;
             14'h17c8 	:	val_out <= 16'h8d17;
             14'h17c9 	:	val_out <= 16'h8d1c;
             14'h17ca 	:	val_out <= 16'h8d21;
             14'h17cb 	:	val_out <= 16'h8d27;
             14'h17cc 	:	val_out <= 16'h8d2c;
             14'h17cd 	:	val_out <= 16'h8d31;
             14'h17ce 	:	val_out <= 16'h8d36;
             14'h17cf 	:	val_out <= 16'h8d3c;
             14'h17d0 	:	val_out <= 16'h8d41;
             14'h17d1 	:	val_out <= 16'h8d46;
             14'h17d2 	:	val_out <= 16'h8d4b;
             14'h17d3 	:	val_out <= 16'h8d51;
             14'h17d4 	:	val_out <= 16'h8d56;
             14'h17d5 	:	val_out <= 16'h8d5b;
             14'h17d6 	:	val_out <= 16'h8d60;
             14'h17d7 	:	val_out <= 16'h8d65;
             14'h17d8 	:	val_out <= 16'h8d6b;
             14'h17d9 	:	val_out <= 16'h8d70;
             14'h17da 	:	val_out <= 16'h8d75;
             14'h17db 	:	val_out <= 16'h8d7a;
             14'h17dc 	:	val_out <= 16'h8d80;
             14'h17dd 	:	val_out <= 16'h8d85;
             14'h17de 	:	val_out <= 16'h8d8a;
             14'h17df 	:	val_out <= 16'h8d8f;
             14'h17e0 	:	val_out <= 16'h8d95;
             14'h17e1 	:	val_out <= 16'h8d9a;
             14'h17e2 	:	val_out <= 16'h8d9f;
             14'h17e3 	:	val_out <= 16'h8da4;
             14'h17e4 	:	val_out <= 16'h8daa;
             14'h17e5 	:	val_out <= 16'h8daf;
             14'h17e6 	:	val_out <= 16'h8db4;
             14'h17e7 	:	val_out <= 16'h8db9;
             14'h17e8 	:	val_out <= 16'h8dbe;
             14'h17e9 	:	val_out <= 16'h8dc4;
             14'h17ea 	:	val_out <= 16'h8dc9;
             14'h17eb 	:	val_out <= 16'h8dce;
             14'h17ec 	:	val_out <= 16'h8dd3;
             14'h17ed 	:	val_out <= 16'h8dd9;
             14'h17ee 	:	val_out <= 16'h8dde;
             14'h17ef 	:	val_out <= 16'h8de3;
             14'h17f0 	:	val_out <= 16'h8de8;
             14'h17f1 	:	val_out <= 16'h8dee;
             14'h17f2 	:	val_out <= 16'h8df3;
             14'h17f3 	:	val_out <= 16'h8df8;
             14'h17f4 	:	val_out <= 16'h8dfd;
             14'h17f5 	:	val_out <= 16'h8e02;
             14'h17f6 	:	val_out <= 16'h8e08;
             14'h17f7 	:	val_out <= 16'h8e0d;
             14'h17f8 	:	val_out <= 16'h8e12;
             14'h17f9 	:	val_out <= 16'h8e17;
             14'h17fa 	:	val_out <= 16'h8e1d;
             14'h17fb 	:	val_out <= 16'h8e22;
             14'h17fc 	:	val_out <= 16'h8e27;
             14'h17fd 	:	val_out <= 16'h8e2c;
             14'h17fe 	:	val_out <= 16'h8e32;
             14'h17ff 	:	val_out <= 16'h8e37;
             14'h1800 	:	val_out <= 16'h8e3c;
             14'h1801 	:	val_out <= 16'h8e41;
             14'h1802 	:	val_out <= 16'h8e46;
             14'h1803 	:	val_out <= 16'h8e4c;
             14'h1804 	:	val_out <= 16'h8e51;
             14'h1805 	:	val_out <= 16'h8e56;
             14'h1806 	:	val_out <= 16'h8e5b;
             14'h1807 	:	val_out <= 16'h8e61;
             14'h1808 	:	val_out <= 16'h8e66;
             14'h1809 	:	val_out <= 16'h8e6b;
             14'h180a 	:	val_out <= 16'h8e70;
             14'h180b 	:	val_out <= 16'h8e75;
             14'h180c 	:	val_out <= 16'h8e7b;
             14'h180d 	:	val_out <= 16'h8e80;
             14'h180e 	:	val_out <= 16'h8e85;
             14'h180f 	:	val_out <= 16'h8e8a;
             14'h1810 	:	val_out <= 16'h8e90;
             14'h1811 	:	val_out <= 16'h8e95;
             14'h1812 	:	val_out <= 16'h8e9a;
             14'h1813 	:	val_out <= 16'h8e9f;
             14'h1814 	:	val_out <= 16'h8ea4;
             14'h1815 	:	val_out <= 16'h8eaa;
             14'h1816 	:	val_out <= 16'h8eaf;
             14'h1817 	:	val_out <= 16'h8eb4;
             14'h1818 	:	val_out <= 16'h8eb9;
             14'h1819 	:	val_out <= 16'h8ebe;
             14'h181a 	:	val_out <= 16'h8ec4;
             14'h181b 	:	val_out <= 16'h8ec9;
             14'h181c 	:	val_out <= 16'h8ece;
             14'h181d 	:	val_out <= 16'h8ed3;
             14'h181e 	:	val_out <= 16'h8ed9;
             14'h181f 	:	val_out <= 16'h8ede;
             14'h1820 	:	val_out <= 16'h8ee3;
             14'h1821 	:	val_out <= 16'h8ee8;
             14'h1822 	:	val_out <= 16'h8eed;
             14'h1823 	:	val_out <= 16'h8ef3;
             14'h1824 	:	val_out <= 16'h8ef8;
             14'h1825 	:	val_out <= 16'h8efd;
             14'h1826 	:	val_out <= 16'h8f02;
             14'h1827 	:	val_out <= 16'h8f07;
             14'h1828 	:	val_out <= 16'h8f0d;
             14'h1829 	:	val_out <= 16'h8f12;
             14'h182a 	:	val_out <= 16'h8f17;
             14'h182b 	:	val_out <= 16'h8f1c;
             14'h182c 	:	val_out <= 16'h8f21;
             14'h182d 	:	val_out <= 16'h8f27;
             14'h182e 	:	val_out <= 16'h8f2c;
             14'h182f 	:	val_out <= 16'h8f31;
             14'h1830 	:	val_out <= 16'h8f36;
             14'h1831 	:	val_out <= 16'h8f3c;
             14'h1832 	:	val_out <= 16'h8f41;
             14'h1833 	:	val_out <= 16'h8f46;
             14'h1834 	:	val_out <= 16'h8f4b;
             14'h1835 	:	val_out <= 16'h8f50;
             14'h1836 	:	val_out <= 16'h8f56;
             14'h1837 	:	val_out <= 16'h8f5b;
             14'h1838 	:	val_out <= 16'h8f60;
             14'h1839 	:	val_out <= 16'h8f65;
             14'h183a 	:	val_out <= 16'h8f6a;
             14'h183b 	:	val_out <= 16'h8f70;
             14'h183c 	:	val_out <= 16'h8f75;
             14'h183d 	:	val_out <= 16'h8f7a;
             14'h183e 	:	val_out <= 16'h8f7f;
             14'h183f 	:	val_out <= 16'h8f84;
             14'h1840 	:	val_out <= 16'h8f8a;
             14'h1841 	:	val_out <= 16'h8f8f;
             14'h1842 	:	val_out <= 16'h8f94;
             14'h1843 	:	val_out <= 16'h8f99;
             14'h1844 	:	val_out <= 16'h8f9e;
             14'h1845 	:	val_out <= 16'h8fa4;
             14'h1846 	:	val_out <= 16'h8fa9;
             14'h1847 	:	val_out <= 16'h8fae;
             14'h1848 	:	val_out <= 16'h8fb3;
             14'h1849 	:	val_out <= 16'h8fb8;
             14'h184a 	:	val_out <= 16'h8fbe;
             14'h184b 	:	val_out <= 16'h8fc3;
             14'h184c 	:	val_out <= 16'h8fc8;
             14'h184d 	:	val_out <= 16'h8fcd;
             14'h184e 	:	val_out <= 16'h8fd2;
             14'h184f 	:	val_out <= 16'h8fd8;
             14'h1850 	:	val_out <= 16'h8fdd;
             14'h1851 	:	val_out <= 16'h8fe2;
             14'h1852 	:	val_out <= 16'h8fe7;
             14'h1853 	:	val_out <= 16'h8fec;
             14'h1854 	:	val_out <= 16'h8ff2;
             14'h1855 	:	val_out <= 16'h8ff7;
             14'h1856 	:	val_out <= 16'h8ffc;
             14'h1857 	:	val_out <= 16'h9001;
             14'h1858 	:	val_out <= 16'h9006;
             14'h1859 	:	val_out <= 16'h900c;
             14'h185a 	:	val_out <= 16'h9011;
             14'h185b 	:	val_out <= 16'h9016;
             14'h185c 	:	val_out <= 16'h901b;
             14'h185d 	:	val_out <= 16'h9020;
             14'h185e 	:	val_out <= 16'h9026;
             14'h185f 	:	val_out <= 16'h902b;
             14'h1860 	:	val_out <= 16'h9030;
             14'h1861 	:	val_out <= 16'h9035;
             14'h1862 	:	val_out <= 16'h903a;
             14'h1863 	:	val_out <= 16'h9040;
             14'h1864 	:	val_out <= 16'h9045;
             14'h1865 	:	val_out <= 16'h904a;
             14'h1866 	:	val_out <= 16'h904f;
             14'h1867 	:	val_out <= 16'h9054;
             14'h1868 	:	val_out <= 16'h9059;
             14'h1869 	:	val_out <= 16'h905f;
             14'h186a 	:	val_out <= 16'h9064;
             14'h186b 	:	val_out <= 16'h9069;
             14'h186c 	:	val_out <= 16'h906e;
             14'h186d 	:	val_out <= 16'h9073;
             14'h186e 	:	val_out <= 16'h9079;
             14'h186f 	:	val_out <= 16'h907e;
             14'h1870 	:	val_out <= 16'h9083;
             14'h1871 	:	val_out <= 16'h9088;
             14'h1872 	:	val_out <= 16'h908d;
             14'h1873 	:	val_out <= 16'h9093;
             14'h1874 	:	val_out <= 16'h9098;
             14'h1875 	:	val_out <= 16'h909d;
             14'h1876 	:	val_out <= 16'h90a2;
             14'h1877 	:	val_out <= 16'h90a7;
             14'h1878 	:	val_out <= 16'h90ac;
             14'h1879 	:	val_out <= 16'h90b2;
             14'h187a 	:	val_out <= 16'h90b7;
             14'h187b 	:	val_out <= 16'h90bc;
             14'h187c 	:	val_out <= 16'h90c1;
             14'h187d 	:	val_out <= 16'h90c6;
             14'h187e 	:	val_out <= 16'h90cc;
             14'h187f 	:	val_out <= 16'h90d1;
             14'h1880 	:	val_out <= 16'h90d6;
             14'h1881 	:	val_out <= 16'h90db;
             14'h1882 	:	val_out <= 16'h90e0;
             14'h1883 	:	val_out <= 16'h90e5;
             14'h1884 	:	val_out <= 16'h90eb;
             14'h1885 	:	val_out <= 16'h90f0;
             14'h1886 	:	val_out <= 16'h90f5;
             14'h1887 	:	val_out <= 16'h90fa;
             14'h1888 	:	val_out <= 16'h90ff;
             14'h1889 	:	val_out <= 16'h9105;
             14'h188a 	:	val_out <= 16'h910a;
             14'h188b 	:	val_out <= 16'h910f;
             14'h188c 	:	val_out <= 16'h9114;
             14'h188d 	:	val_out <= 16'h9119;
             14'h188e 	:	val_out <= 16'h911e;
             14'h188f 	:	val_out <= 16'h9124;
             14'h1890 	:	val_out <= 16'h9129;
             14'h1891 	:	val_out <= 16'h912e;
             14'h1892 	:	val_out <= 16'h9133;
             14'h1893 	:	val_out <= 16'h9138;
             14'h1894 	:	val_out <= 16'h913d;
             14'h1895 	:	val_out <= 16'h9143;
             14'h1896 	:	val_out <= 16'h9148;
             14'h1897 	:	val_out <= 16'h914d;
             14'h1898 	:	val_out <= 16'h9152;
             14'h1899 	:	val_out <= 16'h9157;
             14'h189a 	:	val_out <= 16'h915c;
             14'h189b 	:	val_out <= 16'h9162;
             14'h189c 	:	val_out <= 16'h9167;
             14'h189d 	:	val_out <= 16'h916c;
             14'h189e 	:	val_out <= 16'h9171;
             14'h189f 	:	val_out <= 16'h9176;
             14'h18a0 	:	val_out <= 16'h917c;
             14'h18a1 	:	val_out <= 16'h9181;
             14'h18a2 	:	val_out <= 16'h9186;
             14'h18a3 	:	val_out <= 16'h918b;
             14'h18a4 	:	val_out <= 16'h9190;
             14'h18a5 	:	val_out <= 16'h9195;
             14'h18a6 	:	val_out <= 16'h919b;
             14'h18a7 	:	val_out <= 16'h91a0;
             14'h18a8 	:	val_out <= 16'h91a5;
             14'h18a9 	:	val_out <= 16'h91aa;
             14'h18aa 	:	val_out <= 16'h91af;
             14'h18ab 	:	val_out <= 16'h91b4;
             14'h18ac 	:	val_out <= 16'h91ba;
             14'h18ad 	:	val_out <= 16'h91bf;
             14'h18ae 	:	val_out <= 16'h91c4;
             14'h18af 	:	val_out <= 16'h91c9;
             14'h18b0 	:	val_out <= 16'h91ce;
             14'h18b1 	:	val_out <= 16'h91d3;
             14'h18b2 	:	val_out <= 16'h91d9;
             14'h18b3 	:	val_out <= 16'h91de;
             14'h18b4 	:	val_out <= 16'h91e3;
             14'h18b5 	:	val_out <= 16'h91e8;
             14'h18b6 	:	val_out <= 16'h91ed;
             14'h18b7 	:	val_out <= 16'h91f2;
             14'h18b8 	:	val_out <= 16'h91f7;
             14'h18b9 	:	val_out <= 16'h91fd;
             14'h18ba 	:	val_out <= 16'h9202;
             14'h18bb 	:	val_out <= 16'h9207;
             14'h18bc 	:	val_out <= 16'h920c;
             14'h18bd 	:	val_out <= 16'h9211;
             14'h18be 	:	val_out <= 16'h9216;
             14'h18bf 	:	val_out <= 16'h921c;
             14'h18c0 	:	val_out <= 16'h9221;
             14'h18c1 	:	val_out <= 16'h9226;
             14'h18c2 	:	val_out <= 16'h922b;
             14'h18c3 	:	val_out <= 16'h9230;
             14'h18c4 	:	val_out <= 16'h9235;
             14'h18c5 	:	val_out <= 16'h923b;
             14'h18c6 	:	val_out <= 16'h9240;
             14'h18c7 	:	val_out <= 16'h9245;
             14'h18c8 	:	val_out <= 16'h924a;
             14'h18c9 	:	val_out <= 16'h924f;
             14'h18ca 	:	val_out <= 16'h9254;
             14'h18cb 	:	val_out <= 16'h9259;
             14'h18cc 	:	val_out <= 16'h925f;
             14'h18cd 	:	val_out <= 16'h9264;
             14'h18ce 	:	val_out <= 16'h9269;
             14'h18cf 	:	val_out <= 16'h926e;
             14'h18d0 	:	val_out <= 16'h9273;
             14'h18d1 	:	val_out <= 16'h9278;
             14'h18d2 	:	val_out <= 16'h927e;
             14'h18d3 	:	val_out <= 16'h9283;
             14'h18d4 	:	val_out <= 16'h9288;
             14'h18d5 	:	val_out <= 16'h928d;
             14'h18d6 	:	val_out <= 16'h9292;
             14'h18d7 	:	val_out <= 16'h9297;
             14'h18d8 	:	val_out <= 16'h929c;
             14'h18d9 	:	val_out <= 16'h92a2;
             14'h18da 	:	val_out <= 16'h92a7;
             14'h18db 	:	val_out <= 16'h92ac;
             14'h18dc 	:	val_out <= 16'h92b1;
             14'h18dd 	:	val_out <= 16'h92b6;
             14'h18de 	:	val_out <= 16'h92bb;
             14'h18df 	:	val_out <= 16'h92c1;
             14'h18e0 	:	val_out <= 16'h92c6;
             14'h18e1 	:	val_out <= 16'h92cb;
             14'h18e2 	:	val_out <= 16'h92d0;
             14'h18e3 	:	val_out <= 16'h92d5;
             14'h18e4 	:	val_out <= 16'h92da;
             14'h18e5 	:	val_out <= 16'h92df;
             14'h18e6 	:	val_out <= 16'h92e5;
             14'h18e7 	:	val_out <= 16'h92ea;
             14'h18e8 	:	val_out <= 16'h92ef;
             14'h18e9 	:	val_out <= 16'h92f4;
             14'h18ea 	:	val_out <= 16'h92f9;
             14'h18eb 	:	val_out <= 16'h92fe;
             14'h18ec 	:	val_out <= 16'h9303;
             14'h18ed 	:	val_out <= 16'h9309;
             14'h18ee 	:	val_out <= 16'h930e;
             14'h18ef 	:	val_out <= 16'h9313;
             14'h18f0 	:	val_out <= 16'h9318;
             14'h18f1 	:	val_out <= 16'h931d;
             14'h18f2 	:	val_out <= 16'h9322;
             14'h18f3 	:	val_out <= 16'h9327;
             14'h18f4 	:	val_out <= 16'h932d;
             14'h18f5 	:	val_out <= 16'h9332;
             14'h18f6 	:	val_out <= 16'h9337;
             14'h18f7 	:	val_out <= 16'h933c;
             14'h18f8 	:	val_out <= 16'h9341;
             14'h18f9 	:	val_out <= 16'h9346;
             14'h18fa 	:	val_out <= 16'h934b;
             14'h18fb 	:	val_out <= 16'h9351;
             14'h18fc 	:	val_out <= 16'h9356;
             14'h18fd 	:	val_out <= 16'h935b;
             14'h18fe 	:	val_out <= 16'h9360;
             14'h18ff 	:	val_out <= 16'h9365;
             14'h1900 	:	val_out <= 16'h936a;
             14'h1901 	:	val_out <= 16'h936f;
             14'h1902 	:	val_out <= 16'h9375;
             14'h1903 	:	val_out <= 16'h937a;
             14'h1904 	:	val_out <= 16'h937f;
             14'h1905 	:	val_out <= 16'h9384;
             14'h1906 	:	val_out <= 16'h9389;
             14'h1907 	:	val_out <= 16'h938e;
             14'h1908 	:	val_out <= 16'h9393;
             14'h1909 	:	val_out <= 16'h9398;
             14'h190a 	:	val_out <= 16'h939e;
             14'h190b 	:	val_out <= 16'h93a3;
             14'h190c 	:	val_out <= 16'h93a8;
             14'h190d 	:	val_out <= 16'h93ad;
             14'h190e 	:	val_out <= 16'h93b2;
             14'h190f 	:	val_out <= 16'h93b7;
             14'h1910 	:	val_out <= 16'h93bc;
             14'h1911 	:	val_out <= 16'h93c2;
             14'h1912 	:	val_out <= 16'h93c7;
             14'h1913 	:	val_out <= 16'h93cc;
             14'h1914 	:	val_out <= 16'h93d1;
             14'h1915 	:	val_out <= 16'h93d6;
             14'h1916 	:	val_out <= 16'h93db;
             14'h1917 	:	val_out <= 16'h93e0;
             14'h1918 	:	val_out <= 16'h93e5;
             14'h1919 	:	val_out <= 16'h93eb;
             14'h191a 	:	val_out <= 16'h93f0;
             14'h191b 	:	val_out <= 16'h93f5;
             14'h191c 	:	val_out <= 16'h93fa;
             14'h191d 	:	val_out <= 16'h93ff;
             14'h191e 	:	val_out <= 16'h9404;
             14'h191f 	:	val_out <= 16'h9409;
             14'h1920 	:	val_out <= 16'h940e;
             14'h1921 	:	val_out <= 16'h9414;
             14'h1922 	:	val_out <= 16'h9419;
             14'h1923 	:	val_out <= 16'h941e;
             14'h1924 	:	val_out <= 16'h9423;
             14'h1925 	:	val_out <= 16'h9428;
             14'h1926 	:	val_out <= 16'h942d;
             14'h1927 	:	val_out <= 16'h9432;
             14'h1928 	:	val_out <= 16'h9437;
             14'h1929 	:	val_out <= 16'h943d;
             14'h192a 	:	val_out <= 16'h9442;
             14'h192b 	:	val_out <= 16'h9447;
             14'h192c 	:	val_out <= 16'h944c;
             14'h192d 	:	val_out <= 16'h9451;
             14'h192e 	:	val_out <= 16'h9456;
             14'h192f 	:	val_out <= 16'h945b;
             14'h1930 	:	val_out <= 16'h9460;
             14'h1931 	:	val_out <= 16'h9466;
             14'h1932 	:	val_out <= 16'h946b;
             14'h1933 	:	val_out <= 16'h9470;
             14'h1934 	:	val_out <= 16'h9475;
             14'h1935 	:	val_out <= 16'h947a;
             14'h1936 	:	val_out <= 16'h947f;
             14'h1937 	:	val_out <= 16'h9484;
             14'h1938 	:	val_out <= 16'h9489;
             14'h1939 	:	val_out <= 16'h948e;
             14'h193a 	:	val_out <= 16'h9494;
             14'h193b 	:	val_out <= 16'h9499;
             14'h193c 	:	val_out <= 16'h949e;
             14'h193d 	:	val_out <= 16'h94a3;
             14'h193e 	:	val_out <= 16'h94a8;
             14'h193f 	:	val_out <= 16'h94ad;
             14'h1940 	:	val_out <= 16'h94b2;
             14'h1941 	:	val_out <= 16'h94b7;
             14'h1942 	:	val_out <= 16'h94bd;
             14'h1943 	:	val_out <= 16'h94c2;
             14'h1944 	:	val_out <= 16'h94c7;
             14'h1945 	:	val_out <= 16'h94cc;
             14'h1946 	:	val_out <= 16'h94d1;
             14'h1947 	:	val_out <= 16'h94d6;
             14'h1948 	:	val_out <= 16'h94db;
             14'h1949 	:	val_out <= 16'h94e0;
             14'h194a 	:	val_out <= 16'h94e5;
             14'h194b 	:	val_out <= 16'h94eb;
             14'h194c 	:	val_out <= 16'h94f0;
             14'h194d 	:	val_out <= 16'h94f5;
             14'h194e 	:	val_out <= 16'h94fa;
             14'h194f 	:	val_out <= 16'h94ff;
             14'h1950 	:	val_out <= 16'h9504;
             14'h1951 	:	val_out <= 16'h9509;
             14'h1952 	:	val_out <= 16'h950e;
             14'h1953 	:	val_out <= 16'h9513;
             14'h1954 	:	val_out <= 16'h9519;
             14'h1955 	:	val_out <= 16'h951e;
             14'h1956 	:	val_out <= 16'h9523;
             14'h1957 	:	val_out <= 16'h9528;
             14'h1958 	:	val_out <= 16'h952d;
             14'h1959 	:	val_out <= 16'h9532;
             14'h195a 	:	val_out <= 16'h9537;
             14'h195b 	:	val_out <= 16'h953c;
             14'h195c 	:	val_out <= 16'h9541;
             14'h195d 	:	val_out <= 16'h9546;
             14'h195e 	:	val_out <= 16'h954c;
             14'h195f 	:	val_out <= 16'h9551;
             14'h1960 	:	val_out <= 16'h9556;
             14'h1961 	:	val_out <= 16'h955b;
             14'h1962 	:	val_out <= 16'h9560;
             14'h1963 	:	val_out <= 16'h9565;
             14'h1964 	:	val_out <= 16'h956a;
             14'h1965 	:	val_out <= 16'h956f;
             14'h1966 	:	val_out <= 16'h9574;
             14'h1967 	:	val_out <= 16'h9579;
             14'h1968 	:	val_out <= 16'h957f;
             14'h1969 	:	val_out <= 16'h9584;
             14'h196a 	:	val_out <= 16'h9589;
             14'h196b 	:	val_out <= 16'h958e;
             14'h196c 	:	val_out <= 16'h9593;
             14'h196d 	:	val_out <= 16'h9598;
             14'h196e 	:	val_out <= 16'h959d;
             14'h196f 	:	val_out <= 16'h95a2;
             14'h1970 	:	val_out <= 16'h95a7;
             14'h1971 	:	val_out <= 16'h95ac;
             14'h1972 	:	val_out <= 16'h95b2;
             14'h1973 	:	val_out <= 16'h95b7;
             14'h1974 	:	val_out <= 16'h95bc;
             14'h1975 	:	val_out <= 16'h95c1;
             14'h1976 	:	val_out <= 16'h95c6;
             14'h1977 	:	val_out <= 16'h95cb;
             14'h1978 	:	val_out <= 16'h95d0;
             14'h1979 	:	val_out <= 16'h95d5;
             14'h197a 	:	val_out <= 16'h95da;
             14'h197b 	:	val_out <= 16'h95df;
             14'h197c 	:	val_out <= 16'h95e5;
             14'h197d 	:	val_out <= 16'h95ea;
             14'h197e 	:	val_out <= 16'h95ef;
             14'h197f 	:	val_out <= 16'h95f4;
             14'h1980 	:	val_out <= 16'h95f9;
             14'h1981 	:	val_out <= 16'h95fe;
             14'h1982 	:	val_out <= 16'h9603;
             14'h1983 	:	val_out <= 16'h9608;
             14'h1984 	:	val_out <= 16'h960d;
             14'h1985 	:	val_out <= 16'h9612;
             14'h1986 	:	val_out <= 16'h9617;
             14'h1987 	:	val_out <= 16'h961d;
             14'h1988 	:	val_out <= 16'h9622;
             14'h1989 	:	val_out <= 16'h9627;
             14'h198a 	:	val_out <= 16'h962c;
             14'h198b 	:	val_out <= 16'h9631;
             14'h198c 	:	val_out <= 16'h9636;
             14'h198d 	:	val_out <= 16'h963b;
             14'h198e 	:	val_out <= 16'h9640;
             14'h198f 	:	val_out <= 16'h9645;
             14'h1990 	:	val_out <= 16'h964a;
             14'h1991 	:	val_out <= 16'h964f;
             14'h1992 	:	val_out <= 16'h9654;
             14'h1993 	:	val_out <= 16'h965a;
             14'h1994 	:	val_out <= 16'h965f;
             14'h1995 	:	val_out <= 16'h9664;
             14'h1996 	:	val_out <= 16'h9669;
             14'h1997 	:	val_out <= 16'h966e;
             14'h1998 	:	val_out <= 16'h9673;
             14'h1999 	:	val_out <= 16'h9678;
             14'h199a 	:	val_out <= 16'h967d;
             14'h199b 	:	val_out <= 16'h9682;
             14'h199c 	:	val_out <= 16'h9687;
             14'h199d 	:	val_out <= 16'h968c;
             14'h199e 	:	val_out <= 16'h9691;
             14'h199f 	:	val_out <= 16'h9697;
             14'h19a0 	:	val_out <= 16'h969c;
             14'h19a1 	:	val_out <= 16'h96a1;
             14'h19a2 	:	val_out <= 16'h96a6;
             14'h19a3 	:	val_out <= 16'h96ab;
             14'h19a4 	:	val_out <= 16'h96b0;
             14'h19a5 	:	val_out <= 16'h96b5;
             14'h19a6 	:	val_out <= 16'h96ba;
             14'h19a7 	:	val_out <= 16'h96bf;
             14'h19a8 	:	val_out <= 16'h96c4;
             14'h19a9 	:	val_out <= 16'h96c9;
             14'h19aa 	:	val_out <= 16'h96ce;
             14'h19ab 	:	val_out <= 16'h96d4;
             14'h19ac 	:	val_out <= 16'h96d9;
             14'h19ad 	:	val_out <= 16'h96de;
             14'h19ae 	:	val_out <= 16'h96e3;
             14'h19af 	:	val_out <= 16'h96e8;
             14'h19b0 	:	val_out <= 16'h96ed;
             14'h19b1 	:	val_out <= 16'h96f2;
             14'h19b2 	:	val_out <= 16'h96f7;
             14'h19b3 	:	val_out <= 16'h96fc;
             14'h19b4 	:	val_out <= 16'h9701;
             14'h19b5 	:	val_out <= 16'h9706;
             14'h19b6 	:	val_out <= 16'h970b;
             14'h19b7 	:	val_out <= 16'h9710;
             14'h19b8 	:	val_out <= 16'h9715;
             14'h19b9 	:	val_out <= 16'h971b;
             14'h19ba 	:	val_out <= 16'h9720;
             14'h19bb 	:	val_out <= 16'h9725;
             14'h19bc 	:	val_out <= 16'h972a;
             14'h19bd 	:	val_out <= 16'h972f;
             14'h19be 	:	val_out <= 16'h9734;
             14'h19bf 	:	val_out <= 16'h9739;
             14'h19c0 	:	val_out <= 16'h973e;
             14'h19c1 	:	val_out <= 16'h9743;
             14'h19c2 	:	val_out <= 16'h9748;
             14'h19c3 	:	val_out <= 16'h974d;
             14'h19c4 	:	val_out <= 16'h9752;
             14'h19c5 	:	val_out <= 16'h9757;
             14'h19c6 	:	val_out <= 16'h975c;
             14'h19c7 	:	val_out <= 16'h9762;
             14'h19c8 	:	val_out <= 16'h9767;
             14'h19c9 	:	val_out <= 16'h976c;
             14'h19ca 	:	val_out <= 16'h9771;
             14'h19cb 	:	val_out <= 16'h9776;
             14'h19cc 	:	val_out <= 16'h977b;
             14'h19cd 	:	val_out <= 16'h9780;
             14'h19ce 	:	val_out <= 16'h9785;
             14'h19cf 	:	val_out <= 16'h978a;
             14'h19d0 	:	val_out <= 16'h978f;
             14'h19d1 	:	val_out <= 16'h9794;
             14'h19d2 	:	val_out <= 16'h9799;
             14'h19d3 	:	val_out <= 16'h979e;
             14'h19d4 	:	val_out <= 16'h97a3;
             14'h19d5 	:	val_out <= 16'h97a8;
             14'h19d6 	:	val_out <= 16'h97ae;
             14'h19d7 	:	val_out <= 16'h97b3;
             14'h19d8 	:	val_out <= 16'h97b8;
             14'h19d9 	:	val_out <= 16'h97bd;
             14'h19da 	:	val_out <= 16'h97c2;
             14'h19db 	:	val_out <= 16'h97c7;
             14'h19dc 	:	val_out <= 16'h97cc;
             14'h19dd 	:	val_out <= 16'h97d1;
             14'h19de 	:	val_out <= 16'h97d6;
             14'h19df 	:	val_out <= 16'h97db;
             14'h19e0 	:	val_out <= 16'h97e0;
             14'h19e1 	:	val_out <= 16'h97e5;
             14'h19e2 	:	val_out <= 16'h97ea;
             14'h19e3 	:	val_out <= 16'h97ef;
             14'h19e4 	:	val_out <= 16'h97f4;
             14'h19e5 	:	val_out <= 16'h97f9;
             14'h19e6 	:	val_out <= 16'h97fe;
             14'h19e7 	:	val_out <= 16'h9803;
             14'h19e8 	:	val_out <= 16'h9809;
             14'h19e9 	:	val_out <= 16'h980e;
             14'h19ea 	:	val_out <= 16'h9813;
             14'h19eb 	:	val_out <= 16'h9818;
             14'h19ec 	:	val_out <= 16'h981d;
             14'h19ed 	:	val_out <= 16'h9822;
             14'h19ee 	:	val_out <= 16'h9827;
             14'h19ef 	:	val_out <= 16'h982c;
             14'h19f0 	:	val_out <= 16'h9831;
             14'h19f1 	:	val_out <= 16'h9836;
             14'h19f2 	:	val_out <= 16'h983b;
             14'h19f3 	:	val_out <= 16'h9840;
             14'h19f4 	:	val_out <= 16'h9845;
             14'h19f5 	:	val_out <= 16'h984a;
             14'h19f6 	:	val_out <= 16'h984f;
             14'h19f7 	:	val_out <= 16'h9854;
             14'h19f8 	:	val_out <= 16'h9859;
             14'h19f9 	:	val_out <= 16'h985e;
             14'h19fa 	:	val_out <= 16'h9863;
             14'h19fb 	:	val_out <= 16'h9869;
             14'h19fc 	:	val_out <= 16'h986e;
             14'h19fd 	:	val_out <= 16'h9873;
             14'h19fe 	:	val_out <= 16'h9878;
             14'h19ff 	:	val_out <= 16'h987d;
             14'h1a00 	:	val_out <= 16'h9882;
             14'h1a01 	:	val_out <= 16'h9887;
             14'h1a02 	:	val_out <= 16'h988c;
             14'h1a03 	:	val_out <= 16'h9891;
             14'h1a04 	:	val_out <= 16'h9896;
             14'h1a05 	:	val_out <= 16'h989b;
             14'h1a06 	:	val_out <= 16'h98a0;
             14'h1a07 	:	val_out <= 16'h98a5;
             14'h1a08 	:	val_out <= 16'h98aa;
             14'h1a09 	:	val_out <= 16'h98af;
             14'h1a0a 	:	val_out <= 16'h98b4;
             14'h1a0b 	:	val_out <= 16'h98b9;
             14'h1a0c 	:	val_out <= 16'h98be;
             14'h1a0d 	:	val_out <= 16'h98c3;
             14'h1a0e 	:	val_out <= 16'h98c8;
             14'h1a0f 	:	val_out <= 16'h98cd;
             14'h1a10 	:	val_out <= 16'h98d2;
             14'h1a11 	:	val_out <= 16'h98d8;
             14'h1a12 	:	val_out <= 16'h98dd;
             14'h1a13 	:	val_out <= 16'h98e2;
             14'h1a14 	:	val_out <= 16'h98e7;
             14'h1a15 	:	val_out <= 16'h98ec;
             14'h1a16 	:	val_out <= 16'h98f1;
             14'h1a17 	:	val_out <= 16'h98f6;
             14'h1a18 	:	val_out <= 16'h98fb;
             14'h1a19 	:	val_out <= 16'h9900;
             14'h1a1a 	:	val_out <= 16'h9905;
             14'h1a1b 	:	val_out <= 16'h990a;
             14'h1a1c 	:	val_out <= 16'h990f;
             14'h1a1d 	:	val_out <= 16'h9914;
             14'h1a1e 	:	val_out <= 16'h9919;
             14'h1a1f 	:	val_out <= 16'h991e;
             14'h1a20 	:	val_out <= 16'h9923;
             14'h1a21 	:	val_out <= 16'h9928;
             14'h1a22 	:	val_out <= 16'h992d;
             14'h1a23 	:	val_out <= 16'h9932;
             14'h1a24 	:	val_out <= 16'h9937;
             14'h1a25 	:	val_out <= 16'h993c;
             14'h1a26 	:	val_out <= 16'h9941;
             14'h1a27 	:	val_out <= 16'h9946;
             14'h1a28 	:	val_out <= 16'h994b;
             14'h1a29 	:	val_out <= 16'h9950;
             14'h1a2a 	:	val_out <= 16'h9955;
             14'h1a2b 	:	val_out <= 16'h995a;
             14'h1a2c 	:	val_out <= 16'h995f;
             14'h1a2d 	:	val_out <= 16'h9965;
             14'h1a2e 	:	val_out <= 16'h996a;
             14'h1a2f 	:	val_out <= 16'h996f;
             14'h1a30 	:	val_out <= 16'h9974;
             14'h1a31 	:	val_out <= 16'h9979;
             14'h1a32 	:	val_out <= 16'h997e;
             14'h1a33 	:	val_out <= 16'h9983;
             14'h1a34 	:	val_out <= 16'h9988;
             14'h1a35 	:	val_out <= 16'h998d;
             14'h1a36 	:	val_out <= 16'h9992;
             14'h1a37 	:	val_out <= 16'h9997;
             14'h1a38 	:	val_out <= 16'h999c;
             14'h1a39 	:	val_out <= 16'h99a1;
             14'h1a3a 	:	val_out <= 16'h99a6;
             14'h1a3b 	:	val_out <= 16'h99ab;
             14'h1a3c 	:	val_out <= 16'h99b0;
             14'h1a3d 	:	val_out <= 16'h99b5;
             14'h1a3e 	:	val_out <= 16'h99ba;
             14'h1a3f 	:	val_out <= 16'h99bf;
             14'h1a40 	:	val_out <= 16'h99c4;
             14'h1a41 	:	val_out <= 16'h99c9;
             14'h1a42 	:	val_out <= 16'h99ce;
             14'h1a43 	:	val_out <= 16'h99d3;
             14'h1a44 	:	val_out <= 16'h99d8;
             14'h1a45 	:	val_out <= 16'h99dd;
             14'h1a46 	:	val_out <= 16'h99e2;
             14'h1a47 	:	val_out <= 16'h99e7;
             14'h1a48 	:	val_out <= 16'h99ec;
             14'h1a49 	:	val_out <= 16'h99f1;
             14'h1a4a 	:	val_out <= 16'h99f6;
             14'h1a4b 	:	val_out <= 16'h99fb;
             14'h1a4c 	:	val_out <= 16'h9a00;
             14'h1a4d 	:	val_out <= 16'h9a05;
             14'h1a4e 	:	val_out <= 16'h9a0a;
             14'h1a4f 	:	val_out <= 16'h9a0f;
             14'h1a50 	:	val_out <= 16'h9a14;
             14'h1a51 	:	val_out <= 16'h9a19;
             14'h1a52 	:	val_out <= 16'h9a1e;
             14'h1a53 	:	val_out <= 16'h9a23;
             14'h1a54 	:	val_out <= 16'h9a28;
             14'h1a55 	:	val_out <= 16'h9a2d;
             14'h1a56 	:	val_out <= 16'h9a32;
             14'h1a57 	:	val_out <= 16'h9a37;
             14'h1a58 	:	val_out <= 16'h9a3c;
             14'h1a59 	:	val_out <= 16'h9a41;
             14'h1a5a 	:	val_out <= 16'h9a47;
             14'h1a5b 	:	val_out <= 16'h9a4c;
             14'h1a5c 	:	val_out <= 16'h9a51;
             14'h1a5d 	:	val_out <= 16'h9a56;
             14'h1a5e 	:	val_out <= 16'h9a5b;
             14'h1a5f 	:	val_out <= 16'h9a60;
             14'h1a60 	:	val_out <= 16'h9a65;
             14'h1a61 	:	val_out <= 16'h9a6a;
             14'h1a62 	:	val_out <= 16'h9a6f;
             14'h1a63 	:	val_out <= 16'h9a74;
             14'h1a64 	:	val_out <= 16'h9a79;
             14'h1a65 	:	val_out <= 16'h9a7e;
             14'h1a66 	:	val_out <= 16'h9a83;
             14'h1a67 	:	val_out <= 16'h9a88;
             14'h1a68 	:	val_out <= 16'h9a8d;
             14'h1a69 	:	val_out <= 16'h9a92;
             14'h1a6a 	:	val_out <= 16'h9a97;
             14'h1a6b 	:	val_out <= 16'h9a9c;
             14'h1a6c 	:	val_out <= 16'h9aa1;
             14'h1a6d 	:	val_out <= 16'h9aa6;
             14'h1a6e 	:	val_out <= 16'h9aab;
             14'h1a6f 	:	val_out <= 16'h9ab0;
             14'h1a70 	:	val_out <= 16'h9ab5;
             14'h1a71 	:	val_out <= 16'h9aba;
             14'h1a72 	:	val_out <= 16'h9abf;
             14'h1a73 	:	val_out <= 16'h9ac4;
             14'h1a74 	:	val_out <= 16'h9ac9;
             14'h1a75 	:	val_out <= 16'h9ace;
             14'h1a76 	:	val_out <= 16'h9ad3;
             14'h1a77 	:	val_out <= 16'h9ad8;
             14'h1a78 	:	val_out <= 16'h9add;
             14'h1a79 	:	val_out <= 16'h9ae2;
             14'h1a7a 	:	val_out <= 16'h9ae7;
             14'h1a7b 	:	val_out <= 16'h9aec;
             14'h1a7c 	:	val_out <= 16'h9af1;
             14'h1a7d 	:	val_out <= 16'h9af6;
             14'h1a7e 	:	val_out <= 16'h9afb;
             14'h1a7f 	:	val_out <= 16'h9b00;
             14'h1a80 	:	val_out <= 16'h9b05;
             14'h1a81 	:	val_out <= 16'h9b0a;
             14'h1a82 	:	val_out <= 16'h9b0f;
             14'h1a83 	:	val_out <= 16'h9b14;
             14'h1a84 	:	val_out <= 16'h9b19;
             14'h1a85 	:	val_out <= 16'h9b1e;
             14'h1a86 	:	val_out <= 16'h9b23;
             14'h1a87 	:	val_out <= 16'h9b28;
             14'h1a88 	:	val_out <= 16'h9b2d;
             14'h1a89 	:	val_out <= 16'h9b32;
             14'h1a8a 	:	val_out <= 16'h9b37;
             14'h1a8b 	:	val_out <= 16'h9b3c;
             14'h1a8c 	:	val_out <= 16'h9b41;
             14'h1a8d 	:	val_out <= 16'h9b46;
             14'h1a8e 	:	val_out <= 16'h9b4b;
             14'h1a8f 	:	val_out <= 16'h9b50;
             14'h1a90 	:	val_out <= 16'h9b55;
             14'h1a91 	:	val_out <= 16'h9b5a;
             14'h1a92 	:	val_out <= 16'h9b5f;
             14'h1a93 	:	val_out <= 16'h9b64;
             14'h1a94 	:	val_out <= 16'h9b69;
             14'h1a95 	:	val_out <= 16'h9b6e;
             14'h1a96 	:	val_out <= 16'h9b73;
             14'h1a97 	:	val_out <= 16'h9b78;
             14'h1a98 	:	val_out <= 16'h9b7d;
             14'h1a99 	:	val_out <= 16'h9b82;
             14'h1a9a 	:	val_out <= 16'h9b87;
             14'h1a9b 	:	val_out <= 16'h9b8c;
             14'h1a9c 	:	val_out <= 16'h9b91;
             14'h1a9d 	:	val_out <= 16'h9b96;
             14'h1a9e 	:	val_out <= 16'h9b9b;
             14'h1a9f 	:	val_out <= 16'h9ba0;
             14'h1aa0 	:	val_out <= 16'h9ba5;
             14'h1aa1 	:	val_out <= 16'h9baa;
             14'h1aa2 	:	val_out <= 16'h9baf;
             14'h1aa3 	:	val_out <= 16'h9bb4;
             14'h1aa4 	:	val_out <= 16'h9bb9;
             14'h1aa5 	:	val_out <= 16'h9bbe;
             14'h1aa6 	:	val_out <= 16'h9bc3;
             14'h1aa7 	:	val_out <= 16'h9bc8;
             14'h1aa8 	:	val_out <= 16'h9bcc;
             14'h1aa9 	:	val_out <= 16'h9bd1;
             14'h1aaa 	:	val_out <= 16'h9bd6;
             14'h1aab 	:	val_out <= 16'h9bdb;
             14'h1aac 	:	val_out <= 16'h9be0;
             14'h1aad 	:	val_out <= 16'h9be5;
             14'h1aae 	:	val_out <= 16'h9bea;
             14'h1aaf 	:	val_out <= 16'h9bef;
             14'h1ab0 	:	val_out <= 16'h9bf4;
             14'h1ab1 	:	val_out <= 16'h9bf9;
             14'h1ab2 	:	val_out <= 16'h9bfe;
             14'h1ab3 	:	val_out <= 16'h9c03;
             14'h1ab4 	:	val_out <= 16'h9c08;
             14'h1ab5 	:	val_out <= 16'h9c0d;
             14'h1ab6 	:	val_out <= 16'h9c12;
             14'h1ab7 	:	val_out <= 16'h9c17;
             14'h1ab8 	:	val_out <= 16'h9c1c;
             14'h1ab9 	:	val_out <= 16'h9c21;
             14'h1aba 	:	val_out <= 16'h9c26;
             14'h1abb 	:	val_out <= 16'h9c2b;
             14'h1abc 	:	val_out <= 16'h9c30;
             14'h1abd 	:	val_out <= 16'h9c35;
             14'h1abe 	:	val_out <= 16'h9c3a;
             14'h1abf 	:	val_out <= 16'h9c3f;
             14'h1ac0 	:	val_out <= 16'h9c44;
             14'h1ac1 	:	val_out <= 16'h9c49;
             14'h1ac2 	:	val_out <= 16'h9c4e;
             14'h1ac3 	:	val_out <= 16'h9c53;
             14'h1ac4 	:	val_out <= 16'h9c58;
             14'h1ac5 	:	val_out <= 16'h9c5d;
             14'h1ac6 	:	val_out <= 16'h9c62;
             14'h1ac7 	:	val_out <= 16'h9c67;
             14'h1ac8 	:	val_out <= 16'h9c6c;
             14'h1ac9 	:	val_out <= 16'h9c71;
             14'h1aca 	:	val_out <= 16'h9c76;
             14'h1acb 	:	val_out <= 16'h9c7b;
             14'h1acc 	:	val_out <= 16'h9c80;
             14'h1acd 	:	val_out <= 16'h9c85;
             14'h1ace 	:	val_out <= 16'h9c8a;
             14'h1acf 	:	val_out <= 16'h9c8f;
             14'h1ad0 	:	val_out <= 16'h9c94;
             14'h1ad1 	:	val_out <= 16'h9c99;
             14'h1ad2 	:	val_out <= 16'h9c9e;
             14'h1ad3 	:	val_out <= 16'h9ca3;
             14'h1ad4 	:	val_out <= 16'h9ca7;
             14'h1ad5 	:	val_out <= 16'h9cac;
             14'h1ad6 	:	val_out <= 16'h9cb1;
             14'h1ad7 	:	val_out <= 16'h9cb6;
             14'h1ad8 	:	val_out <= 16'h9cbb;
             14'h1ad9 	:	val_out <= 16'h9cc0;
             14'h1ada 	:	val_out <= 16'h9cc5;
             14'h1adb 	:	val_out <= 16'h9cca;
             14'h1adc 	:	val_out <= 16'h9ccf;
             14'h1add 	:	val_out <= 16'h9cd4;
             14'h1ade 	:	val_out <= 16'h9cd9;
             14'h1adf 	:	val_out <= 16'h9cde;
             14'h1ae0 	:	val_out <= 16'h9ce3;
             14'h1ae1 	:	val_out <= 16'h9ce8;
             14'h1ae2 	:	val_out <= 16'h9ced;
             14'h1ae3 	:	val_out <= 16'h9cf2;
             14'h1ae4 	:	val_out <= 16'h9cf7;
             14'h1ae5 	:	val_out <= 16'h9cfc;
             14'h1ae6 	:	val_out <= 16'h9d01;
             14'h1ae7 	:	val_out <= 16'h9d06;
             14'h1ae8 	:	val_out <= 16'h9d0b;
             14'h1ae9 	:	val_out <= 16'h9d10;
             14'h1aea 	:	val_out <= 16'h9d15;
             14'h1aeb 	:	val_out <= 16'h9d1a;
             14'h1aec 	:	val_out <= 16'h9d1f;
             14'h1aed 	:	val_out <= 16'h9d24;
             14'h1aee 	:	val_out <= 16'h9d29;
             14'h1aef 	:	val_out <= 16'h9d2e;
             14'h1af0 	:	val_out <= 16'h9d32;
             14'h1af1 	:	val_out <= 16'h9d37;
             14'h1af2 	:	val_out <= 16'h9d3c;
             14'h1af3 	:	val_out <= 16'h9d41;
             14'h1af4 	:	val_out <= 16'h9d46;
             14'h1af5 	:	val_out <= 16'h9d4b;
             14'h1af6 	:	val_out <= 16'h9d50;
             14'h1af7 	:	val_out <= 16'h9d55;
             14'h1af8 	:	val_out <= 16'h9d5a;
             14'h1af9 	:	val_out <= 16'h9d5f;
             14'h1afa 	:	val_out <= 16'h9d64;
             14'h1afb 	:	val_out <= 16'h9d69;
             14'h1afc 	:	val_out <= 16'h9d6e;
             14'h1afd 	:	val_out <= 16'h9d73;
             14'h1afe 	:	val_out <= 16'h9d78;
             14'h1aff 	:	val_out <= 16'h9d7d;
             14'h1b00 	:	val_out <= 16'h9d82;
             14'h1b01 	:	val_out <= 16'h9d87;
             14'h1b02 	:	val_out <= 16'h9d8c;
             14'h1b03 	:	val_out <= 16'h9d91;
             14'h1b04 	:	val_out <= 16'h9d96;
             14'h1b05 	:	val_out <= 16'h9d9b;
             14'h1b06 	:	val_out <= 16'h9da0;
             14'h1b07 	:	val_out <= 16'h9da4;
             14'h1b08 	:	val_out <= 16'h9da9;
             14'h1b09 	:	val_out <= 16'h9dae;
             14'h1b0a 	:	val_out <= 16'h9db3;
             14'h1b0b 	:	val_out <= 16'h9db8;
             14'h1b0c 	:	val_out <= 16'h9dbd;
             14'h1b0d 	:	val_out <= 16'h9dc2;
             14'h1b0e 	:	val_out <= 16'h9dc7;
             14'h1b0f 	:	val_out <= 16'h9dcc;
             14'h1b10 	:	val_out <= 16'h9dd1;
             14'h1b11 	:	val_out <= 16'h9dd6;
             14'h1b12 	:	val_out <= 16'h9ddb;
             14'h1b13 	:	val_out <= 16'h9de0;
             14'h1b14 	:	val_out <= 16'h9de5;
             14'h1b15 	:	val_out <= 16'h9dea;
             14'h1b16 	:	val_out <= 16'h9def;
             14'h1b17 	:	val_out <= 16'h9df4;
             14'h1b18 	:	val_out <= 16'h9df9;
             14'h1b19 	:	val_out <= 16'h9dfe;
             14'h1b1a 	:	val_out <= 16'h9e02;
             14'h1b1b 	:	val_out <= 16'h9e07;
             14'h1b1c 	:	val_out <= 16'h9e0c;
             14'h1b1d 	:	val_out <= 16'h9e11;
             14'h1b1e 	:	val_out <= 16'h9e16;
             14'h1b1f 	:	val_out <= 16'h9e1b;
             14'h1b20 	:	val_out <= 16'h9e20;
             14'h1b21 	:	val_out <= 16'h9e25;
             14'h1b22 	:	val_out <= 16'h9e2a;
             14'h1b23 	:	val_out <= 16'h9e2f;
             14'h1b24 	:	val_out <= 16'h9e34;
             14'h1b25 	:	val_out <= 16'h9e39;
             14'h1b26 	:	val_out <= 16'h9e3e;
             14'h1b27 	:	val_out <= 16'h9e43;
             14'h1b28 	:	val_out <= 16'h9e48;
             14'h1b29 	:	val_out <= 16'h9e4d;
             14'h1b2a 	:	val_out <= 16'h9e51;
             14'h1b2b 	:	val_out <= 16'h9e56;
             14'h1b2c 	:	val_out <= 16'h9e5b;
             14'h1b2d 	:	val_out <= 16'h9e60;
             14'h1b2e 	:	val_out <= 16'h9e65;
             14'h1b2f 	:	val_out <= 16'h9e6a;
             14'h1b30 	:	val_out <= 16'h9e6f;
             14'h1b31 	:	val_out <= 16'h9e74;
             14'h1b32 	:	val_out <= 16'h9e79;
             14'h1b33 	:	val_out <= 16'h9e7e;
             14'h1b34 	:	val_out <= 16'h9e83;
             14'h1b35 	:	val_out <= 16'h9e88;
             14'h1b36 	:	val_out <= 16'h9e8d;
             14'h1b37 	:	val_out <= 16'h9e92;
             14'h1b38 	:	val_out <= 16'h9e97;
             14'h1b39 	:	val_out <= 16'h9e9c;
             14'h1b3a 	:	val_out <= 16'h9ea0;
             14'h1b3b 	:	val_out <= 16'h9ea5;
             14'h1b3c 	:	val_out <= 16'h9eaa;
             14'h1b3d 	:	val_out <= 16'h9eaf;
             14'h1b3e 	:	val_out <= 16'h9eb4;
             14'h1b3f 	:	val_out <= 16'h9eb9;
             14'h1b40 	:	val_out <= 16'h9ebe;
             14'h1b41 	:	val_out <= 16'h9ec3;
             14'h1b42 	:	val_out <= 16'h9ec8;
             14'h1b43 	:	val_out <= 16'h9ecd;
             14'h1b44 	:	val_out <= 16'h9ed2;
             14'h1b45 	:	val_out <= 16'h9ed7;
             14'h1b46 	:	val_out <= 16'h9edc;
             14'h1b47 	:	val_out <= 16'h9ee1;
             14'h1b48 	:	val_out <= 16'h9ee5;
             14'h1b49 	:	val_out <= 16'h9eea;
             14'h1b4a 	:	val_out <= 16'h9eef;
             14'h1b4b 	:	val_out <= 16'h9ef4;
             14'h1b4c 	:	val_out <= 16'h9ef9;
             14'h1b4d 	:	val_out <= 16'h9efe;
             14'h1b4e 	:	val_out <= 16'h9f03;
             14'h1b4f 	:	val_out <= 16'h9f08;
             14'h1b50 	:	val_out <= 16'h9f0d;
             14'h1b51 	:	val_out <= 16'h9f12;
             14'h1b52 	:	val_out <= 16'h9f17;
             14'h1b53 	:	val_out <= 16'h9f1c;
             14'h1b54 	:	val_out <= 16'h9f21;
             14'h1b55 	:	val_out <= 16'h9f25;
             14'h1b56 	:	val_out <= 16'h9f2a;
             14'h1b57 	:	val_out <= 16'h9f2f;
             14'h1b58 	:	val_out <= 16'h9f34;
             14'h1b59 	:	val_out <= 16'h9f39;
             14'h1b5a 	:	val_out <= 16'h9f3e;
             14'h1b5b 	:	val_out <= 16'h9f43;
             14'h1b5c 	:	val_out <= 16'h9f48;
             14'h1b5d 	:	val_out <= 16'h9f4d;
             14'h1b5e 	:	val_out <= 16'h9f52;
             14'h1b5f 	:	val_out <= 16'h9f57;
             14'h1b60 	:	val_out <= 16'h9f5c;
             14'h1b61 	:	val_out <= 16'h9f60;
             14'h1b62 	:	val_out <= 16'h9f65;
             14'h1b63 	:	val_out <= 16'h9f6a;
             14'h1b64 	:	val_out <= 16'h9f6f;
             14'h1b65 	:	val_out <= 16'h9f74;
             14'h1b66 	:	val_out <= 16'h9f79;
             14'h1b67 	:	val_out <= 16'h9f7e;
             14'h1b68 	:	val_out <= 16'h9f83;
             14'h1b69 	:	val_out <= 16'h9f88;
             14'h1b6a 	:	val_out <= 16'h9f8d;
             14'h1b6b 	:	val_out <= 16'h9f92;
             14'h1b6c 	:	val_out <= 16'h9f97;
             14'h1b6d 	:	val_out <= 16'h9f9b;
             14'h1b6e 	:	val_out <= 16'h9fa0;
             14'h1b6f 	:	val_out <= 16'h9fa5;
             14'h1b70 	:	val_out <= 16'h9faa;
             14'h1b71 	:	val_out <= 16'h9faf;
             14'h1b72 	:	val_out <= 16'h9fb4;
             14'h1b73 	:	val_out <= 16'h9fb9;
             14'h1b74 	:	val_out <= 16'h9fbe;
             14'h1b75 	:	val_out <= 16'h9fc3;
             14'h1b76 	:	val_out <= 16'h9fc8;
             14'h1b77 	:	val_out <= 16'h9fcd;
             14'h1b78 	:	val_out <= 16'h9fd1;
             14'h1b79 	:	val_out <= 16'h9fd6;
             14'h1b7a 	:	val_out <= 16'h9fdb;
             14'h1b7b 	:	val_out <= 16'h9fe0;
             14'h1b7c 	:	val_out <= 16'h9fe5;
             14'h1b7d 	:	val_out <= 16'h9fea;
             14'h1b7e 	:	val_out <= 16'h9fef;
             14'h1b7f 	:	val_out <= 16'h9ff4;
             14'h1b80 	:	val_out <= 16'h9ff9;
             14'h1b81 	:	val_out <= 16'h9ffe;
             14'h1b82 	:	val_out <= 16'ha003;
             14'h1b83 	:	val_out <= 16'ha007;
             14'h1b84 	:	val_out <= 16'ha00c;
             14'h1b85 	:	val_out <= 16'ha011;
             14'h1b86 	:	val_out <= 16'ha016;
             14'h1b87 	:	val_out <= 16'ha01b;
             14'h1b88 	:	val_out <= 16'ha020;
             14'h1b89 	:	val_out <= 16'ha025;
             14'h1b8a 	:	val_out <= 16'ha02a;
             14'h1b8b 	:	val_out <= 16'ha02f;
             14'h1b8c 	:	val_out <= 16'ha034;
             14'h1b8d 	:	val_out <= 16'ha038;
             14'h1b8e 	:	val_out <= 16'ha03d;
             14'h1b8f 	:	val_out <= 16'ha042;
             14'h1b90 	:	val_out <= 16'ha047;
             14'h1b91 	:	val_out <= 16'ha04c;
             14'h1b92 	:	val_out <= 16'ha051;
             14'h1b93 	:	val_out <= 16'ha056;
             14'h1b94 	:	val_out <= 16'ha05b;
             14'h1b95 	:	val_out <= 16'ha060;
             14'h1b96 	:	val_out <= 16'ha065;
             14'h1b97 	:	val_out <= 16'ha069;
             14'h1b98 	:	val_out <= 16'ha06e;
             14'h1b99 	:	val_out <= 16'ha073;
             14'h1b9a 	:	val_out <= 16'ha078;
             14'h1b9b 	:	val_out <= 16'ha07d;
             14'h1b9c 	:	val_out <= 16'ha082;
             14'h1b9d 	:	val_out <= 16'ha087;
             14'h1b9e 	:	val_out <= 16'ha08c;
             14'h1b9f 	:	val_out <= 16'ha091;
             14'h1ba0 	:	val_out <= 16'ha096;
             14'h1ba1 	:	val_out <= 16'ha09a;
             14'h1ba2 	:	val_out <= 16'ha09f;
             14'h1ba3 	:	val_out <= 16'ha0a4;
             14'h1ba4 	:	val_out <= 16'ha0a9;
             14'h1ba5 	:	val_out <= 16'ha0ae;
             14'h1ba6 	:	val_out <= 16'ha0b3;
             14'h1ba7 	:	val_out <= 16'ha0b8;
             14'h1ba8 	:	val_out <= 16'ha0bd;
             14'h1ba9 	:	val_out <= 16'ha0c2;
             14'h1baa 	:	val_out <= 16'ha0c6;
             14'h1bab 	:	val_out <= 16'ha0cb;
             14'h1bac 	:	val_out <= 16'ha0d0;
             14'h1bad 	:	val_out <= 16'ha0d5;
             14'h1bae 	:	val_out <= 16'ha0da;
             14'h1baf 	:	val_out <= 16'ha0df;
             14'h1bb0 	:	val_out <= 16'ha0e4;
             14'h1bb1 	:	val_out <= 16'ha0e9;
             14'h1bb2 	:	val_out <= 16'ha0ee;
             14'h1bb3 	:	val_out <= 16'ha0f2;
             14'h1bb4 	:	val_out <= 16'ha0f7;
             14'h1bb5 	:	val_out <= 16'ha0fc;
             14'h1bb6 	:	val_out <= 16'ha101;
             14'h1bb7 	:	val_out <= 16'ha106;
             14'h1bb8 	:	val_out <= 16'ha10b;
             14'h1bb9 	:	val_out <= 16'ha110;
             14'h1bba 	:	val_out <= 16'ha115;
             14'h1bbb 	:	val_out <= 16'ha11a;
             14'h1bbc 	:	val_out <= 16'ha11e;
             14'h1bbd 	:	val_out <= 16'ha123;
             14'h1bbe 	:	val_out <= 16'ha128;
             14'h1bbf 	:	val_out <= 16'ha12d;
             14'h1bc0 	:	val_out <= 16'ha132;
             14'h1bc1 	:	val_out <= 16'ha137;
             14'h1bc2 	:	val_out <= 16'ha13c;
             14'h1bc3 	:	val_out <= 16'ha141;
             14'h1bc4 	:	val_out <= 16'ha145;
             14'h1bc5 	:	val_out <= 16'ha14a;
             14'h1bc6 	:	val_out <= 16'ha14f;
             14'h1bc7 	:	val_out <= 16'ha154;
             14'h1bc8 	:	val_out <= 16'ha159;
             14'h1bc9 	:	val_out <= 16'ha15e;
             14'h1bca 	:	val_out <= 16'ha163;
             14'h1bcb 	:	val_out <= 16'ha168;
             14'h1bcc 	:	val_out <= 16'ha16c;
             14'h1bcd 	:	val_out <= 16'ha171;
             14'h1bce 	:	val_out <= 16'ha176;
             14'h1bcf 	:	val_out <= 16'ha17b;
             14'h1bd0 	:	val_out <= 16'ha180;
             14'h1bd1 	:	val_out <= 16'ha185;
             14'h1bd2 	:	val_out <= 16'ha18a;
             14'h1bd3 	:	val_out <= 16'ha18f;
             14'h1bd4 	:	val_out <= 16'ha193;
             14'h1bd5 	:	val_out <= 16'ha198;
             14'h1bd6 	:	val_out <= 16'ha19d;
             14'h1bd7 	:	val_out <= 16'ha1a2;
             14'h1bd8 	:	val_out <= 16'ha1a7;
             14'h1bd9 	:	val_out <= 16'ha1ac;
             14'h1bda 	:	val_out <= 16'ha1b1;
             14'h1bdb 	:	val_out <= 16'ha1b6;
             14'h1bdc 	:	val_out <= 16'ha1ba;
             14'h1bdd 	:	val_out <= 16'ha1bf;
             14'h1bde 	:	val_out <= 16'ha1c4;
             14'h1bdf 	:	val_out <= 16'ha1c9;
             14'h1be0 	:	val_out <= 16'ha1ce;
             14'h1be1 	:	val_out <= 16'ha1d3;
             14'h1be2 	:	val_out <= 16'ha1d8;
             14'h1be3 	:	val_out <= 16'ha1dd;
             14'h1be4 	:	val_out <= 16'ha1e1;
             14'h1be5 	:	val_out <= 16'ha1e6;
             14'h1be6 	:	val_out <= 16'ha1eb;
             14'h1be7 	:	val_out <= 16'ha1f0;
             14'h1be8 	:	val_out <= 16'ha1f5;
             14'h1be9 	:	val_out <= 16'ha1fa;
             14'h1bea 	:	val_out <= 16'ha1ff;
             14'h1beb 	:	val_out <= 16'ha203;
             14'h1bec 	:	val_out <= 16'ha208;
             14'h1bed 	:	val_out <= 16'ha20d;
             14'h1bee 	:	val_out <= 16'ha212;
             14'h1bef 	:	val_out <= 16'ha217;
             14'h1bf0 	:	val_out <= 16'ha21c;
             14'h1bf1 	:	val_out <= 16'ha221;
             14'h1bf2 	:	val_out <= 16'ha225;
             14'h1bf3 	:	val_out <= 16'ha22a;
             14'h1bf4 	:	val_out <= 16'ha22f;
             14'h1bf5 	:	val_out <= 16'ha234;
             14'h1bf6 	:	val_out <= 16'ha239;
             14'h1bf7 	:	val_out <= 16'ha23e;
             14'h1bf8 	:	val_out <= 16'ha243;
             14'h1bf9 	:	val_out <= 16'ha248;
             14'h1bfa 	:	val_out <= 16'ha24c;
             14'h1bfb 	:	val_out <= 16'ha251;
             14'h1bfc 	:	val_out <= 16'ha256;
             14'h1bfd 	:	val_out <= 16'ha25b;
             14'h1bfe 	:	val_out <= 16'ha260;
             14'h1bff 	:	val_out <= 16'ha265;
             14'h1c00 	:	val_out <= 16'ha26a;
             14'h1c01 	:	val_out <= 16'ha26e;
             14'h1c02 	:	val_out <= 16'ha273;
             14'h1c03 	:	val_out <= 16'ha278;
             14'h1c04 	:	val_out <= 16'ha27d;
             14'h1c05 	:	val_out <= 16'ha282;
             14'h1c06 	:	val_out <= 16'ha287;
             14'h1c07 	:	val_out <= 16'ha28c;
             14'h1c08 	:	val_out <= 16'ha290;
             14'h1c09 	:	val_out <= 16'ha295;
             14'h1c0a 	:	val_out <= 16'ha29a;
             14'h1c0b 	:	val_out <= 16'ha29f;
             14'h1c0c 	:	val_out <= 16'ha2a4;
             14'h1c0d 	:	val_out <= 16'ha2a9;
             14'h1c0e 	:	val_out <= 16'ha2ad;
             14'h1c0f 	:	val_out <= 16'ha2b2;
             14'h1c10 	:	val_out <= 16'ha2b7;
             14'h1c11 	:	val_out <= 16'ha2bc;
             14'h1c12 	:	val_out <= 16'ha2c1;
             14'h1c13 	:	val_out <= 16'ha2c6;
             14'h1c14 	:	val_out <= 16'ha2cb;
             14'h1c15 	:	val_out <= 16'ha2cf;
             14'h1c16 	:	val_out <= 16'ha2d4;
             14'h1c17 	:	val_out <= 16'ha2d9;
             14'h1c18 	:	val_out <= 16'ha2de;
             14'h1c19 	:	val_out <= 16'ha2e3;
             14'h1c1a 	:	val_out <= 16'ha2e8;
             14'h1c1b 	:	val_out <= 16'ha2ed;
             14'h1c1c 	:	val_out <= 16'ha2f1;
             14'h1c1d 	:	val_out <= 16'ha2f6;
             14'h1c1e 	:	val_out <= 16'ha2fb;
             14'h1c1f 	:	val_out <= 16'ha300;
             14'h1c20 	:	val_out <= 16'ha305;
             14'h1c21 	:	val_out <= 16'ha30a;
             14'h1c22 	:	val_out <= 16'ha30e;
             14'h1c23 	:	val_out <= 16'ha313;
             14'h1c24 	:	val_out <= 16'ha318;
             14'h1c25 	:	val_out <= 16'ha31d;
             14'h1c26 	:	val_out <= 16'ha322;
             14'h1c27 	:	val_out <= 16'ha327;
             14'h1c28 	:	val_out <= 16'ha32b;
             14'h1c29 	:	val_out <= 16'ha330;
             14'h1c2a 	:	val_out <= 16'ha335;
             14'h1c2b 	:	val_out <= 16'ha33a;
             14'h1c2c 	:	val_out <= 16'ha33f;
             14'h1c2d 	:	val_out <= 16'ha344;
             14'h1c2e 	:	val_out <= 16'ha349;
             14'h1c2f 	:	val_out <= 16'ha34d;
             14'h1c30 	:	val_out <= 16'ha352;
             14'h1c31 	:	val_out <= 16'ha357;
             14'h1c32 	:	val_out <= 16'ha35c;
             14'h1c33 	:	val_out <= 16'ha361;
             14'h1c34 	:	val_out <= 16'ha366;
             14'h1c35 	:	val_out <= 16'ha36a;
             14'h1c36 	:	val_out <= 16'ha36f;
             14'h1c37 	:	val_out <= 16'ha374;
             14'h1c38 	:	val_out <= 16'ha379;
             14'h1c39 	:	val_out <= 16'ha37e;
             14'h1c3a 	:	val_out <= 16'ha383;
             14'h1c3b 	:	val_out <= 16'ha387;
             14'h1c3c 	:	val_out <= 16'ha38c;
             14'h1c3d 	:	val_out <= 16'ha391;
             14'h1c3e 	:	val_out <= 16'ha396;
             14'h1c3f 	:	val_out <= 16'ha39b;
             14'h1c40 	:	val_out <= 16'ha3a0;
             14'h1c41 	:	val_out <= 16'ha3a4;
             14'h1c42 	:	val_out <= 16'ha3a9;
             14'h1c43 	:	val_out <= 16'ha3ae;
             14'h1c44 	:	val_out <= 16'ha3b3;
             14'h1c45 	:	val_out <= 16'ha3b8;
             14'h1c46 	:	val_out <= 16'ha3bd;
             14'h1c47 	:	val_out <= 16'ha3c1;
             14'h1c48 	:	val_out <= 16'ha3c6;
             14'h1c49 	:	val_out <= 16'ha3cb;
             14'h1c4a 	:	val_out <= 16'ha3d0;
             14'h1c4b 	:	val_out <= 16'ha3d5;
             14'h1c4c 	:	val_out <= 16'ha3da;
             14'h1c4d 	:	val_out <= 16'ha3de;
             14'h1c4e 	:	val_out <= 16'ha3e3;
             14'h1c4f 	:	val_out <= 16'ha3e8;
             14'h1c50 	:	val_out <= 16'ha3ed;
             14'h1c51 	:	val_out <= 16'ha3f2;
             14'h1c52 	:	val_out <= 16'ha3f6;
             14'h1c53 	:	val_out <= 16'ha3fb;
             14'h1c54 	:	val_out <= 16'ha400;
             14'h1c55 	:	val_out <= 16'ha405;
             14'h1c56 	:	val_out <= 16'ha40a;
             14'h1c57 	:	val_out <= 16'ha40f;
             14'h1c58 	:	val_out <= 16'ha413;
             14'h1c59 	:	val_out <= 16'ha418;
             14'h1c5a 	:	val_out <= 16'ha41d;
             14'h1c5b 	:	val_out <= 16'ha422;
             14'h1c5c 	:	val_out <= 16'ha427;
             14'h1c5d 	:	val_out <= 16'ha42c;
             14'h1c5e 	:	val_out <= 16'ha430;
             14'h1c5f 	:	val_out <= 16'ha435;
             14'h1c60 	:	val_out <= 16'ha43a;
             14'h1c61 	:	val_out <= 16'ha43f;
             14'h1c62 	:	val_out <= 16'ha444;
             14'h1c63 	:	val_out <= 16'ha448;
             14'h1c64 	:	val_out <= 16'ha44d;
             14'h1c65 	:	val_out <= 16'ha452;
             14'h1c66 	:	val_out <= 16'ha457;
             14'h1c67 	:	val_out <= 16'ha45c;
             14'h1c68 	:	val_out <= 16'ha461;
             14'h1c69 	:	val_out <= 16'ha465;
             14'h1c6a 	:	val_out <= 16'ha46a;
             14'h1c6b 	:	val_out <= 16'ha46f;
             14'h1c6c 	:	val_out <= 16'ha474;
             14'h1c6d 	:	val_out <= 16'ha479;
             14'h1c6e 	:	val_out <= 16'ha47d;
             14'h1c6f 	:	val_out <= 16'ha482;
             14'h1c70 	:	val_out <= 16'ha487;
             14'h1c71 	:	val_out <= 16'ha48c;
             14'h1c72 	:	val_out <= 16'ha491;
             14'h1c73 	:	val_out <= 16'ha496;
             14'h1c74 	:	val_out <= 16'ha49a;
             14'h1c75 	:	val_out <= 16'ha49f;
             14'h1c76 	:	val_out <= 16'ha4a4;
             14'h1c77 	:	val_out <= 16'ha4a9;
             14'h1c78 	:	val_out <= 16'ha4ae;
             14'h1c79 	:	val_out <= 16'ha4b2;
             14'h1c7a 	:	val_out <= 16'ha4b7;
             14'h1c7b 	:	val_out <= 16'ha4bc;
             14'h1c7c 	:	val_out <= 16'ha4c1;
             14'h1c7d 	:	val_out <= 16'ha4c6;
             14'h1c7e 	:	val_out <= 16'ha4ca;
             14'h1c7f 	:	val_out <= 16'ha4cf;
             14'h1c80 	:	val_out <= 16'ha4d4;
             14'h1c81 	:	val_out <= 16'ha4d9;
             14'h1c82 	:	val_out <= 16'ha4de;
             14'h1c83 	:	val_out <= 16'ha4e2;
             14'h1c84 	:	val_out <= 16'ha4e7;
             14'h1c85 	:	val_out <= 16'ha4ec;
             14'h1c86 	:	val_out <= 16'ha4f1;
             14'h1c87 	:	val_out <= 16'ha4f6;
             14'h1c88 	:	val_out <= 16'ha4fa;
             14'h1c89 	:	val_out <= 16'ha4ff;
             14'h1c8a 	:	val_out <= 16'ha504;
             14'h1c8b 	:	val_out <= 16'ha509;
             14'h1c8c 	:	val_out <= 16'ha50e;
             14'h1c8d 	:	val_out <= 16'ha513;
             14'h1c8e 	:	val_out <= 16'ha517;
             14'h1c8f 	:	val_out <= 16'ha51c;
             14'h1c90 	:	val_out <= 16'ha521;
             14'h1c91 	:	val_out <= 16'ha526;
             14'h1c92 	:	val_out <= 16'ha52b;
             14'h1c93 	:	val_out <= 16'ha52f;
             14'h1c94 	:	val_out <= 16'ha534;
             14'h1c95 	:	val_out <= 16'ha539;
             14'h1c96 	:	val_out <= 16'ha53e;
             14'h1c97 	:	val_out <= 16'ha543;
             14'h1c98 	:	val_out <= 16'ha547;
             14'h1c99 	:	val_out <= 16'ha54c;
             14'h1c9a 	:	val_out <= 16'ha551;
             14'h1c9b 	:	val_out <= 16'ha556;
             14'h1c9c 	:	val_out <= 16'ha55b;
             14'h1c9d 	:	val_out <= 16'ha55f;
             14'h1c9e 	:	val_out <= 16'ha564;
             14'h1c9f 	:	val_out <= 16'ha569;
             14'h1ca0 	:	val_out <= 16'ha56e;
             14'h1ca1 	:	val_out <= 16'ha572;
             14'h1ca2 	:	val_out <= 16'ha577;
             14'h1ca3 	:	val_out <= 16'ha57c;
             14'h1ca4 	:	val_out <= 16'ha581;
             14'h1ca5 	:	val_out <= 16'ha586;
             14'h1ca6 	:	val_out <= 16'ha58a;
             14'h1ca7 	:	val_out <= 16'ha58f;
             14'h1ca8 	:	val_out <= 16'ha594;
             14'h1ca9 	:	val_out <= 16'ha599;
             14'h1caa 	:	val_out <= 16'ha59e;
             14'h1cab 	:	val_out <= 16'ha5a2;
             14'h1cac 	:	val_out <= 16'ha5a7;
             14'h1cad 	:	val_out <= 16'ha5ac;
             14'h1cae 	:	val_out <= 16'ha5b1;
             14'h1caf 	:	val_out <= 16'ha5b6;
             14'h1cb0 	:	val_out <= 16'ha5ba;
             14'h1cb1 	:	val_out <= 16'ha5bf;
             14'h1cb2 	:	val_out <= 16'ha5c4;
             14'h1cb3 	:	val_out <= 16'ha5c9;
             14'h1cb4 	:	val_out <= 16'ha5ce;
             14'h1cb5 	:	val_out <= 16'ha5d2;
             14'h1cb6 	:	val_out <= 16'ha5d7;
             14'h1cb7 	:	val_out <= 16'ha5dc;
             14'h1cb8 	:	val_out <= 16'ha5e1;
             14'h1cb9 	:	val_out <= 16'ha5e5;
             14'h1cba 	:	val_out <= 16'ha5ea;
             14'h1cbb 	:	val_out <= 16'ha5ef;
             14'h1cbc 	:	val_out <= 16'ha5f4;
             14'h1cbd 	:	val_out <= 16'ha5f9;
             14'h1cbe 	:	val_out <= 16'ha5fd;
             14'h1cbf 	:	val_out <= 16'ha602;
             14'h1cc0 	:	val_out <= 16'ha607;
             14'h1cc1 	:	val_out <= 16'ha60c;
             14'h1cc2 	:	val_out <= 16'ha610;
             14'h1cc3 	:	val_out <= 16'ha615;
             14'h1cc4 	:	val_out <= 16'ha61a;
             14'h1cc5 	:	val_out <= 16'ha61f;
             14'h1cc6 	:	val_out <= 16'ha624;
             14'h1cc7 	:	val_out <= 16'ha628;
             14'h1cc8 	:	val_out <= 16'ha62d;
             14'h1cc9 	:	val_out <= 16'ha632;
             14'h1cca 	:	val_out <= 16'ha637;
             14'h1ccb 	:	val_out <= 16'ha63c;
             14'h1ccc 	:	val_out <= 16'ha640;
             14'h1ccd 	:	val_out <= 16'ha645;
             14'h1cce 	:	val_out <= 16'ha64a;
             14'h1ccf 	:	val_out <= 16'ha64f;
             14'h1cd0 	:	val_out <= 16'ha653;
             14'h1cd1 	:	val_out <= 16'ha658;
             14'h1cd2 	:	val_out <= 16'ha65d;
             14'h1cd3 	:	val_out <= 16'ha662;
             14'h1cd4 	:	val_out <= 16'ha667;
             14'h1cd5 	:	val_out <= 16'ha66b;
             14'h1cd6 	:	val_out <= 16'ha670;
             14'h1cd7 	:	val_out <= 16'ha675;
             14'h1cd8 	:	val_out <= 16'ha67a;
             14'h1cd9 	:	val_out <= 16'ha67e;
             14'h1cda 	:	val_out <= 16'ha683;
             14'h1cdb 	:	val_out <= 16'ha688;
             14'h1cdc 	:	val_out <= 16'ha68d;
             14'h1cdd 	:	val_out <= 16'ha691;
             14'h1cde 	:	val_out <= 16'ha696;
             14'h1cdf 	:	val_out <= 16'ha69b;
             14'h1ce0 	:	val_out <= 16'ha6a0;
             14'h1ce1 	:	val_out <= 16'ha6a5;
             14'h1ce2 	:	val_out <= 16'ha6a9;
             14'h1ce3 	:	val_out <= 16'ha6ae;
             14'h1ce4 	:	val_out <= 16'ha6b3;
             14'h1ce5 	:	val_out <= 16'ha6b8;
             14'h1ce6 	:	val_out <= 16'ha6bc;
             14'h1ce7 	:	val_out <= 16'ha6c1;
             14'h1ce8 	:	val_out <= 16'ha6c6;
             14'h1ce9 	:	val_out <= 16'ha6cb;
             14'h1cea 	:	val_out <= 16'ha6cf;
             14'h1ceb 	:	val_out <= 16'ha6d4;
             14'h1cec 	:	val_out <= 16'ha6d9;
             14'h1ced 	:	val_out <= 16'ha6de;
             14'h1cee 	:	val_out <= 16'ha6e3;
             14'h1cef 	:	val_out <= 16'ha6e7;
             14'h1cf0 	:	val_out <= 16'ha6ec;
             14'h1cf1 	:	val_out <= 16'ha6f1;
             14'h1cf2 	:	val_out <= 16'ha6f6;
             14'h1cf3 	:	val_out <= 16'ha6fa;
             14'h1cf4 	:	val_out <= 16'ha6ff;
             14'h1cf5 	:	val_out <= 16'ha704;
             14'h1cf6 	:	val_out <= 16'ha709;
             14'h1cf7 	:	val_out <= 16'ha70d;
             14'h1cf8 	:	val_out <= 16'ha712;
             14'h1cf9 	:	val_out <= 16'ha717;
             14'h1cfa 	:	val_out <= 16'ha71c;
             14'h1cfb 	:	val_out <= 16'ha720;
             14'h1cfc 	:	val_out <= 16'ha725;
             14'h1cfd 	:	val_out <= 16'ha72a;
             14'h1cfe 	:	val_out <= 16'ha72f;
             14'h1cff 	:	val_out <= 16'ha733;
             14'h1d00 	:	val_out <= 16'ha738;
             14'h1d01 	:	val_out <= 16'ha73d;
             14'h1d02 	:	val_out <= 16'ha742;
             14'h1d03 	:	val_out <= 16'ha746;
             14'h1d04 	:	val_out <= 16'ha74b;
             14'h1d05 	:	val_out <= 16'ha750;
             14'h1d06 	:	val_out <= 16'ha755;
             14'h1d07 	:	val_out <= 16'ha75a;
             14'h1d08 	:	val_out <= 16'ha75e;
             14'h1d09 	:	val_out <= 16'ha763;
             14'h1d0a 	:	val_out <= 16'ha768;
             14'h1d0b 	:	val_out <= 16'ha76d;
             14'h1d0c 	:	val_out <= 16'ha771;
             14'h1d0d 	:	val_out <= 16'ha776;
             14'h1d0e 	:	val_out <= 16'ha77b;
             14'h1d0f 	:	val_out <= 16'ha780;
             14'h1d10 	:	val_out <= 16'ha784;
             14'h1d11 	:	val_out <= 16'ha789;
             14'h1d12 	:	val_out <= 16'ha78e;
             14'h1d13 	:	val_out <= 16'ha793;
             14'h1d14 	:	val_out <= 16'ha797;
             14'h1d15 	:	val_out <= 16'ha79c;
             14'h1d16 	:	val_out <= 16'ha7a1;
             14'h1d17 	:	val_out <= 16'ha7a6;
             14'h1d18 	:	val_out <= 16'ha7aa;
             14'h1d19 	:	val_out <= 16'ha7af;
             14'h1d1a 	:	val_out <= 16'ha7b4;
             14'h1d1b 	:	val_out <= 16'ha7b9;
             14'h1d1c 	:	val_out <= 16'ha7bd;
             14'h1d1d 	:	val_out <= 16'ha7c2;
             14'h1d1e 	:	val_out <= 16'ha7c7;
             14'h1d1f 	:	val_out <= 16'ha7cc;
             14'h1d20 	:	val_out <= 16'ha7d0;
             14'h1d21 	:	val_out <= 16'ha7d5;
             14'h1d22 	:	val_out <= 16'ha7da;
             14'h1d23 	:	val_out <= 16'ha7de;
             14'h1d24 	:	val_out <= 16'ha7e3;
             14'h1d25 	:	val_out <= 16'ha7e8;
             14'h1d26 	:	val_out <= 16'ha7ed;
             14'h1d27 	:	val_out <= 16'ha7f1;
             14'h1d28 	:	val_out <= 16'ha7f6;
             14'h1d29 	:	val_out <= 16'ha7fb;
             14'h1d2a 	:	val_out <= 16'ha800;
             14'h1d2b 	:	val_out <= 16'ha804;
             14'h1d2c 	:	val_out <= 16'ha809;
             14'h1d2d 	:	val_out <= 16'ha80e;
             14'h1d2e 	:	val_out <= 16'ha813;
             14'h1d2f 	:	val_out <= 16'ha817;
             14'h1d30 	:	val_out <= 16'ha81c;
             14'h1d31 	:	val_out <= 16'ha821;
             14'h1d32 	:	val_out <= 16'ha826;
             14'h1d33 	:	val_out <= 16'ha82a;
             14'h1d34 	:	val_out <= 16'ha82f;
             14'h1d35 	:	val_out <= 16'ha834;
             14'h1d36 	:	val_out <= 16'ha839;
             14'h1d37 	:	val_out <= 16'ha83d;
             14'h1d38 	:	val_out <= 16'ha842;
             14'h1d39 	:	val_out <= 16'ha847;
             14'h1d3a 	:	val_out <= 16'ha84b;
             14'h1d3b 	:	val_out <= 16'ha850;
             14'h1d3c 	:	val_out <= 16'ha855;
             14'h1d3d 	:	val_out <= 16'ha85a;
             14'h1d3e 	:	val_out <= 16'ha85e;
             14'h1d3f 	:	val_out <= 16'ha863;
             14'h1d40 	:	val_out <= 16'ha868;
             14'h1d41 	:	val_out <= 16'ha86d;
             14'h1d42 	:	val_out <= 16'ha871;
             14'h1d43 	:	val_out <= 16'ha876;
             14'h1d44 	:	val_out <= 16'ha87b;
             14'h1d45 	:	val_out <= 16'ha880;
             14'h1d46 	:	val_out <= 16'ha884;
             14'h1d47 	:	val_out <= 16'ha889;
             14'h1d48 	:	val_out <= 16'ha88e;
             14'h1d49 	:	val_out <= 16'ha892;
             14'h1d4a 	:	val_out <= 16'ha897;
             14'h1d4b 	:	val_out <= 16'ha89c;
             14'h1d4c 	:	val_out <= 16'ha8a1;
             14'h1d4d 	:	val_out <= 16'ha8a5;
             14'h1d4e 	:	val_out <= 16'ha8aa;
             14'h1d4f 	:	val_out <= 16'ha8af;
             14'h1d50 	:	val_out <= 16'ha8b4;
             14'h1d51 	:	val_out <= 16'ha8b8;
             14'h1d52 	:	val_out <= 16'ha8bd;
             14'h1d53 	:	val_out <= 16'ha8c2;
             14'h1d54 	:	val_out <= 16'ha8c6;
             14'h1d55 	:	val_out <= 16'ha8cb;
             14'h1d56 	:	val_out <= 16'ha8d0;
             14'h1d57 	:	val_out <= 16'ha8d5;
             14'h1d58 	:	val_out <= 16'ha8d9;
             14'h1d59 	:	val_out <= 16'ha8de;
             14'h1d5a 	:	val_out <= 16'ha8e3;
             14'h1d5b 	:	val_out <= 16'ha8e8;
             14'h1d5c 	:	val_out <= 16'ha8ec;
             14'h1d5d 	:	val_out <= 16'ha8f1;
             14'h1d5e 	:	val_out <= 16'ha8f6;
             14'h1d5f 	:	val_out <= 16'ha8fa;
             14'h1d60 	:	val_out <= 16'ha8ff;
             14'h1d61 	:	val_out <= 16'ha904;
             14'h1d62 	:	val_out <= 16'ha909;
             14'h1d63 	:	val_out <= 16'ha90d;
             14'h1d64 	:	val_out <= 16'ha912;
             14'h1d65 	:	val_out <= 16'ha917;
             14'h1d66 	:	val_out <= 16'ha91b;
             14'h1d67 	:	val_out <= 16'ha920;
             14'h1d68 	:	val_out <= 16'ha925;
             14'h1d69 	:	val_out <= 16'ha92a;
             14'h1d6a 	:	val_out <= 16'ha92e;
             14'h1d6b 	:	val_out <= 16'ha933;
             14'h1d6c 	:	val_out <= 16'ha938;
             14'h1d6d 	:	val_out <= 16'ha93c;
             14'h1d6e 	:	val_out <= 16'ha941;
             14'h1d6f 	:	val_out <= 16'ha946;
             14'h1d70 	:	val_out <= 16'ha94b;
             14'h1d71 	:	val_out <= 16'ha94f;
             14'h1d72 	:	val_out <= 16'ha954;
             14'h1d73 	:	val_out <= 16'ha959;
             14'h1d74 	:	val_out <= 16'ha95d;
             14'h1d75 	:	val_out <= 16'ha962;
             14'h1d76 	:	val_out <= 16'ha967;
             14'h1d77 	:	val_out <= 16'ha96c;
             14'h1d78 	:	val_out <= 16'ha970;
             14'h1d79 	:	val_out <= 16'ha975;
             14'h1d7a 	:	val_out <= 16'ha97a;
             14'h1d7b 	:	val_out <= 16'ha97e;
             14'h1d7c 	:	val_out <= 16'ha983;
             14'h1d7d 	:	val_out <= 16'ha988;
             14'h1d7e 	:	val_out <= 16'ha98d;
             14'h1d7f 	:	val_out <= 16'ha991;
             14'h1d80 	:	val_out <= 16'ha996;
             14'h1d81 	:	val_out <= 16'ha99b;
             14'h1d82 	:	val_out <= 16'ha99f;
             14'h1d83 	:	val_out <= 16'ha9a4;
             14'h1d84 	:	val_out <= 16'ha9a9;
             14'h1d85 	:	val_out <= 16'ha9ad;
             14'h1d86 	:	val_out <= 16'ha9b2;
             14'h1d87 	:	val_out <= 16'ha9b7;
             14'h1d88 	:	val_out <= 16'ha9bc;
             14'h1d89 	:	val_out <= 16'ha9c0;
             14'h1d8a 	:	val_out <= 16'ha9c5;
             14'h1d8b 	:	val_out <= 16'ha9ca;
             14'h1d8c 	:	val_out <= 16'ha9ce;
             14'h1d8d 	:	val_out <= 16'ha9d3;
             14'h1d8e 	:	val_out <= 16'ha9d8;
             14'h1d8f 	:	val_out <= 16'ha9dc;
             14'h1d90 	:	val_out <= 16'ha9e1;
             14'h1d91 	:	val_out <= 16'ha9e6;
             14'h1d92 	:	val_out <= 16'ha9eb;
             14'h1d93 	:	val_out <= 16'ha9ef;
             14'h1d94 	:	val_out <= 16'ha9f4;
             14'h1d95 	:	val_out <= 16'ha9f9;
             14'h1d96 	:	val_out <= 16'ha9fd;
             14'h1d97 	:	val_out <= 16'haa02;
             14'h1d98 	:	val_out <= 16'haa07;
             14'h1d99 	:	val_out <= 16'haa0b;
             14'h1d9a 	:	val_out <= 16'haa10;
             14'h1d9b 	:	val_out <= 16'haa15;
             14'h1d9c 	:	val_out <= 16'haa1a;
             14'h1d9d 	:	val_out <= 16'haa1e;
             14'h1d9e 	:	val_out <= 16'haa23;
             14'h1d9f 	:	val_out <= 16'haa28;
             14'h1da0 	:	val_out <= 16'haa2c;
             14'h1da1 	:	val_out <= 16'haa31;
             14'h1da2 	:	val_out <= 16'haa36;
             14'h1da3 	:	val_out <= 16'haa3a;
             14'h1da4 	:	val_out <= 16'haa3f;
             14'h1da5 	:	val_out <= 16'haa44;
             14'h1da6 	:	val_out <= 16'haa49;
             14'h1da7 	:	val_out <= 16'haa4d;
             14'h1da8 	:	val_out <= 16'haa52;
             14'h1da9 	:	val_out <= 16'haa57;
             14'h1daa 	:	val_out <= 16'haa5b;
             14'h1dab 	:	val_out <= 16'haa60;
             14'h1dac 	:	val_out <= 16'haa65;
             14'h1dad 	:	val_out <= 16'haa69;
             14'h1dae 	:	val_out <= 16'haa6e;
             14'h1daf 	:	val_out <= 16'haa73;
             14'h1db0 	:	val_out <= 16'haa77;
             14'h1db1 	:	val_out <= 16'haa7c;
             14'h1db2 	:	val_out <= 16'haa81;
             14'h1db3 	:	val_out <= 16'haa85;
             14'h1db4 	:	val_out <= 16'haa8a;
             14'h1db5 	:	val_out <= 16'haa8f;
             14'h1db6 	:	val_out <= 16'haa94;
             14'h1db7 	:	val_out <= 16'haa98;
             14'h1db8 	:	val_out <= 16'haa9d;
             14'h1db9 	:	val_out <= 16'haaa2;
             14'h1dba 	:	val_out <= 16'haaa6;
             14'h1dbb 	:	val_out <= 16'haaab;
             14'h1dbc 	:	val_out <= 16'haab0;
             14'h1dbd 	:	val_out <= 16'haab4;
             14'h1dbe 	:	val_out <= 16'haab9;
             14'h1dbf 	:	val_out <= 16'haabe;
             14'h1dc0 	:	val_out <= 16'haac2;
             14'h1dc1 	:	val_out <= 16'haac7;
             14'h1dc2 	:	val_out <= 16'haacc;
             14'h1dc3 	:	val_out <= 16'haad0;
             14'h1dc4 	:	val_out <= 16'haad5;
             14'h1dc5 	:	val_out <= 16'haada;
             14'h1dc6 	:	val_out <= 16'haade;
             14'h1dc7 	:	val_out <= 16'haae3;
             14'h1dc8 	:	val_out <= 16'haae8;
             14'h1dc9 	:	val_out <= 16'haaec;
             14'h1dca 	:	val_out <= 16'haaf1;
             14'h1dcb 	:	val_out <= 16'haaf6;
             14'h1dcc 	:	val_out <= 16'haafa;
             14'h1dcd 	:	val_out <= 16'haaff;
             14'h1dce 	:	val_out <= 16'hab04;
             14'h1dcf 	:	val_out <= 16'hab09;
             14'h1dd0 	:	val_out <= 16'hab0d;
             14'h1dd1 	:	val_out <= 16'hab12;
             14'h1dd2 	:	val_out <= 16'hab17;
             14'h1dd3 	:	val_out <= 16'hab1b;
             14'h1dd4 	:	val_out <= 16'hab20;
             14'h1dd5 	:	val_out <= 16'hab25;
             14'h1dd6 	:	val_out <= 16'hab29;
             14'h1dd7 	:	val_out <= 16'hab2e;
             14'h1dd8 	:	val_out <= 16'hab33;
             14'h1dd9 	:	val_out <= 16'hab37;
             14'h1dda 	:	val_out <= 16'hab3c;
             14'h1ddb 	:	val_out <= 16'hab41;
             14'h1ddc 	:	val_out <= 16'hab45;
             14'h1ddd 	:	val_out <= 16'hab4a;
             14'h1dde 	:	val_out <= 16'hab4f;
             14'h1ddf 	:	val_out <= 16'hab53;
             14'h1de0 	:	val_out <= 16'hab58;
             14'h1de1 	:	val_out <= 16'hab5d;
             14'h1de2 	:	val_out <= 16'hab61;
             14'h1de3 	:	val_out <= 16'hab66;
             14'h1de4 	:	val_out <= 16'hab6b;
             14'h1de5 	:	val_out <= 16'hab6f;
             14'h1de6 	:	val_out <= 16'hab74;
             14'h1de7 	:	val_out <= 16'hab79;
             14'h1de8 	:	val_out <= 16'hab7d;
             14'h1de9 	:	val_out <= 16'hab82;
             14'h1dea 	:	val_out <= 16'hab87;
             14'h1deb 	:	val_out <= 16'hab8b;
             14'h1dec 	:	val_out <= 16'hab90;
             14'h1ded 	:	val_out <= 16'hab95;
             14'h1dee 	:	val_out <= 16'hab99;
             14'h1def 	:	val_out <= 16'hab9e;
             14'h1df0 	:	val_out <= 16'haba3;
             14'h1df1 	:	val_out <= 16'haba7;
             14'h1df2 	:	val_out <= 16'habac;
             14'h1df3 	:	val_out <= 16'habb1;
             14'h1df4 	:	val_out <= 16'habb5;
             14'h1df5 	:	val_out <= 16'habba;
             14'h1df6 	:	val_out <= 16'habbf;
             14'h1df7 	:	val_out <= 16'habc3;
             14'h1df8 	:	val_out <= 16'habc8;
             14'h1df9 	:	val_out <= 16'habcd;
             14'h1dfa 	:	val_out <= 16'habd1;
             14'h1dfb 	:	val_out <= 16'habd6;
             14'h1dfc 	:	val_out <= 16'habda;
             14'h1dfd 	:	val_out <= 16'habdf;
             14'h1dfe 	:	val_out <= 16'habe4;
             14'h1dff 	:	val_out <= 16'habe8;
             14'h1e00 	:	val_out <= 16'habed;
             14'h1e01 	:	val_out <= 16'habf2;
             14'h1e02 	:	val_out <= 16'habf6;
             14'h1e03 	:	val_out <= 16'habfb;
             14'h1e04 	:	val_out <= 16'hac00;
             14'h1e05 	:	val_out <= 16'hac04;
             14'h1e06 	:	val_out <= 16'hac09;
             14'h1e07 	:	val_out <= 16'hac0e;
             14'h1e08 	:	val_out <= 16'hac12;
             14'h1e09 	:	val_out <= 16'hac17;
             14'h1e0a 	:	val_out <= 16'hac1c;
             14'h1e0b 	:	val_out <= 16'hac20;
             14'h1e0c 	:	val_out <= 16'hac25;
             14'h1e0d 	:	val_out <= 16'hac2a;
             14'h1e0e 	:	val_out <= 16'hac2e;
             14'h1e0f 	:	val_out <= 16'hac33;
             14'h1e10 	:	val_out <= 16'hac38;
             14'h1e11 	:	val_out <= 16'hac3c;
             14'h1e12 	:	val_out <= 16'hac41;
             14'h1e13 	:	val_out <= 16'hac45;
             14'h1e14 	:	val_out <= 16'hac4a;
             14'h1e15 	:	val_out <= 16'hac4f;
             14'h1e16 	:	val_out <= 16'hac53;
             14'h1e17 	:	val_out <= 16'hac58;
             14'h1e18 	:	val_out <= 16'hac5d;
             14'h1e19 	:	val_out <= 16'hac61;
             14'h1e1a 	:	val_out <= 16'hac66;
             14'h1e1b 	:	val_out <= 16'hac6b;
             14'h1e1c 	:	val_out <= 16'hac6f;
             14'h1e1d 	:	val_out <= 16'hac74;
             14'h1e1e 	:	val_out <= 16'hac79;
             14'h1e1f 	:	val_out <= 16'hac7d;
             14'h1e20 	:	val_out <= 16'hac82;
             14'h1e21 	:	val_out <= 16'hac87;
             14'h1e22 	:	val_out <= 16'hac8b;
             14'h1e23 	:	val_out <= 16'hac90;
             14'h1e24 	:	val_out <= 16'hac94;
             14'h1e25 	:	val_out <= 16'hac99;
             14'h1e26 	:	val_out <= 16'hac9e;
             14'h1e27 	:	val_out <= 16'haca2;
             14'h1e28 	:	val_out <= 16'haca7;
             14'h1e29 	:	val_out <= 16'hacac;
             14'h1e2a 	:	val_out <= 16'hacb0;
             14'h1e2b 	:	val_out <= 16'hacb5;
             14'h1e2c 	:	val_out <= 16'hacba;
             14'h1e2d 	:	val_out <= 16'hacbe;
             14'h1e2e 	:	val_out <= 16'hacc3;
             14'h1e2f 	:	val_out <= 16'hacc7;
             14'h1e30 	:	val_out <= 16'haccc;
             14'h1e31 	:	val_out <= 16'hacd1;
             14'h1e32 	:	val_out <= 16'hacd5;
             14'h1e33 	:	val_out <= 16'hacda;
             14'h1e34 	:	val_out <= 16'hacdf;
             14'h1e35 	:	val_out <= 16'hace3;
             14'h1e36 	:	val_out <= 16'hace8;
             14'h1e37 	:	val_out <= 16'haced;
             14'h1e38 	:	val_out <= 16'hacf1;
             14'h1e39 	:	val_out <= 16'hacf6;
             14'h1e3a 	:	val_out <= 16'hacfa;
             14'h1e3b 	:	val_out <= 16'hacff;
             14'h1e3c 	:	val_out <= 16'had04;
             14'h1e3d 	:	val_out <= 16'had08;
             14'h1e3e 	:	val_out <= 16'had0d;
             14'h1e3f 	:	val_out <= 16'had12;
             14'h1e40 	:	val_out <= 16'had16;
             14'h1e41 	:	val_out <= 16'had1b;
             14'h1e42 	:	val_out <= 16'had1f;
             14'h1e43 	:	val_out <= 16'had24;
             14'h1e44 	:	val_out <= 16'had29;
             14'h1e45 	:	val_out <= 16'had2d;
             14'h1e46 	:	val_out <= 16'had32;
             14'h1e47 	:	val_out <= 16'had37;
             14'h1e48 	:	val_out <= 16'had3b;
             14'h1e49 	:	val_out <= 16'had40;
             14'h1e4a 	:	val_out <= 16'had44;
             14'h1e4b 	:	val_out <= 16'had49;
             14'h1e4c 	:	val_out <= 16'had4e;
             14'h1e4d 	:	val_out <= 16'had52;
             14'h1e4e 	:	val_out <= 16'had57;
             14'h1e4f 	:	val_out <= 16'had5c;
             14'h1e50 	:	val_out <= 16'had60;
             14'h1e51 	:	val_out <= 16'had65;
             14'h1e52 	:	val_out <= 16'had69;
             14'h1e53 	:	val_out <= 16'had6e;
             14'h1e54 	:	val_out <= 16'had73;
             14'h1e55 	:	val_out <= 16'had77;
             14'h1e56 	:	val_out <= 16'had7c;
             14'h1e57 	:	val_out <= 16'had81;
             14'h1e58 	:	val_out <= 16'had85;
             14'h1e59 	:	val_out <= 16'had8a;
             14'h1e5a 	:	val_out <= 16'had8e;
             14'h1e5b 	:	val_out <= 16'had93;
             14'h1e5c 	:	val_out <= 16'had98;
             14'h1e5d 	:	val_out <= 16'had9c;
             14'h1e5e 	:	val_out <= 16'hada1;
             14'h1e5f 	:	val_out <= 16'hada6;
             14'h1e60 	:	val_out <= 16'hadaa;
             14'h1e61 	:	val_out <= 16'hadaf;
             14'h1e62 	:	val_out <= 16'hadb3;
             14'h1e63 	:	val_out <= 16'hadb8;
             14'h1e64 	:	val_out <= 16'hadbd;
             14'h1e65 	:	val_out <= 16'hadc1;
             14'h1e66 	:	val_out <= 16'hadc6;
             14'h1e67 	:	val_out <= 16'hadca;
             14'h1e68 	:	val_out <= 16'hadcf;
             14'h1e69 	:	val_out <= 16'hadd4;
             14'h1e6a 	:	val_out <= 16'hadd8;
             14'h1e6b 	:	val_out <= 16'haddd;
             14'h1e6c 	:	val_out <= 16'hade2;
             14'h1e6d 	:	val_out <= 16'hade6;
             14'h1e6e 	:	val_out <= 16'hadeb;
             14'h1e6f 	:	val_out <= 16'hadef;
             14'h1e70 	:	val_out <= 16'hadf4;
             14'h1e71 	:	val_out <= 16'hadf9;
             14'h1e72 	:	val_out <= 16'hadfd;
             14'h1e73 	:	val_out <= 16'hae02;
             14'h1e74 	:	val_out <= 16'hae06;
             14'h1e75 	:	val_out <= 16'hae0b;
             14'h1e76 	:	val_out <= 16'hae10;
             14'h1e77 	:	val_out <= 16'hae14;
             14'h1e78 	:	val_out <= 16'hae19;
             14'h1e79 	:	val_out <= 16'hae1d;
             14'h1e7a 	:	val_out <= 16'hae22;
             14'h1e7b 	:	val_out <= 16'hae27;
             14'h1e7c 	:	val_out <= 16'hae2b;
             14'h1e7d 	:	val_out <= 16'hae30;
             14'h1e7e 	:	val_out <= 16'hae34;
             14'h1e7f 	:	val_out <= 16'hae39;
             14'h1e80 	:	val_out <= 16'hae3e;
             14'h1e81 	:	val_out <= 16'hae42;
             14'h1e82 	:	val_out <= 16'hae47;
             14'h1e83 	:	val_out <= 16'hae4b;
             14'h1e84 	:	val_out <= 16'hae50;
             14'h1e85 	:	val_out <= 16'hae55;
             14'h1e86 	:	val_out <= 16'hae59;
             14'h1e87 	:	val_out <= 16'hae5e;
             14'h1e88 	:	val_out <= 16'hae62;
             14'h1e89 	:	val_out <= 16'hae67;
             14'h1e8a 	:	val_out <= 16'hae6c;
             14'h1e8b 	:	val_out <= 16'hae70;
             14'h1e8c 	:	val_out <= 16'hae75;
             14'h1e8d 	:	val_out <= 16'hae79;
             14'h1e8e 	:	val_out <= 16'hae7e;
             14'h1e8f 	:	val_out <= 16'hae83;
             14'h1e90 	:	val_out <= 16'hae87;
             14'h1e91 	:	val_out <= 16'hae8c;
             14'h1e92 	:	val_out <= 16'hae90;
             14'h1e93 	:	val_out <= 16'hae95;
             14'h1e94 	:	val_out <= 16'hae9a;
             14'h1e95 	:	val_out <= 16'hae9e;
             14'h1e96 	:	val_out <= 16'haea3;
             14'h1e97 	:	val_out <= 16'haea7;
             14'h1e98 	:	val_out <= 16'haeac;
             14'h1e99 	:	val_out <= 16'haeb1;
             14'h1e9a 	:	val_out <= 16'haeb5;
             14'h1e9b 	:	val_out <= 16'haeba;
             14'h1e9c 	:	val_out <= 16'haebe;
             14'h1e9d 	:	val_out <= 16'haec3;
             14'h1e9e 	:	val_out <= 16'haec8;
             14'h1e9f 	:	val_out <= 16'haecc;
             14'h1ea0 	:	val_out <= 16'haed1;
             14'h1ea1 	:	val_out <= 16'haed5;
             14'h1ea2 	:	val_out <= 16'haeda;
             14'h1ea3 	:	val_out <= 16'haedf;
             14'h1ea4 	:	val_out <= 16'haee3;
             14'h1ea5 	:	val_out <= 16'haee8;
             14'h1ea6 	:	val_out <= 16'haeec;
             14'h1ea7 	:	val_out <= 16'haef1;
             14'h1ea8 	:	val_out <= 16'haef5;
             14'h1ea9 	:	val_out <= 16'haefa;
             14'h1eaa 	:	val_out <= 16'haeff;
             14'h1eab 	:	val_out <= 16'haf03;
             14'h1eac 	:	val_out <= 16'haf08;
             14'h1ead 	:	val_out <= 16'haf0c;
             14'h1eae 	:	val_out <= 16'haf11;
             14'h1eaf 	:	val_out <= 16'haf16;
             14'h1eb0 	:	val_out <= 16'haf1a;
             14'h1eb1 	:	val_out <= 16'haf1f;
             14'h1eb2 	:	val_out <= 16'haf23;
             14'h1eb3 	:	val_out <= 16'haf28;
             14'h1eb4 	:	val_out <= 16'haf2c;
             14'h1eb5 	:	val_out <= 16'haf31;
             14'h1eb6 	:	val_out <= 16'haf36;
             14'h1eb7 	:	val_out <= 16'haf3a;
             14'h1eb8 	:	val_out <= 16'haf3f;
             14'h1eb9 	:	val_out <= 16'haf43;
             14'h1eba 	:	val_out <= 16'haf48;
             14'h1ebb 	:	val_out <= 16'haf4d;
             14'h1ebc 	:	val_out <= 16'haf51;
             14'h1ebd 	:	val_out <= 16'haf56;
             14'h1ebe 	:	val_out <= 16'haf5a;
             14'h1ebf 	:	val_out <= 16'haf5f;
             14'h1ec0 	:	val_out <= 16'haf63;
             14'h1ec1 	:	val_out <= 16'haf68;
             14'h1ec2 	:	val_out <= 16'haf6d;
             14'h1ec3 	:	val_out <= 16'haf71;
             14'h1ec4 	:	val_out <= 16'haf76;
             14'h1ec5 	:	val_out <= 16'haf7a;
             14'h1ec6 	:	val_out <= 16'haf7f;
             14'h1ec7 	:	val_out <= 16'haf83;
             14'h1ec8 	:	val_out <= 16'haf88;
             14'h1ec9 	:	val_out <= 16'haf8d;
             14'h1eca 	:	val_out <= 16'haf91;
             14'h1ecb 	:	val_out <= 16'haf96;
             14'h1ecc 	:	val_out <= 16'haf9a;
             14'h1ecd 	:	val_out <= 16'haf9f;
             14'h1ece 	:	val_out <= 16'hafa3;
             14'h1ecf 	:	val_out <= 16'hafa8;
             14'h1ed0 	:	val_out <= 16'hafad;
             14'h1ed1 	:	val_out <= 16'hafb1;
             14'h1ed2 	:	val_out <= 16'hafb6;
             14'h1ed3 	:	val_out <= 16'hafba;
             14'h1ed4 	:	val_out <= 16'hafbf;
             14'h1ed5 	:	val_out <= 16'hafc3;
             14'h1ed6 	:	val_out <= 16'hafc8;
             14'h1ed7 	:	val_out <= 16'hafcd;
             14'h1ed8 	:	val_out <= 16'hafd1;
             14'h1ed9 	:	val_out <= 16'hafd6;
             14'h1eda 	:	val_out <= 16'hafda;
             14'h1edb 	:	val_out <= 16'hafdf;
             14'h1edc 	:	val_out <= 16'hafe3;
             14'h1edd 	:	val_out <= 16'hafe8;
             14'h1ede 	:	val_out <= 16'hafed;
             14'h1edf 	:	val_out <= 16'haff1;
             14'h1ee0 	:	val_out <= 16'haff6;
             14'h1ee1 	:	val_out <= 16'haffa;
             14'h1ee2 	:	val_out <= 16'hafff;
             14'h1ee3 	:	val_out <= 16'hb003;
             14'h1ee4 	:	val_out <= 16'hb008;
             14'h1ee5 	:	val_out <= 16'hb00c;
             14'h1ee6 	:	val_out <= 16'hb011;
             14'h1ee7 	:	val_out <= 16'hb016;
             14'h1ee8 	:	val_out <= 16'hb01a;
             14'h1ee9 	:	val_out <= 16'hb01f;
             14'h1eea 	:	val_out <= 16'hb023;
             14'h1eeb 	:	val_out <= 16'hb028;
             14'h1eec 	:	val_out <= 16'hb02c;
             14'h1eed 	:	val_out <= 16'hb031;
             14'h1eee 	:	val_out <= 16'hb036;
             14'h1eef 	:	val_out <= 16'hb03a;
             14'h1ef0 	:	val_out <= 16'hb03f;
             14'h1ef1 	:	val_out <= 16'hb043;
             14'h1ef2 	:	val_out <= 16'hb048;
             14'h1ef3 	:	val_out <= 16'hb04c;
             14'h1ef4 	:	val_out <= 16'hb051;
             14'h1ef5 	:	val_out <= 16'hb055;
             14'h1ef6 	:	val_out <= 16'hb05a;
             14'h1ef7 	:	val_out <= 16'hb05f;
             14'h1ef8 	:	val_out <= 16'hb063;
             14'h1ef9 	:	val_out <= 16'hb068;
             14'h1efa 	:	val_out <= 16'hb06c;
             14'h1efb 	:	val_out <= 16'hb071;
             14'h1efc 	:	val_out <= 16'hb075;
             14'h1efd 	:	val_out <= 16'hb07a;
             14'h1efe 	:	val_out <= 16'hb07e;
             14'h1eff 	:	val_out <= 16'hb083;
             14'h1f00 	:	val_out <= 16'hb088;
             14'h1f01 	:	val_out <= 16'hb08c;
             14'h1f02 	:	val_out <= 16'hb091;
             14'h1f03 	:	val_out <= 16'hb095;
             14'h1f04 	:	val_out <= 16'hb09a;
             14'h1f05 	:	val_out <= 16'hb09e;
             14'h1f06 	:	val_out <= 16'hb0a3;
             14'h1f07 	:	val_out <= 16'hb0a7;
             14'h1f08 	:	val_out <= 16'hb0ac;
             14'h1f09 	:	val_out <= 16'hb0b0;
             14'h1f0a 	:	val_out <= 16'hb0b5;
             14'h1f0b 	:	val_out <= 16'hb0ba;
             14'h1f0c 	:	val_out <= 16'hb0be;
             14'h1f0d 	:	val_out <= 16'hb0c3;
             14'h1f0e 	:	val_out <= 16'hb0c7;
             14'h1f0f 	:	val_out <= 16'hb0cc;
             14'h1f10 	:	val_out <= 16'hb0d0;
             14'h1f11 	:	val_out <= 16'hb0d5;
             14'h1f12 	:	val_out <= 16'hb0d9;
             14'h1f13 	:	val_out <= 16'hb0de;
             14'h1f14 	:	val_out <= 16'hb0e2;
             14'h1f15 	:	val_out <= 16'hb0e7;
             14'h1f16 	:	val_out <= 16'hb0ec;
             14'h1f17 	:	val_out <= 16'hb0f0;
             14'h1f18 	:	val_out <= 16'hb0f5;
             14'h1f19 	:	val_out <= 16'hb0f9;
             14'h1f1a 	:	val_out <= 16'hb0fe;
             14'h1f1b 	:	val_out <= 16'hb102;
             14'h1f1c 	:	val_out <= 16'hb107;
             14'h1f1d 	:	val_out <= 16'hb10b;
             14'h1f1e 	:	val_out <= 16'hb110;
             14'h1f1f 	:	val_out <= 16'hb114;
             14'h1f20 	:	val_out <= 16'hb119;
             14'h1f21 	:	val_out <= 16'hb11d;
             14'h1f22 	:	val_out <= 16'hb122;
             14'h1f23 	:	val_out <= 16'hb127;
             14'h1f24 	:	val_out <= 16'hb12b;
             14'h1f25 	:	val_out <= 16'hb130;
             14'h1f26 	:	val_out <= 16'hb134;
             14'h1f27 	:	val_out <= 16'hb139;
             14'h1f28 	:	val_out <= 16'hb13d;
             14'h1f29 	:	val_out <= 16'hb142;
             14'h1f2a 	:	val_out <= 16'hb146;
             14'h1f2b 	:	val_out <= 16'hb14b;
             14'h1f2c 	:	val_out <= 16'hb14f;
             14'h1f2d 	:	val_out <= 16'hb154;
             14'h1f2e 	:	val_out <= 16'hb158;
             14'h1f2f 	:	val_out <= 16'hb15d;
             14'h1f30 	:	val_out <= 16'hb161;
             14'h1f31 	:	val_out <= 16'hb166;
             14'h1f32 	:	val_out <= 16'hb16b;
             14'h1f33 	:	val_out <= 16'hb16f;
             14'h1f34 	:	val_out <= 16'hb174;
             14'h1f35 	:	val_out <= 16'hb178;
             14'h1f36 	:	val_out <= 16'hb17d;
             14'h1f37 	:	val_out <= 16'hb181;
             14'h1f38 	:	val_out <= 16'hb186;
             14'h1f39 	:	val_out <= 16'hb18a;
             14'h1f3a 	:	val_out <= 16'hb18f;
             14'h1f3b 	:	val_out <= 16'hb193;
             14'h1f3c 	:	val_out <= 16'hb198;
             14'h1f3d 	:	val_out <= 16'hb19c;
             14'h1f3e 	:	val_out <= 16'hb1a1;
             14'h1f3f 	:	val_out <= 16'hb1a5;
             14'h1f40 	:	val_out <= 16'hb1aa;
             14'h1f41 	:	val_out <= 16'hb1ae;
             14'h1f42 	:	val_out <= 16'hb1b3;
             14'h1f43 	:	val_out <= 16'hb1b7;
             14'h1f44 	:	val_out <= 16'hb1bc;
             14'h1f45 	:	val_out <= 16'hb1c0;
             14'h1f46 	:	val_out <= 16'hb1c5;
             14'h1f47 	:	val_out <= 16'hb1ca;
             14'h1f48 	:	val_out <= 16'hb1ce;
             14'h1f49 	:	val_out <= 16'hb1d3;
             14'h1f4a 	:	val_out <= 16'hb1d7;
             14'h1f4b 	:	val_out <= 16'hb1dc;
             14'h1f4c 	:	val_out <= 16'hb1e0;
             14'h1f4d 	:	val_out <= 16'hb1e5;
             14'h1f4e 	:	val_out <= 16'hb1e9;
             14'h1f4f 	:	val_out <= 16'hb1ee;
             14'h1f50 	:	val_out <= 16'hb1f2;
             14'h1f51 	:	val_out <= 16'hb1f7;
             14'h1f52 	:	val_out <= 16'hb1fb;
             14'h1f53 	:	val_out <= 16'hb200;
             14'h1f54 	:	val_out <= 16'hb204;
             14'h1f55 	:	val_out <= 16'hb209;
             14'h1f56 	:	val_out <= 16'hb20d;
             14'h1f57 	:	val_out <= 16'hb212;
             14'h1f58 	:	val_out <= 16'hb216;
             14'h1f59 	:	val_out <= 16'hb21b;
             14'h1f5a 	:	val_out <= 16'hb21f;
             14'h1f5b 	:	val_out <= 16'hb224;
             14'h1f5c 	:	val_out <= 16'hb228;
             14'h1f5d 	:	val_out <= 16'hb22d;
             14'h1f5e 	:	val_out <= 16'hb231;
             14'h1f5f 	:	val_out <= 16'hb236;
             14'h1f60 	:	val_out <= 16'hb23a;
             14'h1f61 	:	val_out <= 16'hb23f;
             14'h1f62 	:	val_out <= 16'hb243;
             14'h1f63 	:	val_out <= 16'hb248;
             14'h1f64 	:	val_out <= 16'hb24c;
             14'h1f65 	:	val_out <= 16'hb251;
             14'h1f66 	:	val_out <= 16'hb255;
             14'h1f67 	:	val_out <= 16'hb25a;
             14'h1f68 	:	val_out <= 16'hb25e;
             14'h1f69 	:	val_out <= 16'hb263;
             14'h1f6a 	:	val_out <= 16'hb268;
             14'h1f6b 	:	val_out <= 16'hb26c;
             14'h1f6c 	:	val_out <= 16'hb271;
             14'h1f6d 	:	val_out <= 16'hb275;
             14'h1f6e 	:	val_out <= 16'hb27a;
             14'h1f6f 	:	val_out <= 16'hb27e;
             14'h1f70 	:	val_out <= 16'hb283;
             14'h1f71 	:	val_out <= 16'hb287;
             14'h1f72 	:	val_out <= 16'hb28c;
             14'h1f73 	:	val_out <= 16'hb290;
             14'h1f74 	:	val_out <= 16'hb295;
             14'h1f75 	:	val_out <= 16'hb299;
             14'h1f76 	:	val_out <= 16'hb29e;
             14'h1f77 	:	val_out <= 16'hb2a2;
             14'h1f78 	:	val_out <= 16'hb2a7;
             14'h1f79 	:	val_out <= 16'hb2ab;
             14'h1f7a 	:	val_out <= 16'hb2b0;
             14'h1f7b 	:	val_out <= 16'hb2b4;
             14'h1f7c 	:	val_out <= 16'hb2b9;
             14'h1f7d 	:	val_out <= 16'hb2bd;
             14'h1f7e 	:	val_out <= 16'hb2c2;
             14'h1f7f 	:	val_out <= 16'hb2c6;
             14'h1f80 	:	val_out <= 16'hb2cb;
             14'h1f81 	:	val_out <= 16'hb2cf;
             14'h1f82 	:	val_out <= 16'hb2d4;
             14'h1f83 	:	val_out <= 16'hb2d8;
             14'h1f84 	:	val_out <= 16'hb2dd;
             14'h1f85 	:	val_out <= 16'hb2e1;
             14'h1f86 	:	val_out <= 16'hb2e6;
             14'h1f87 	:	val_out <= 16'hb2ea;
             14'h1f88 	:	val_out <= 16'hb2ee;
             14'h1f89 	:	val_out <= 16'hb2f3;
             14'h1f8a 	:	val_out <= 16'hb2f7;
             14'h1f8b 	:	val_out <= 16'hb2fc;
             14'h1f8c 	:	val_out <= 16'hb300;
             14'h1f8d 	:	val_out <= 16'hb305;
             14'h1f8e 	:	val_out <= 16'hb309;
             14'h1f8f 	:	val_out <= 16'hb30e;
             14'h1f90 	:	val_out <= 16'hb312;
             14'h1f91 	:	val_out <= 16'hb317;
             14'h1f92 	:	val_out <= 16'hb31b;
             14'h1f93 	:	val_out <= 16'hb320;
             14'h1f94 	:	val_out <= 16'hb324;
             14'h1f95 	:	val_out <= 16'hb329;
             14'h1f96 	:	val_out <= 16'hb32d;
             14'h1f97 	:	val_out <= 16'hb332;
             14'h1f98 	:	val_out <= 16'hb336;
             14'h1f99 	:	val_out <= 16'hb33b;
             14'h1f9a 	:	val_out <= 16'hb33f;
             14'h1f9b 	:	val_out <= 16'hb344;
             14'h1f9c 	:	val_out <= 16'hb348;
             14'h1f9d 	:	val_out <= 16'hb34d;
             14'h1f9e 	:	val_out <= 16'hb351;
             14'h1f9f 	:	val_out <= 16'hb356;
             14'h1fa0 	:	val_out <= 16'hb35a;
             14'h1fa1 	:	val_out <= 16'hb35f;
             14'h1fa2 	:	val_out <= 16'hb363;
             14'h1fa3 	:	val_out <= 16'hb368;
             14'h1fa4 	:	val_out <= 16'hb36c;
             14'h1fa5 	:	val_out <= 16'hb371;
             14'h1fa6 	:	val_out <= 16'hb375;
             14'h1fa7 	:	val_out <= 16'hb37a;
             14'h1fa8 	:	val_out <= 16'hb37e;
             14'h1fa9 	:	val_out <= 16'hb383;
             14'h1faa 	:	val_out <= 16'hb387;
             14'h1fab 	:	val_out <= 16'hb38c;
             14'h1fac 	:	val_out <= 16'hb390;
             14'h1fad 	:	val_out <= 16'hb394;
             14'h1fae 	:	val_out <= 16'hb399;
             14'h1faf 	:	val_out <= 16'hb39d;
             14'h1fb0 	:	val_out <= 16'hb3a2;
             14'h1fb1 	:	val_out <= 16'hb3a6;
             14'h1fb2 	:	val_out <= 16'hb3ab;
             14'h1fb3 	:	val_out <= 16'hb3af;
             14'h1fb4 	:	val_out <= 16'hb3b4;
             14'h1fb5 	:	val_out <= 16'hb3b8;
             14'h1fb6 	:	val_out <= 16'hb3bd;
             14'h1fb7 	:	val_out <= 16'hb3c1;
             14'h1fb8 	:	val_out <= 16'hb3c6;
             14'h1fb9 	:	val_out <= 16'hb3ca;
             14'h1fba 	:	val_out <= 16'hb3cf;
             14'h1fbb 	:	val_out <= 16'hb3d3;
             14'h1fbc 	:	val_out <= 16'hb3d8;
             14'h1fbd 	:	val_out <= 16'hb3dc;
             14'h1fbe 	:	val_out <= 16'hb3e1;
             14'h1fbf 	:	val_out <= 16'hb3e5;
             14'h1fc0 	:	val_out <= 16'hb3e9;
             14'h1fc1 	:	val_out <= 16'hb3ee;
             14'h1fc2 	:	val_out <= 16'hb3f2;
             14'h1fc3 	:	val_out <= 16'hb3f7;
             14'h1fc4 	:	val_out <= 16'hb3fb;
             14'h1fc5 	:	val_out <= 16'hb400;
             14'h1fc6 	:	val_out <= 16'hb404;
             14'h1fc7 	:	val_out <= 16'hb409;
             14'h1fc8 	:	val_out <= 16'hb40d;
             14'h1fc9 	:	val_out <= 16'hb412;
             14'h1fca 	:	val_out <= 16'hb416;
             14'h1fcb 	:	val_out <= 16'hb41b;
             14'h1fcc 	:	val_out <= 16'hb41f;
             14'h1fcd 	:	val_out <= 16'hb424;
             14'h1fce 	:	val_out <= 16'hb428;
             14'h1fcf 	:	val_out <= 16'hb42c;
             14'h1fd0 	:	val_out <= 16'hb431;
             14'h1fd1 	:	val_out <= 16'hb435;
             14'h1fd2 	:	val_out <= 16'hb43a;
             14'h1fd3 	:	val_out <= 16'hb43e;
             14'h1fd4 	:	val_out <= 16'hb443;
             14'h1fd5 	:	val_out <= 16'hb447;
             14'h1fd6 	:	val_out <= 16'hb44c;
             14'h1fd7 	:	val_out <= 16'hb450;
             14'h1fd8 	:	val_out <= 16'hb455;
             14'h1fd9 	:	val_out <= 16'hb459;
             14'h1fda 	:	val_out <= 16'hb45e;
             14'h1fdb 	:	val_out <= 16'hb462;
             14'h1fdc 	:	val_out <= 16'hb466;
             14'h1fdd 	:	val_out <= 16'hb46b;
             14'h1fde 	:	val_out <= 16'hb46f;
             14'h1fdf 	:	val_out <= 16'hb474;
             14'h1fe0 	:	val_out <= 16'hb478;
             14'h1fe1 	:	val_out <= 16'hb47d;
             14'h1fe2 	:	val_out <= 16'hb481;
             14'h1fe3 	:	val_out <= 16'hb486;
             14'h1fe4 	:	val_out <= 16'hb48a;
             14'h1fe5 	:	val_out <= 16'hb48f;
             14'h1fe6 	:	val_out <= 16'hb493;
             14'h1fe7 	:	val_out <= 16'hb497;
             14'h1fe8 	:	val_out <= 16'hb49c;
             14'h1fe9 	:	val_out <= 16'hb4a0;
             14'h1fea 	:	val_out <= 16'hb4a5;
             14'h1feb 	:	val_out <= 16'hb4a9;
             14'h1fec 	:	val_out <= 16'hb4ae;
             14'h1fed 	:	val_out <= 16'hb4b2;
             14'h1fee 	:	val_out <= 16'hb4b7;
             14'h1fef 	:	val_out <= 16'hb4bb;
             14'h1ff0 	:	val_out <= 16'hb4c0;
             14'h1ff1 	:	val_out <= 16'hb4c4;
             14'h1ff2 	:	val_out <= 16'hb4c8;
             14'h1ff3 	:	val_out <= 16'hb4cd;
             14'h1ff4 	:	val_out <= 16'hb4d1;
             14'h1ff5 	:	val_out <= 16'hb4d6;
             14'h1ff6 	:	val_out <= 16'hb4da;
             14'h1ff7 	:	val_out <= 16'hb4df;
             14'h1ff8 	:	val_out <= 16'hb4e3;
             14'h1ff9 	:	val_out <= 16'hb4e8;
             14'h1ffa 	:	val_out <= 16'hb4ec;
             14'h1ffb 	:	val_out <= 16'hb4f0;
             14'h1ffc 	:	val_out <= 16'hb4f5;
             14'h1ffd 	:	val_out <= 16'hb4f9;
             14'h1ffe 	:	val_out <= 16'hb4fe;
             14'h1fff 	:	val_out <= 16'hb502;
             14'h2000 	:	val_out <= 16'hb507;
             14'h2001 	:	val_out <= 16'hb50b;
             14'h2002 	:	val_out <= 16'hb510;
             14'h2003 	:	val_out <= 16'hb514;
             14'h2004 	:	val_out <= 16'hb518;
             14'h2005 	:	val_out <= 16'hb51d;
             14'h2006 	:	val_out <= 16'hb521;
             14'h2007 	:	val_out <= 16'hb526;
             14'h2008 	:	val_out <= 16'hb52a;
             14'h2009 	:	val_out <= 16'hb52f;
             14'h200a 	:	val_out <= 16'hb533;
             14'h200b 	:	val_out <= 16'hb538;
             14'h200c 	:	val_out <= 16'hb53c;
             14'h200d 	:	val_out <= 16'hb540;
             14'h200e 	:	val_out <= 16'hb545;
             14'h200f 	:	val_out <= 16'hb549;
             14'h2010 	:	val_out <= 16'hb54e;
             14'h2011 	:	val_out <= 16'hb552;
             14'h2012 	:	val_out <= 16'hb557;
             14'h2013 	:	val_out <= 16'hb55b;
             14'h2014 	:	val_out <= 16'hb55f;
             14'h2015 	:	val_out <= 16'hb564;
             14'h2016 	:	val_out <= 16'hb568;
             14'h2017 	:	val_out <= 16'hb56d;
             14'h2018 	:	val_out <= 16'hb571;
             14'h2019 	:	val_out <= 16'hb576;
             14'h201a 	:	val_out <= 16'hb57a;
             14'h201b 	:	val_out <= 16'hb57e;
             14'h201c 	:	val_out <= 16'hb583;
             14'h201d 	:	val_out <= 16'hb587;
             14'h201e 	:	val_out <= 16'hb58c;
             14'h201f 	:	val_out <= 16'hb590;
             14'h2020 	:	val_out <= 16'hb595;
             14'h2021 	:	val_out <= 16'hb599;
             14'h2022 	:	val_out <= 16'hb59d;
             14'h2023 	:	val_out <= 16'hb5a2;
             14'h2024 	:	val_out <= 16'hb5a6;
             14'h2025 	:	val_out <= 16'hb5ab;
             14'h2026 	:	val_out <= 16'hb5af;
             14'h2027 	:	val_out <= 16'hb5b4;
             14'h2028 	:	val_out <= 16'hb5b8;
             14'h2029 	:	val_out <= 16'hb5bc;
             14'h202a 	:	val_out <= 16'hb5c1;
             14'h202b 	:	val_out <= 16'hb5c5;
             14'h202c 	:	val_out <= 16'hb5ca;
             14'h202d 	:	val_out <= 16'hb5ce;
             14'h202e 	:	val_out <= 16'hb5d3;
             14'h202f 	:	val_out <= 16'hb5d7;
             14'h2030 	:	val_out <= 16'hb5db;
             14'h2031 	:	val_out <= 16'hb5e0;
             14'h2032 	:	val_out <= 16'hb5e4;
             14'h2033 	:	val_out <= 16'hb5e9;
             14'h2034 	:	val_out <= 16'hb5ed;
             14'h2035 	:	val_out <= 16'hb5f2;
             14'h2036 	:	val_out <= 16'hb5f6;
             14'h2037 	:	val_out <= 16'hb5fa;
             14'h2038 	:	val_out <= 16'hb5ff;
             14'h2039 	:	val_out <= 16'hb603;
             14'h203a 	:	val_out <= 16'hb608;
             14'h203b 	:	val_out <= 16'hb60c;
             14'h203c 	:	val_out <= 16'hb610;
             14'h203d 	:	val_out <= 16'hb615;
             14'h203e 	:	val_out <= 16'hb619;
             14'h203f 	:	val_out <= 16'hb61e;
             14'h2040 	:	val_out <= 16'hb622;
             14'h2041 	:	val_out <= 16'hb627;
             14'h2042 	:	val_out <= 16'hb62b;
             14'h2043 	:	val_out <= 16'hb62f;
             14'h2044 	:	val_out <= 16'hb634;
             14'h2045 	:	val_out <= 16'hb638;
             14'h2046 	:	val_out <= 16'hb63d;
             14'h2047 	:	val_out <= 16'hb641;
             14'h2048 	:	val_out <= 16'hb645;
             14'h2049 	:	val_out <= 16'hb64a;
             14'h204a 	:	val_out <= 16'hb64e;
             14'h204b 	:	val_out <= 16'hb653;
             14'h204c 	:	val_out <= 16'hb657;
             14'h204d 	:	val_out <= 16'hb65b;
             14'h204e 	:	val_out <= 16'hb660;
             14'h204f 	:	val_out <= 16'hb664;
             14'h2050 	:	val_out <= 16'hb669;
             14'h2051 	:	val_out <= 16'hb66d;
             14'h2052 	:	val_out <= 16'hb672;
             14'h2053 	:	val_out <= 16'hb676;
             14'h2054 	:	val_out <= 16'hb67a;
             14'h2055 	:	val_out <= 16'hb67f;
             14'h2056 	:	val_out <= 16'hb683;
             14'h2057 	:	val_out <= 16'hb688;
             14'h2058 	:	val_out <= 16'hb68c;
             14'h2059 	:	val_out <= 16'hb690;
             14'h205a 	:	val_out <= 16'hb695;
             14'h205b 	:	val_out <= 16'hb699;
             14'h205c 	:	val_out <= 16'hb69e;
             14'h205d 	:	val_out <= 16'hb6a2;
             14'h205e 	:	val_out <= 16'hb6a6;
             14'h205f 	:	val_out <= 16'hb6ab;
             14'h2060 	:	val_out <= 16'hb6af;
             14'h2061 	:	val_out <= 16'hb6b4;
             14'h2062 	:	val_out <= 16'hb6b8;
             14'h2063 	:	val_out <= 16'hb6bc;
             14'h2064 	:	val_out <= 16'hb6c1;
             14'h2065 	:	val_out <= 16'hb6c5;
             14'h2066 	:	val_out <= 16'hb6ca;
             14'h2067 	:	val_out <= 16'hb6ce;
             14'h2068 	:	val_out <= 16'hb6d2;
             14'h2069 	:	val_out <= 16'hb6d7;
             14'h206a 	:	val_out <= 16'hb6db;
             14'h206b 	:	val_out <= 16'hb6e0;
             14'h206c 	:	val_out <= 16'hb6e4;
             14'h206d 	:	val_out <= 16'hb6e8;
             14'h206e 	:	val_out <= 16'hb6ed;
             14'h206f 	:	val_out <= 16'hb6f1;
             14'h2070 	:	val_out <= 16'hb6f6;
             14'h2071 	:	val_out <= 16'hb6fa;
             14'h2072 	:	val_out <= 16'hb6fe;
             14'h2073 	:	val_out <= 16'hb703;
             14'h2074 	:	val_out <= 16'hb707;
             14'h2075 	:	val_out <= 16'hb70c;
             14'h2076 	:	val_out <= 16'hb710;
             14'h2077 	:	val_out <= 16'hb714;
             14'h2078 	:	val_out <= 16'hb719;
             14'h2079 	:	val_out <= 16'hb71d;
             14'h207a 	:	val_out <= 16'hb721;
             14'h207b 	:	val_out <= 16'hb726;
             14'h207c 	:	val_out <= 16'hb72a;
             14'h207d 	:	val_out <= 16'hb72f;
             14'h207e 	:	val_out <= 16'hb733;
             14'h207f 	:	val_out <= 16'hb737;
             14'h2080 	:	val_out <= 16'hb73c;
             14'h2081 	:	val_out <= 16'hb740;
             14'h2082 	:	val_out <= 16'hb745;
             14'h2083 	:	val_out <= 16'hb749;
             14'h2084 	:	val_out <= 16'hb74d;
             14'h2085 	:	val_out <= 16'hb752;
             14'h2086 	:	val_out <= 16'hb756;
             14'h2087 	:	val_out <= 16'hb75b;
             14'h2088 	:	val_out <= 16'hb75f;
             14'h2089 	:	val_out <= 16'hb763;
             14'h208a 	:	val_out <= 16'hb768;
             14'h208b 	:	val_out <= 16'hb76c;
             14'h208c 	:	val_out <= 16'hb770;
             14'h208d 	:	val_out <= 16'hb775;
             14'h208e 	:	val_out <= 16'hb779;
             14'h208f 	:	val_out <= 16'hb77e;
             14'h2090 	:	val_out <= 16'hb782;
             14'h2091 	:	val_out <= 16'hb786;
             14'h2092 	:	val_out <= 16'hb78b;
             14'h2093 	:	val_out <= 16'hb78f;
             14'h2094 	:	val_out <= 16'hb793;
             14'h2095 	:	val_out <= 16'hb798;
             14'h2096 	:	val_out <= 16'hb79c;
             14'h2097 	:	val_out <= 16'hb7a1;
             14'h2098 	:	val_out <= 16'hb7a5;
             14'h2099 	:	val_out <= 16'hb7a9;
             14'h209a 	:	val_out <= 16'hb7ae;
             14'h209b 	:	val_out <= 16'hb7b2;
             14'h209c 	:	val_out <= 16'hb7b7;
             14'h209d 	:	val_out <= 16'hb7bb;
             14'h209e 	:	val_out <= 16'hb7bf;
             14'h209f 	:	val_out <= 16'hb7c4;
             14'h20a0 	:	val_out <= 16'hb7c8;
             14'h20a1 	:	val_out <= 16'hb7cc;
             14'h20a2 	:	val_out <= 16'hb7d1;
             14'h20a3 	:	val_out <= 16'hb7d5;
             14'h20a4 	:	val_out <= 16'hb7da;
             14'h20a5 	:	val_out <= 16'hb7de;
             14'h20a6 	:	val_out <= 16'hb7e2;
             14'h20a7 	:	val_out <= 16'hb7e7;
             14'h20a8 	:	val_out <= 16'hb7eb;
             14'h20a9 	:	val_out <= 16'hb7ef;
             14'h20aa 	:	val_out <= 16'hb7f4;
             14'h20ab 	:	val_out <= 16'hb7f8;
             14'h20ac 	:	val_out <= 16'hb7fc;
             14'h20ad 	:	val_out <= 16'hb801;
             14'h20ae 	:	val_out <= 16'hb805;
             14'h20af 	:	val_out <= 16'hb80a;
             14'h20b0 	:	val_out <= 16'hb80e;
             14'h20b1 	:	val_out <= 16'hb812;
             14'h20b2 	:	val_out <= 16'hb817;
             14'h20b3 	:	val_out <= 16'hb81b;
             14'h20b4 	:	val_out <= 16'hb81f;
             14'h20b5 	:	val_out <= 16'hb824;
             14'h20b6 	:	val_out <= 16'hb828;
             14'h20b7 	:	val_out <= 16'hb82d;
             14'h20b8 	:	val_out <= 16'hb831;
             14'h20b9 	:	val_out <= 16'hb835;
             14'h20ba 	:	val_out <= 16'hb83a;
             14'h20bb 	:	val_out <= 16'hb83e;
             14'h20bc 	:	val_out <= 16'hb842;
             14'h20bd 	:	val_out <= 16'hb847;
             14'h20be 	:	val_out <= 16'hb84b;
             14'h20bf 	:	val_out <= 16'hb84f;
             14'h20c0 	:	val_out <= 16'hb854;
             14'h20c1 	:	val_out <= 16'hb858;
             14'h20c2 	:	val_out <= 16'hb85c;
             14'h20c3 	:	val_out <= 16'hb861;
             14'h20c4 	:	val_out <= 16'hb865;
             14'h20c5 	:	val_out <= 16'hb86a;
             14'h20c6 	:	val_out <= 16'hb86e;
             14'h20c7 	:	val_out <= 16'hb872;
             14'h20c8 	:	val_out <= 16'hb877;
             14'h20c9 	:	val_out <= 16'hb87b;
             14'h20ca 	:	val_out <= 16'hb87f;
             14'h20cb 	:	val_out <= 16'hb884;
             14'h20cc 	:	val_out <= 16'hb888;
             14'h20cd 	:	val_out <= 16'hb88c;
             14'h20ce 	:	val_out <= 16'hb891;
             14'h20cf 	:	val_out <= 16'hb895;
             14'h20d0 	:	val_out <= 16'hb899;
             14'h20d1 	:	val_out <= 16'hb89e;
             14'h20d2 	:	val_out <= 16'hb8a2;
             14'h20d3 	:	val_out <= 16'hb8a7;
             14'h20d4 	:	val_out <= 16'hb8ab;
             14'h20d5 	:	val_out <= 16'hb8af;
             14'h20d6 	:	val_out <= 16'hb8b4;
             14'h20d7 	:	val_out <= 16'hb8b8;
             14'h20d8 	:	val_out <= 16'hb8bc;
             14'h20d9 	:	val_out <= 16'hb8c1;
             14'h20da 	:	val_out <= 16'hb8c5;
             14'h20db 	:	val_out <= 16'hb8c9;
             14'h20dc 	:	val_out <= 16'hb8ce;
             14'h20dd 	:	val_out <= 16'hb8d2;
             14'h20de 	:	val_out <= 16'hb8d6;
             14'h20df 	:	val_out <= 16'hb8db;
             14'h20e0 	:	val_out <= 16'hb8df;
             14'h20e1 	:	val_out <= 16'hb8e3;
             14'h20e2 	:	val_out <= 16'hb8e8;
             14'h20e3 	:	val_out <= 16'hb8ec;
             14'h20e4 	:	val_out <= 16'hb8f0;
             14'h20e5 	:	val_out <= 16'hb8f5;
             14'h20e6 	:	val_out <= 16'hb8f9;
             14'h20e7 	:	val_out <= 16'hb8fd;
             14'h20e8 	:	val_out <= 16'hb902;
             14'h20e9 	:	val_out <= 16'hb906;
             14'h20ea 	:	val_out <= 16'hb90b;
             14'h20eb 	:	val_out <= 16'hb90f;
             14'h20ec 	:	val_out <= 16'hb913;
             14'h20ed 	:	val_out <= 16'hb918;
             14'h20ee 	:	val_out <= 16'hb91c;
             14'h20ef 	:	val_out <= 16'hb920;
             14'h20f0 	:	val_out <= 16'hb925;
             14'h20f1 	:	val_out <= 16'hb929;
             14'h20f2 	:	val_out <= 16'hb92d;
             14'h20f3 	:	val_out <= 16'hb932;
             14'h20f4 	:	val_out <= 16'hb936;
             14'h20f5 	:	val_out <= 16'hb93a;
             14'h20f6 	:	val_out <= 16'hb93f;
             14'h20f7 	:	val_out <= 16'hb943;
             14'h20f8 	:	val_out <= 16'hb947;
             14'h20f9 	:	val_out <= 16'hb94c;
             14'h20fa 	:	val_out <= 16'hb950;
             14'h20fb 	:	val_out <= 16'hb954;
             14'h20fc 	:	val_out <= 16'hb959;
             14'h20fd 	:	val_out <= 16'hb95d;
             14'h20fe 	:	val_out <= 16'hb961;
             14'h20ff 	:	val_out <= 16'hb966;
             14'h2100 	:	val_out <= 16'hb96a;
             14'h2101 	:	val_out <= 16'hb96e;
             14'h2102 	:	val_out <= 16'hb973;
             14'h2103 	:	val_out <= 16'hb977;
             14'h2104 	:	val_out <= 16'hb97b;
             14'h2105 	:	val_out <= 16'hb980;
             14'h2106 	:	val_out <= 16'hb984;
             14'h2107 	:	val_out <= 16'hb988;
             14'h2108 	:	val_out <= 16'hb98d;
             14'h2109 	:	val_out <= 16'hb991;
             14'h210a 	:	val_out <= 16'hb995;
             14'h210b 	:	val_out <= 16'hb99a;
             14'h210c 	:	val_out <= 16'hb99e;
             14'h210d 	:	val_out <= 16'hb9a2;
             14'h210e 	:	val_out <= 16'hb9a7;
             14'h210f 	:	val_out <= 16'hb9ab;
             14'h2110 	:	val_out <= 16'hb9af;
             14'h2111 	:	val_out <= 16'hb9b4;
             14'h2112 	:	val_out <= 16'hb9b8;
             14'h2113 	:	val_out <= 16'hb9bc;
             14'h2114 	:	val_out <= 16'hb9c0;
             14'h2115 	:	val_out <= 16'hb9c5;
             14'h2116 	:	val_out <= 16'hb9c9;
             14'h2117 	:	val_out <= 16'hb9cd;
             14'h2118 	:	val_out <= 16'hb9d2;
             14'h2119 	:	val_out <= 16'hb9d6;
             14'h211a 	:	val_out <= 16'hb9da;
             14'h211b 	:	val_out <= 16'hb9df;
             14'h211c 	:	val_out <= 16'hb9e3;
             14'h211d 	:	val_out <= 16'hb9e7;
             14'h211e 	:	val_out <= 16'hb9ec;
             14'h211f 	:	val_out <= 16'hb9f0;
             14'h2120 	:	val_out <= 16'hb9f4;
             14'h2121 	:	val_out <= 16'hb9f9;
             14'h2122 	:	val_out <= 16'hb9fd;
             14'h2123 	:	val_out <= 16'hba01;
             14'h2124 	:	val_out <= 16'hba06;
             14'h2125 	:	val_out <= 16'hba0a;
             14'h2126 	:	val_out <= 16'hba0e;
             14'h2127 	:	val_out <= 16'hba13;
             14'h2128 	:	val_out <= 16'hba17;
             14'h2129 	:	val_out <= 16'hba1b;
             14'h212a 	:	val_out <= 16'hba1f;
             14'h212b 	:	val_out <= 16'hba24;
             14'h212c 	:	val_out <= 16'hba28;
             14'h212d 	:	val_out <= 16'hba2c;
             14'h212e 	:	val_out <= 16'hba31;
             14'h212f 	:	val_out <= 16'hba35;
             14'h2130 	:	val_out <= 16'hba39;
             14'h2131 	:	val_out <= 16'hba3e;
             14'h2132 	:	val_out <= 16'hba42;
             14'h2133 	:	val_out <= 16'hba46;
             14'h2134 	:	val_out <= 16'hba4b;
             14'h2135 	:	val_out <= 16'hba4f;
             14'h2136 	:	val_out <= 16'hba53;
             14'h2137 	:	val_out <= 16'hba58;
             14'h2138 	:	val_out <= 16'hba5c;
             14'h2139 	:	val_out <= 16'hba60;
             14'h213a 	:	val_out <= 16'hba64;
             14'h213b 	:	val_out <= 16'hba69;
             14'h213c 	:	val_out <= 16'hba6d;
             14'h213d 	:	val_out <= 16'hba71;
             14'h213e 	:	val_out <= 16'hba76;
             14'h213f 	:	val_out <= 16'hba7a;
             14'h2140 	:	val_out <= 16'hba7e;
             14'h2141 	:	val_out <= 16'hba83;
             14'h2142 	:	val_out <= 16'hba87;
             14'h2143 	:	val_out <= 16'hba8b;
             14'h2144 	:	val_out <= 16'hba90;
             14'h2145 	:	val_out <= 16'hba94;
             14'h2146 	:	val_out <= 16'hba98;
             14'h2147 	:	val_out <= 16'hba9c;
             14'h2148 	:	val_out <= 16'hbaa1;
             14'h2149 	:	val_out <= 16'hbaa5;
             14'h214a 	:	val_out <= 16'hbaa9;
             14'h214b 	:	val_out <= 16'hbaae;
             14'h214c 	:	val_out <= 16'hbab2;
             14'h214d 	:	val_out <= 16'hbab6;
             14'h214e 	:	val_out <= 16'hbabb;
             14'h214f 	:	val_out <= 16'hbabf;
             14'h2150 	:	val_out <= 16'hbac3;
             14'h2151 	:	val_out <= 16'hbac7;
             14'h2152 	:	val_out <= 16'hbacc;
             14'h2153 	:	val_out <= 16'hbad0;
             14'h2154 	:	val_out <= 16'hbad4;
             14'h2155 	:	val_out <= 16'hbad9;
             14'h2156 	:	val_out <= 16'hbadd;
             14'h2157 	:	val_out <= 16'hbae1;
             14'h2158 	:	val_out <= 16'hbae5;
             14'h2159 	:	val_out <= 16'hbaea;
             14'h215a 	:	val_out <= 16'hbaee;
             14'h215b 	:	val_out <= 16'hbaf2;
             14'h215c 	:	val_out <= 16'hbaf7;
             14'h215d 	:	val_out <= 16'hbafb;
             14'h215e 	:	val_out <= 16'hbaff;
             14'h215f 	:	val_out <= 16'hbb04;
             14'h2160 	:	val_out <= 16'hbb08;
             14'h2161 	:	val_out <= 16'hbb0c;
             14'h2162 	:	val_out <= 16'hbb10;
             14'h2163 	:	val_out <= 16'hbb15;
             14'h2164 	:	val_out <= 16'hbb19;
             14'h2165 	:	val_out <= 16'hbb1d;
             14'h2166 	:	val_out <= 16'hbb22;
             14'h2167 	:	val_out <= 16'hbb26;
             14'h2168 	:	val_out <= 16'hbb2a;
             14'h2169 	:	val_out <= 16'hbb2e;
             14'h216a 	:	val_out <= 16'hbb33;
             14'h216b 	:	val_out <= 16'hbb37;
             14'h216c 	:	val_out <= 16'hbb3b;
             14'h216d 	:	val_out <= 16'hbb40;
             14'h216e 	:	val_out <= 16'hbb44;
             14'h216f 	:	val_out <= 16'hbb48;
             14'h2170 	:	val_out <= 16'hbb4c;
             14'h2171 	:	val_out <= 16'hbb51;
             14'h2172 	:	val_out <= 16'hbb55;
             14'h2173 	:	val_out <= 16'hbb59;
             14'h2174 	:	val_out <= 16'hbb5e;
             14'h2175 	:	val_out <= 16'hbb62;
             14'h2176 	:	val_out <= 16'hbb66;
             14'h2177 	:	val_out <= 16'hbb6a;
             14'h2178 	:	val_out <= 16'hbb6f;
             14'h2179 	:	val_out <= 16'hbb73;
             14'h217a 	:	val_out <= 16'hbb77;
             14'h217b 	:	val_out <= 16'hbb7b;
             14'h217c 	:	val_out <= 16'hbb80;
             14'h217d 	:	val_out <= 16'hbb84;
             14'h217e 	:	val_out <= 16'hbb88;
             14'h217f 	:	val_out <= 16'hbb8d;
             14'h2180 	:	val_out <= 16'hbb91;
             14'h2181 	:	val_out <= 16'hbb95;
             14'h2182 	:	val_out <= 16'hbb99;
             14'h2183 	:	val_out <= 16'hbb9e;
             14'h2184 	:	val_out <= 16'hbba2;
             14'h2185 	:	val_out <= 16'hbba6;
             14'h2186 	:	val_out <= 16'hbbab;
             14'h2187 	:	val_out <= 16'hbbaf;
             14'h2188 	:	val_out <= 16'hbbb3;
             14'h2189 	:	val_out <= 16'hbbb7;
             14'h218a 	:	val_out <= 16'hbbbc;
             14'h218b 	:	val_out <= 16'hbbc0;
             14'h218c 	:	val_out <= 16'hbbc4;
             14'h218d 	:	val_out <= 16'hbbc8;
             14'h218e 	:	val_out <= 16'hbbcd;
             14'h218f 	:	val_out <= 16'hbbd1;
             14'h2190 	:	val_out <= 16'hbbd5;
             14'h2191 	:	val_out <= 16'hbbd9;
             14'h2192 	:	val_out <= 16'hbbde;
             14'h2193 	:	val_out <= 16'hbbe2;
             14'h2194 	:	val_out <= 16'hbbe6;
             14'h2195 	:	val_out <= 16'hbbeb;
             14'h2196 	:	val_out <= 16'hbbef;
             14'h2197 	:	val_out <= 16'hbbf3;
             14'h2198 	:	val_out <= 16'hbbf7;
             14'h2199 	:	val_out <= 16'hbbfc;
             14'h219a 	:	val_out <= 16'hbc00;
             14'h219b 	:	val_out <= 16'hbc04;
             14'h219c 	:	val_out <= 16'hbc08;
             14'h219d 	:	val_out <= 16'hbc0d;
             14'h219e 	:	val_out <= 16'hbc11;
             14'h219f 	:	val_out <= 16'hbc15;
             14'h21a0 	:	val_out <= 16'hbc19;
             14'h21a1 	:	val_out <= 16'hbc1e;
             14'h21a2 	:	val_out <= 16'hbc22;
             14'h21a3 	:	val_out <= 16'hbc26;
             14'h21a4 	:	val_out <= 16'hbc2b;
             14'h21a5 	:	val_out <= 16'hbc2f;
             14'h21a6 	:	val_out <= 16'hbc33;
             14'h21a7 	:	val_out <= 16'hbc37;
             14'h21a8 	:	val_out <= 16'hbc3c;
             14'h21a9 	:	val_out <= 16'hbc40;
             14'h21aa 	:	val_out <= 16'hbc44;
             14'h21ab 	:	val_out <= 16'hbc48;
             14'h21ac 	:	val_out <= 16'hbc4d;
             14'h21ad 	:	val_out <= 16'hbc51;
             14'h21ae 	:	val_out <= 16'hbc55;
             14'h21af 	:	val_out <= 16'hbc59;
             14'h21b0 	:	val_out <= 16'hbc5e;
             14'h21b1 	:	val_out <= 16'hbc62;
             14'h21b2 	:	val_out <= 16'hbc66;
             14'h21b3 	:	val_out <= 16'hbc6a;
             14'h21b4 	:	val_out <= 16'hbc6f;
             14'h21b5 	:	val_out <= 16'hbc73;
             14'h21b6 	:	val_out <= 16'hbc77;
             14'h21b7 	:	val_out <= 16'hbc7b;
             14'h21b8 	:	val_out <= 16'hbc80;
             14'h21b9 	:	val_out <= 16'hbc84;
             14'h21ba 	:	val_out <= 16'hbc88;
             14'h21bb 	:	val_out <= 16'hbc8c;
             14'h21bc 	:	val_out <= 16'hbc91;
             14'h21bd 	:	val_out <= 16'hbc95;
             14'h21be 	:	val_out <= 16'hbc99;
             14'h21bf 	:	val_out <= 16'hbc9d;
             14'h21c0 	:	val_out <= 16'hbca2;
             14'h21c1 	:	val_out <= 16'hbca6;
             14'h21c2 	:	val_out <= 16'hbcaa;
             14'h21c3 	:	val_out <= 16'hbcae;
             14'h21c4 	:	val_out <= 16'hbcb3;
             14'h21c5 	:	val_out <= 16'hbcb7;
             14'h21c6 	:	val_out <= 16'hbcbb;
             14'h21c7 	:	val_out <= 16'hbcbf;
             14'h21c8 	:	val_out <= 16'hbcc4;
             14'h21c9 	:	val_out <= 16'hbcc8;
             14'h21ca 	:	val_out <= 16'hbccc;
             14'h21cb 	:	val_out <= 16'hbcd0;
             14'h21cc 	:	val_out <= 16'hbcd5;
             14'h21cd 	:	val_out <= 16'hbcd9;
             14'h21ce 	:	val_out <= 16'hbcdd;
             14'h21cf 	:	val_out <= 16'hbce1;
             14'h21d0 	:	val_out <= 16'hbce6;
             14'h21d1 	:	val_out <= 16'hbcea;
             14'h21d2 	:	val_out <= 16'hbcee;
             14'h21d3 	:	val_out <= 16'hbcf2;
             14'h21d4 	:	val_out <= 16'hbcf7;
             14'h21d5 	:	val_out <= 16'hbcfb;
             14'h21d6 	:	val_out <= 16'hbcff;
             14'h21d7 	:	val_out <= 16'hbd03;
             14'h21d8 	:	val_out <= 16'hbd07;
             14'h21d9 	:	val_out <= 16'hbd0c;
             14'h21da 	:	val_out <= 16'hbd10;
             14'h21db 	:	val_out <= 16'hbd14;
             14'h21dc 	:	val_out <= 16'hbd18;
             14'h21dd 	:	val_out <= 16'hbd1d;
             14'h21de 	:	val_out <= 16'hbd21;
             14'h21df 	:	val_out <= 16'hbd25;
             14'h21e0 	:	val_out <= 16'hbd29;
             14'h21e1 	:	val_out <= 16'hbd2e;
             14'h21e2 	:	val_out <= 16'hbd32;
             14'h21e3 	:	val_out <= 16'hbd36;
             14'h21e4 	:	val_out <= 16'hbd3a;
             14'h21e5 	:	val_out <= 16'hbd3e;
             14'h21e6 	:	val_out <= 16'hbd43;
             14'h21e7 	:	val_out <= 16'hbd47;
             14'h21e8 	:	val_out <= 16'hbd4b;
             14'h21e9 	:	val_out <= 16'hbd4f;
             14'h21ea 	:	val_out <= 16'hbd54;
             14'h21eb 	:	val_out <= 16'hbd58;
             14'h21ec 	:	val_out <= 16'hbd5c;
             14'h21ed 	:	val_out <= 16'hbd60;
             14'h21ee 	:	val_out <= 16'hbd65;
             14'h21ef 	:	val_out <= 16'hbd69;
             14'h21f0 	:	val_out <= 16'hbd6d;
             14'h21f1 	:	val_out <= 16'hbd71;
             14'h21f2 	:	val_out <= 16'hbd75;
             14'h21f3 	:	val_out <= 16'hbd7a;
             14'h21f4 	:	val_out <= 16'hbd7e;
             14'h21f5 	:	val_out <= 16'hbd82;
             14'h21f6 	:	val_out <= 16'hbd86;
             14'h21f7 	:	val_out <= 16'hbd8b;
             14'h21f8 	:	val_out <= 16'hbd8f;
             14'h21f9 	:	val_out <= 16'hbd93;
             14'h21fa 	:	val_out <= 16'hbd97;
             14'h21fb 	:	val_out <= 16'hbd9b;
             14'h21fc 	:	val_out <= 16'hbda0;
             14'h21fd 	:	val_out <= 16'hbda4;
             14'h21fe 	:	val_out <= 16'hbda8;
             14'h21ff 	:	val_out <= 16'hbdac;
             14'h2200 	:	val_out <= 16'hbdb1;
             14'h2201 	:	val_out <= 16'hbdb5;
             14'h2202 	:	val_out <= 16'hbdb9;
             14'h2203 	:	val_out <= 16'hbdbd;
             14'h2204 	:	val_out <= 16'hbdc1;
             14'h2205 	:	val_out <= 16'hbdc6;
             14'h2206 	:	val_out <= 16'hbdca;
             14'h2207 	:	val_out <= 16'hbdce;
             14'h2208 	:	val_out <= 16'hbdd2;
             14'h2209 	:	val_out <= 16'hbdd7;
             14'h220a 	:	val_out <= 16'hbddb;
             14'h220b 	:	val_out <= 16'hbddf;
             14'h220c 	:	val_out <= 16'hbde3;
             14'h220d 	:	val_out <= 16'hbde7;
             14'h220e 	:	val_out <= 16'hbdec;
             14'h220f 	:	val_out <= 16'hbdf0;
             14'h2210 	:	val_out <= 16'hbdf4;
             14'h2211 	:	val_out <= 16'hbdf8;
             14'h2212 	:	val_out <= 16'hbdfc;
             14'h2213 	:	val_out <= 16'hbe01;
             14'h2214 	:	val_out <= 16'hbe05;
             14'h2215 	:	val_out <= 16'hbe09;
             14'h2216 	:	val_out <= 16'hbe0d;
             14'h2217 	:	val_out <= 16'hbe12;
             14'h2218 	:	val_out <= 16'hbe16;
             14'h2219 	:	val_out <= 16'hbe1a;
             14'h221a 	:	val_out <= 16'hbe1e;
             14'h221b 	:	val_out <= 16'hbe22;
             14'h221c 	:	val_out <= 16'hbe27;
             14'h221d 	:	val_out <= 16'hbe2b;
             14'h221e 	:	val_out <= 16'hbe2f;
             14'h221f 	:	val_out <= 16'hbe33;
             14'h2220 	:	val_out <= 16'hbe37;
             14'h2221 	:	val_out <= 16'hbe3c;
             14'h2222 	:	val_out <= 16'hbe40;
             14'h2223 	:	val_out <= 16'hbe44;
             14'h2224 	:	val_out <= 16'hbe48;
             14'h2225 	:	val_out <= 16'hbe4c;
             14'h2226 	:	val_out <= 16'hbe51;
             14'h2227 	:	val_out <= 16'hbe55;
             14'h2228 	:	val_out <= 16'hbe59;
             14'h2229 	:	val_out <= 16'hbe5d;
             14'h222a 	:	val_out <= 16'hbe61;
             14'h222b 	:	val_out <= 16'hbe66;
             14'h222c 	:	val_out <= 16'hbe6a;
             14'h222d 	:	val_out <= 16'hbe6e;
             14'h222e 	:	val_out <= 16'hbe72;
             14'h222f 	:	val_out <= 16'hbe76;
             14'h2230 	:	val_out <= 16'hbe7b;
             14'h2231 	:	val_out <= 16'hbe7f;
             14'h2232 	:	val_out <= 16'hbe83;
             14'h2233 	:	val_out <= 16'hbe87;
             14'h2234 	:	val_out <= 16'hbe8b;
             14'h2235 	:	val_out <= 16'hbe90;
             14'h2236 	:	val_out <= 16'hbe94;
             14'h2237 	:	val_out <= 16'hbe98;
             14'h2238 	:	val_out <= 16'hbe9c;
             14'h2239 	:	val_out <= 16'hbea0;
             14'h223a 	:	val_out <= 16'hbea5;
             14'h223b 	:	val_out <= 16'hbea9;
             14'h223c 	:	val_out <= 16'hbead;
             14'h223d 	:	val_out <= 16'hbeb1;
             14'h223e 	:	val_out <= 16'hbeb5;
             14'h223f 	:	val_out <= 16'hbeba;
             14'h2240 	:	val_out <= 16'hbebe;
             14'h2241 	:	val_out <= 16'hbec2;
             14'h2242 	:	val_out <= 16'hbec6;
             14'h2243 	:	val_out <= 16'hbeca;
             14'h2244 	:	val_out <= 16'hbece;
             14'h2245 	:	val_out <= 16'hbed3;
             14'h2246 	:	val_out <= 16'hbed7;
             14'h2247 	:	val_out <= 16'hbedb;
             14'h2248 	:	val_out <= 16'hbedf;
             14'h2249 	:	val_out <= 16'hbee3;
             14'h224a 	:	val_out <= 16'hbee8;
             14'h224b 	:	val_out <= 16'hbeec;
             14'h224c 	:	val_out <= 16'hbef0;
             14'h224d 	:	val_out <= 16'hbef4;
             14'h224e 	:	val_out <= 16'hbef8;
             14'h224f 	:	val_out <= 16'hbefd;
             14'h2250 	:	val_out <= 16'hbf01;
             14'h2251 	:	val_out <= 16'hbf05;
             14'h2252 	:	val_out <= 16'hbf09;
             14'h2253 	:	val_out <= 16'hbf0d;
             14'h2254 	:	val_out <= 16'hbf11;
             14'h2255 	:	val_out <= 16'hbf16;
             14'h2256 	:	val_out <= 16'hbf1a;
             14'h2257 	:	val_out <= 16'hbf1e;
             14'h2258 	:	val_out <= 16'hbf22;
             14'h2259 	:	val_out <= 16'hbf26;
             14'h225a 	:	val_out <= 16'hbf2b;
             14'h225b 	:	val_out <= 16'hbf2f;
             14'h225c 	:	val_out <= 16'hbf33;
             14'h225d 	:	val_out <= 16'hbf37;
             14'h225e 	:	val_out <= 16'hbf3b;
             14'h225f 	:	val_out <= 16'hbf3f;
             14'h2260 	:	val_out <= 16'hbf44;
             14'h2261 	:	val_out <= 16'hbf48;
             14'h2262 	:	val_out <= 16'hbf4c;
             14'h2263 	:	val_out <= 16'hbf50;
             14'h2264 	:	val_out <= 16'hbf54;
             14'h2265 	:	val_out <= 16'hbf58;
             14'h2266 	:	val_out <= 16'hbf5d;
             14'h2267 	:	val_out <= 16'hbf61;
             14'h2268 	:	val_out <= 16'hbf65;
             14'h2269 	:	val_out <= 16'hbf69;
             14'h226a 	:	val_out <= 16'hbf6d;
             14'h226b 	:	val_out <= 16'hbf71;
             14'h226c 	:	val_out <= 16'hbf76;
             14'h226d 	:	val_out <= 16'hbf7a;
             14'h226e 	:	val_out <= 16'hbf7e;
             14'h226f 	:	val_out <= 16'hbf82;
             14'h2270 	:	val_out <= 16'hbf86;
             14'h2271 	:	val_out <= 16'hbf8b;
             14'h2272 	:	val_out <= 16'hbf8f;
             14'h2273 	:	val_out <= 16'hbf93;
             14'h2274 	:	val_out <= 16'hbf97;
             14'h2275 	:	val_out <= 16'hbf9b;
             14'h2276 	:	val_out <= 16'hbf9f;
             14'h2277 	:	val_out <= 16'hbfa4;
             14'h2278 	:	val_out <= 16'hbfa8;
             14'h2279 	:	val_out <= 16'hbfac;
             14'h227a 	:	val_out <= 16'hbfb0;
             14'h227b 	:	val_out <= 16'hbfb4;
             14'h227c 	:	val_out <= 16'hbfb8;
             14'h227d 	:	val_out <= 16'hbfbc;
             14'h227e 	:	val_out <= 16'hbfc1;
             14'h227f 	:	val_out <= 16'hbfc5;
             14'h2280 	:	val_out <= 16'hbfc9;
             14'h2281 	:	val_out <= 16'hbfcd;
             14'h2282 	:	val_out <= 16'hbfd1;
             14'h2283 	:	val_out <= 16'hbfd5;
             14'h2284 	:	val_out <= 16'hbfda;
             14'h2285 	:	val_out <= 16'hbfde;
             14'h2286 	:	val_out <= 16'hbfe2;
             14'h2287 	:	val_out <= 16'hbfe6;
             14'h2288 	:	val_out <= 16'hbfea;
             14'h2289 	:	val_out <= 16'hbfee;
             14'h228a 	:	val_out <= 16'hbff3;
             14'h228b 	:	val_out <= 16'hbff7;
             14'h228c 	:	val_out <= 16'hbffb;
             14'h228d 	:	val_out <= 16'hbfff;
             14'h228e 	:	val_out <= 16'hc003;
             14'h228f 	:	val_out <= 16'hc007;
             14'h2290 	:	val_out <= 16'hc00c;
             14'h2291 	:	val_out <= 16'hc010;
             14'h2292 	:	val_out <= 16'hc014;
             14'h2293 	:	val_out <= 16'hc018;
             14'h2294 	:	val_out <= 16'hc01c;
             14'h2295 	:	val_out <= 16'hc020;
             14'h2296 	:	val_out <= 16'hc024;
             14'h2297 	:	val_out <= 16'hc029;
             14'h2298 	:	val_out <= 16'hc02d;
             14'h2299 	:	val_out <= 16'hc031;
             14'h229a 	:	val_out <= 16'hc035;
             14'h229b 	:	val_out <= 16'hc039;
             14'h229c 	:	val_out <= 16'hc03d;
             14'h229d 	:	val_out <= 16'hc041;
             14'h229e 	:	val_out <= 16'hc046;
             14'h229f 	:	val_out <= 16'hc04a;
             14'h22a0 	:	val_out <= 16'hc04e;
             14'h22a1 	:	val_out <= 16'hc052;
             14'h22a2 	:	val_out <= 16'hc056;
             14'h22a3 	:	val_out <= 16'hc05a;
             14'h22a4 	:	val_out <= 16'hc05f;
             14'h22a5 	:	val_out <= 16'hc063;
             14'h22a6 	:	val_out <= 16'hc067;
             14'h22a7 	:	val_out <= 16'hc06b;
             14'h22a8 	:	val_out <= 16'hc06f;
             14'h22a9 	:	val_out <= 16'hc073;
             14'h22aa 	:	val_out <= 16'hc077;
             14'h22ab 	:	val_out <= 16'hc07c;
             14'h22ac 	:	val_out <= 16'hc080;
             14'h22ad 	:	val_out <= 16'hc084;
             14'h22ae 	:	val_out <= 16'hc088;
             14'h22af 	:	val_out <= 16'hc08c;
             14'h22b0 	:	val_out <= 16'hc090;
             14'h22b1 	:	val_out <= 16'hc094;
             14'h22b2 	:	val_out <= 16'hc099;
             14'h22b3 	:	val_out <= 16'hc09d;
             14'h22b4 	:	val_out <= 16'hc0a1;
             14'h22b5 	:	val_out <= 16'hc0a5;
             14'h22b6 	:	val_out <= 16'hc0a9;
             14'h22b7 	:	val_out <= 16'hc0ad;
             14'h22b8 	:	val_out <= 16'hc0b1;
             14'h22b9 	:	val_out <= 16'hc0b5;
             14'h22ba 	:	val_out <= 16'hc0ba;
             14'h22bb 	:	val_out <= 16'hc0be;
             14'h22bc 	:	val_out <= 16'hc0c2;
             14'h22bd 	:	val_out <= 16'hc0c6;
             14'h22be 	:	val_out <= 16'hc0ca;
             14'h22bf 	:	val_out <= 16'hc0ce;
             14'h22c0 	:	val_out <= 16'hc0d2;
             14'h22c1 	:	val_out <= 16'hc0d7;
             14'h22c2 	:	val_out <= 16'hc0db;
             14'h22c3 	:	val_out <= 16'hc0df;
             14'h22c4 	:	val_out <= 16'hc0e3;
             14'h22c5 	:	val_out <= 16'hc0e7;
             14'h22c6 	:	val_out <= 16'hc0eb;
             14'h22c7 	:	val_out <= 16'hc0ef;
             14'h22c8 	:	val_out <= 16'hc0f3;
             14'h22c9 	:	val_out <= 16'hc0f8;
             14'h22ca 	:	val_out <= 16'hc0fc;
             14'h22cb 	:	val_out <= 16'hc100;
             14'h22cc 	:	val_out <= 16'hc104;
             14'h22cd 	:	val_out <= 16'hc108;
             14'h22ce 	:	val_out <= 16'hc10c;
             14'h22cf 	:	val_out <= 16'hc110;
             14'h22d0 	:	val_out <= 16'hc114;
             14'h22d1 	:	val_out <= 16'hc119;
             14'h22d2 	:	val_out <= 16'hc11d;
             14'h22d3 	:	val_out <= 16'hc121;
             14'h22d4 	:	val_out <= 16'hc125;
             14'h22d5 	:	val_out <= 16'hc129;
             14'h22d6 	:	val_out <= 16'hc12d;
             14'h22d7 	:	val_out <= 16'hc131;
             14'h22d8 	:	val_out <= 16'hc135;
             14'h22d9 	:	val_out <= 16'hc13a;
             14'h22da 	:	val_out <= 16'hc13e;
             14'h22db 	:	val_out <= 16'hc142;
             14'h22dc 	:	val_out <= 16'hc146;
             14'h22dd 	:	val_out <= 16'hc14a;
             14'h22de 	:	val_out <= 16'hc14e;
             14'h22df 	:	val_out <= 16'hc152;
             14'h22e0 	:	val_out <= 16'hc156;
             14'h22e1 	:	val_out <= 16'hc15b;
             14'h22e2 	:	val_out <= 16'hc15f;
             14'h22e3 	:	val_out <= 16'hc163;
             14'h22e4 	:	val_out <= 16'hc167;
             14'h22e5 	:	val_out <= 16'hc16b;
             14'h22e6 	:	val_out <= 16'hc16f;
             14'h22e7 	:	val_out <= 16'hc173;
             14'h22e8 	:	val_out <= 16'hc177;
             14'h22e9 	:	val_out <= 16'hc17b;
             14'h22ea 	:	val_out <= 16'hc180;
             14'h22eb 	:	val_out <= 16'hc184;
             14'h22ec 	:	val_out <= 16'hc188;
             14'h22ed 	:	val_out <= 16'hc18c;
             14'h22ee 	:	val_out <= 16'hc190;
             14'h22ef 	:	val_out <= 16'hc194;
             14'h22f0 	:	val_out <= 16'hc198;
             14'h22f1 	:	val_out <= 16'hc19c;
             14'h22f2 	:	val_out <= 16'hc1a0;
             14'h22f3 	:	val_out <= 16'hc1a5;
             14'h22f4 	:	val_out <= 16'hc1a9;
             14'h22f5 	:	val_out <= 16'hc1ad;
             14'h22f6 	:	val_out <= 16'hc1b1;
             14'h22f7 	:	val_out <= 16'hc1b5;
             14'h22f8 	:	val_out <= 16'hc1b9;
             14'h22f9 	:	val_out <= 16'hc1bd;
             14'h22fa 	:	val_out <= 16'hc1c1;
             14'h22fb 	:	val_out <= 16'hc1c5;
             14'h22fc 	:	val_out <= 16'hc1ca;
             14'h22fd 	:	val_out <= 16'hc1ce;
             14'h22fe 	:	val_out <= 16'hc1d2;
             14'h22ff 	:	val_out <= 16'hc1d6;
             14'h2300 	:	val_out <= 16'hc1da;
             14'h2301 	:	val_out <= 16'hc1de;
             14'h2302 	:	val_out <= 16'hc1e2;
             14'h2303 	:	val_out <= 16'hc1e6;
             14'h2304 	:	val_out <= 16'hc1ea;
             14'h2305 	:	val_out <= 16'hc1ef;
             14'h2306 	:	val_out <= 16'hc1f3;
             14'h2307 	:	val_out <= 16'hc1f7;
             14'h2308 	:	val_out <= 16'hc1fb;
             14'h2309 	:	val_out <= 16'hc1ff;
             14'h230a 	:	val_out <= 16'hc203;
             14'h230b 	:	val_out <= 16'hc207;
             14'h230c 	:	val_out <= 16'hc20b;
             14'h230d 	:	val_out <= 16'hc20f;
             14'h230e 	:	val_out <= 16'hc213;
             14'h230f 	:	val_out <= 16'hc217;
             14'h2310 	:	val_out <= 16'hc21c;
             14'h2311 	:	val_out <= 16'hc220;
             14'h2312 	:	val_out <= 16'hc224;
             14'h2313 	:	val_out <= 16'hc228;
             14'h2314 	:	val_out <= 16'hc22c;
             14'h2315 	:	val_out <= 16'hc230;
             14'h2316 	:	val_out <= 16'hc234;
             14'h2317 	:	val_out <= 16'hc238;
             14'h2318 	:	val_out <= 16'hc23c;
             14'h2319 	:	val_out <= 16'hc240;
             14'h231a 	:	val_out <= 16'hc245;
             14'h231b 	:	val_out <= 16'hc249;
             14'h231c 	:	val_out <= 16'hc24d;
             14'h231d 	:	val_out <= 16'hc251;
             14'h231e 	:	val_out <= 16'hc255;
             14'h231f 	:	val_out <= 16'hc259;
             14'h2320 	:	val_out <= 16'hc25d;
             14'h2321 	:	val_out <= 16'hc261;
             14'h2322 	:	val_out <= 16'hc265;
             14'h2323 	:	val_out <= 16'hc269;
             14'h2324 	:	val_out <= 16'hc26d;
             14'h2325 	:	val_out <= 16'hc272;
             14'h2326 	:	val_out <= 16'hc276;
             14'h2327 	:	val_out <= 16'hc27a;
             14'h2328 	:	val_out <= 16'hc27e;
             14'h2329 	:	val_out <= 16'hc282;
             14'h232a 	:	val_out <= 16'hc286;
             14'h232b 	:	val_out <= 16'hc28a;
             14'h232c 	:	val_out <= 16'hc28e;
             14'h232d 	:	val_out <= 16'hc292;
             14'h232e 	:	val_out <= 16'hc296;
             14'h232f 	:	val_out <= 16'hc29a;
             14'h2330 	:	val_out <= 16'hc29e;
             14'h2331 	:	val_out <= 16'hc2a3;
             14'h2332 	:	val_out <= 16'hc2a7;
             14'h2333 	:	val_out <= 16'hc2ab;
             14'h2334 	:	val_out <= 16'hc2af;
             14'h2335 	:	val_out <= 16'hc2b3;
             14'h2336 	:	val_out <= 16'hc2b7;
             14'h2337 	:	val_out <= 16'hc2bb;
             14'h2338 	:	val_out <= 16'hc2bf;
             14'h2339 	:	val_out <= 16'hc2c3;
             14'h233a 	:	val_out <= 16'hc2c7;
             14'h233b 	:	val_out <= 16'hc2cb;
             14'h233c 	:	val_out <= 16'hc2cf;
             14'h233d 	:	val_out <= 16'hc2d3;
             14'h233e 	:	val_out <= 16'hc2d8;
             14'h233f 	:	val_out <= 16'hc2dc;
             14'h2340 	:	val_out <= 16'hc2e0;
             14'h2341 	:	val_out <= 16'hc2e4;
             14'h2342 	:	val_out <= 16'hc2e8;
             14'h2343 	:	val_out <= 16'hc2ec;
             14'h2344 	:	val_out <= 16'hc2f0;
             14'h2345 	:	val_out <= 16'hc2f4;
             14'h2346 	:	val_out <= 16'hc2f8;
             14'h2347 	:	val_out <= 16'hc2fc;
             14'h2348 	:	val_out <= 16'hc300;
             14'h2349 	:	val_out <= 16'hc304;
             14'h234a 	:	val_out <= 16'hc308;
             14'h234b 	:	val_out <= 16'hc30c;
             14'h234c 	:	val_out <= 16'hc311;
             14'h234d 	:	val_out <= 16'hc315;
             14'h234e 	:	val_out <= 16'hc319;
             14'h234f 	:	val_out <= 16'hc31d;
             14'h2350 	:	val_out <= 16'hc321;
             14'h2351 	:	val_out <= 16'hc325;
             14'h2352 	:	val_out <= 16'hc329;
             14'h2353 	:	val_out <= 16'hc32d;
             14'h2354 	:	val_out <= 16'hc331;
             14'h2355 	:	val_out <= 16'hc335;
             14'h2356 	:	val_out <= 16'hc339;
             14'h2357 	:	val_out <= 16'hc33d;
             14'h2358 	:	val_out <= 16'hc341;
             14'h2359 	:	val_out <= 16'hc345;
             14'h235a 	:	val_out <= 16'hc349;
             14'h235b 	:	val_out <= 16'hc34e;
             14'h235c 	:	val_out <= 16'hc352;
             14'h235d 	:	val_out <= 16'hc356;
             14'h235e 	:	val_out <= 16'hc35a;
             14'h235f 	:	val_out <= 16'hc35e;
             14'h2360 	:	val_out <= 16'hc362;
             14'h2361 	:	val_out <= 16'hc366;
             14'h2362 	:	val_out <= 16'hc36a;
             14'h2363 	:	val_out <= 16'hc36e;
             14'h2364 	:	val_out <= 16'hc372;
             14'h2365 	:	val_out <= 16'hc376;
             14'h2366 	:	val_out <= 16'hc37a;
             14'h2367 	:	val_out <= 16'hc37e;
             14'h2368 	:	val_out <= 16'hc382;
             14'h2369 	:	val_out <= 16'hc386;
             14'h236a 	:	val_out <= 16'hc38a;
             14'h236b 	:	val_out <= 16'hc38e;
             14'h236c 	:	val_out <= 16'hc393;
             14'h236d 	:	val_out <= 16'hc397;
             14'h236e 	:	val_out <= 16'hc39b;
             14'h236f 	:	val_out <= 16'hc39f;
             14'h2370 	:	val_out <= 16'hc3a3;
             14'h2371 	:	val_out <= 16'hc3a7;
             14'h2372 	:	val_out <= 16'hc3ab;
             14'h2373 	:	val_out <= 16'hc3af;
             14'h2374 	:	val_out <= 16'hc3b3;
             14'h2375 	:	val_out <= 16'hc3b7;
             14'h2376 	:	val_out <= 16'hc3bb;
             14'h2377 	:	val_out <= 16'hc3bf;
             14'h2378 	:	val_out <= 16'hc3c3;
             14'h2379 	:	val_out <= 16'hc3c7;
             14'h237a 	:	val_out <= 16'hc3cb;
             14'h237b 	:	val_out <= 16'hc3cf;
             14'h237c 	:	val_out <= 16'hc3d3;
             14'h237d 	:	val_out <= 16'hc3d7;
             14'h237e 	:	val_out <= 16'hc3db;
             14'h237f 	:	val_out <= 16'hc3df;
             14'h2380 	:	val_out <= 16'hc3e4;
             14'h2381 	:	val_out <= 16'hc3e8;
             14'h2382 	:	val_out <= 16'hc3ec;
             14'h2383 	:	val_out <= 16'hc3f0;
             14'h2384 	:	val_out <= 16'hc3f4;
             14'h2385 	:	val_out <= 16'hc3f8;
             14'h2386 	:	val_out <= 16'hc3fc;
             14'h2387 	:	val_out <= 16'hc400;
             14'h2388 	:	val_out <= 16'hc404;
             14'h2389 	:	val_out <= 16'hc408;
             14'h238a 	:	val_out <= 16'hc40c;
             14'h238b 	:	val_out <= 16'hc410;
             14'h238c 	:	val_out <= 16'hc414;
             14'h238d 	:	val_out <= 16'hc418;
             14'h238e 	:	val_out <= 16'hc41c;
             14'h238f 	:	val_out <= 16'hc420;
             14'h2390 	:	val_out <= 16'hc424;
             14'h2391 	:	val_out <= 16'hc428;
             14'h2392 	:	val_out <= 16'hc42c;
             14'h2393 	:	val_out <= 16'hc430;
             14'h2394 	:	val_out <= 16'hc434;
             14'h2395 	:	val_out <= 16'hc438;
             14'h2396 	:	val_out <= 16'hc43c;
             14'h2397 	:	val_out <= 16'hc440;
             14'h2398 	:	val_out <= 16'hc444;
             14'h2399 	:	val_out <= 16'hc449;
             14'h239a 	:	val_out <= 16'hc44d;
             14'h239b 	:	val_out <= 16'hc451;
             14'h239c 	:	val_out <= 16'hc455;
             14'h239d 	:	val_out <= 16'hc459;
             14'h239e 	:	val_out <= 16'hc45d;
             14'h239f 	:	val_out <= 16'hc461;
             14'h23a0 	:	val_out <= 16'hc465;
             14'h23a1 	:	val_out <= 16'hc469;
             14'h23a2 	:	val_out <= 16'hc46d;
             14'h23a3 	:	val_out <= 16'hc471;
             14'h23a4 	:	val_out <= 16'hc475;
             14'h23a5 	:	val_out <= 16'hc479;
             14'h23a6 	:	val_out <= 16'hc47d;
             14'h23a7 	:	val_out <= 16'hc481;
             14'h23a8 	:	val_out <= 16'hc485;
             14'h23a9 	:	val_out <= 16'hc489;
             14'h23aa 	:	val_out <= 16'hc48d;
             14'h23ab 	:	val_out <= 16'hc491;
             14'h23ac 	:	val_out <= 16'hc495;
             14'h23ad 	:	val_out <= 16'hc499;
             14'h23ae 	:	val_out <= 16'hc49d;
             14'h23af 	:	val_out <= 16'hc4a1;
             14'h23b0 	:	val_out <= 16'hc4a5;
             14'h23b1 	:	val_out <= 16'hc4a9;
             14'h23b2 	:	val_out <= 16'hc4ad;
             14'h23b3 	:	val_out <= 16'hc4b1;
             14'h23b4 	:	val_out <= 16'hc4b5;
             14'h23b5 	:	val_out <= 16'hc4b9;
             14'h23b6 	:	val_out <= 16'hc4bd;
             14'h23b7 	:	val_out <= 16'hc4c1;
             14'h23b8 	:	val_out <= 16'hc4c5;
             14'h23b9 	:	val_out <= 16'hc4c9;
             14'h23ba 	:	val_out <= 16'hc4cd;
             14'h23bb 	:	val_out <= 16'hc4d1;
             14'h23bc 	:	val_out <= 16'hc4d5;
             14'h23bd 	:	val_out <= 16'hc4d9;
             14'h23be 	:	val_out <= 16'hc4dd;
             14'h23bf 	:	val_out <= 16'hc4e1;
             14'h23c0 	:	val_out <= 16'hc4e5;
             14'h23c1 	:	val_out <= 16'hc4e9;
             14'h23c2 	:	val_out <= 16'hc4ed;
             14'h23c3 	:	val_out <= 16'hc4f2;
             14'h23c4 	:	val_out <= 16'hc4f6;
             14'h23c5 	:	val_out <= 16'hc4fa;
             14'h23c6 	:	val_out <= 16'hc4fe;
             14'h23c7 	:	val_out <= 16'hc502;
             14'h23c8 	:	val_out <= 16'hc506;
             14'h23c9 	:	val_out <= 16'hc50a;
             14'h23ca 	:	val_out <= 16'hc50e;
             14'h23cb 	:	val_out <= 16'hc512;
             14'h23cc 	:	val_out <= 16'hc516;
             14'h23cd 	:	val_out <= 16'hc51a;
             14'h23ce 	:	val_out <= 16'hc51e;
             14'h23cf 	:	val_out <= 16'hc522;
             14'h23d0 	:	val_out <= 16'hc526;
             14'h23d1 	:	val_out <= 16'hc52a;
             14'h23d2 	:	val_out <= 16'hc52e;
             14'h23d3 	:	val_out <= 16'hc532;
             14'h23d4 	:	val_out <= 16'hc536;
             14'h23d5 	:	val_out <= 16'hc53a;
             14'h23d6 	:	val_out <= 16'hc53e;
             14'h23d7 	:	val_out <= 16'hc542;
             14'h23d8 	:	val_out <= 16'hc546;
             14'h23d9 	:	val_out <= 16'hc54a;
             14'h23da 	:	val_out <= 16'hc54e;
             14'h23db 	:	val_out <= 16'hc552;
             14'h23dc 	:	val_out <= 16'hc556;
             14'h23dd 	:	val_out <= 16'hc55a;
             14'h23de 	:	val_out <= 16'hc55e;
             14'h23df 	:	val_out <= 16'hc562;
             14'h23e0 	:	val_out <= 16'hc566;
             14'h23e1 	:	val_out <= 16'hc56a;
             14'h23e2 	:	val_out <= 16'hc56e;
             14'h23e3 	:	val_out <= 16'hc572;
             14'h23e4 	:	val_out <= 16'hc576;
             14'h23e5 	:	val_out <= 16'hc57a;
             14'h23e6 	:	val_out <= 16'hc57e;
             14'h23e7 	:	val_out <= 16'hc582;
             14'h23e8 	:	val_out <= 16'hc586;
             14'h23e9 	:	val_out <= 16'hc58a;
             14'h23ea 	:	val_out <= 16'hc58e;
             14'h23eb 	:	val_out <= 16'hc592;
             14'h23ec 	:	val_out <= 16'hc596;
             14'h23ed 	:	val_out <= 16'hc59a;
             14'h23ee 	:	val_out <= 16'hc59e;
             14'h23ef 	:	val_out <= 16'hc5a2;
             14'h23f0 	:	val_out <= 16'hc5a6;
             14'h23f1 	:	val_out <= 16'hc5aa;
             14'h23f2 	:	val_out <= 16'hc5ae;
             14'h23f3 	:	val_out <= 16'hc5b2;
             14'h23f4 	:	val_out <= 16'hc5b6;
             14'h23f5 	:	val_out <= 16'hc5ba;
             14'h23f6 	:	val_out <= 16'hc5be;
             14'h23f7 	:	val_out <= 16'hc5c2;
             14'h23f8 	:	val_out <= 16'hc5c6;
             14'h23f9 	:	val_out <= 16'hc5ca;
             14'h23fa 	:	val_out <= 16'hc5ce;
             14'h23fb 	:	val_out <= 16'hc5d2;
             14'h23fc 	:	val_out <= 16'hc5d6;
             14'h23fd 	:	val_out <= 16'hc5da;
             14'h23fe 	:	val_out <= 16'hc5de;
             14'h23ff 	:	val_out <= 16'hc5e2;
             14'h2400 	:	val_out <= 16'hc5e6;
             14'h2401 	:	val_out <= 16'hc5e9;
             14'h2402 	:	val_out <= 16'hc5ed;
             14'h2403 	:	val_out <= 16'hc5f1;
             14'h2404 	:	val_out <= 16'hc5f5;
             14'h2405 	:	val_out <= 16'hc5f9;
             14'h2406 	:	val_out <= 16'hc5fd;
             14'h2407 	:	val_out <= 16'hc601;
             14'h2408 	:	val_out <= 16'hc605;
             14'h2409 	:	val_out <= 16'hc609;
             14'h240a 	:	val_out <= 16'hc60d;
             14'h240b 	:	val_out <= 16'hc611;
             14'h240c 	:	val_out <= 16'hc615;
             14'h240d 	:	val_out <= 16'hc619;
             14'h240e 	:	val_out <= 16'hc61d;
             14'h240f 	:	val_out <= 16'hc621;
             14'h2410 	:	val_out <= 16'hc625;
             14'h2411 	:	val_out <= 16'hc629;
             14'h2412 	:	val_out <= 16'hc62d;
             14'h2413 	:	val_out <= 16'hc631;
             14'h2414 	:	val_out <= 16'hc635;
             14'h2415 	:	val_out <= 16'hc639;
             14'h2416 	:	val_out <= 16'hc63d;
             14'h2417 	:	val_out <= 16'hc641;
             14'h2418 	:	val_out <= 16'hc645;
             14'h2419 	:	val_out <= 16'hc649;
             14'h241a 	:	val_out <= 16'hc64d;
             14'h241b 	:	val_out <= 16'hc651;
             14'h241c 	:	val_out <= 16'hc655;
             14'h241d 	:	val_out <= 16'hc659;
             14'h241e 	:	val_out <= 16'hc65d;
             14'h241f 	:	val_out <= 16'hc661;
             14'h2420 	:	val_out <= 16'hc665;
             14'h2421 	:	val_out <= 16'hc669;
             14'h2422 	:	val_out <= 16'hc66d;
             14'h2423 	:	val_out <= 16'hc671;
             14'h2424 	:	val_out <= 16'hc675;
             14'h2425 	:	val_out <= 16'hc679;
             14'h2426 	:	val_out <= 16'hc67d;
             14'h2427 	:	val_out <= 16'hc681;
             14'h2428 	:	val_out <= 16'hc685;
             14'h2429 	:	val_out <= 16'hc689;
             14'h242a 	:	val_out <= 16'hc68c;
             14'h242b 	:	val_out <= 16'hc690;
             14'h242c 	:	val_out <= 16'hc694;
             14'h242d 	:	val_out <= 16'hc698;
             14'h242e 	:	val_out <= 16'hc69c;
             14'h242f 	:	val_out <= 16'hc6a0;
             14'h2430 	:	val_out <= 16'hc6a4;
             14'h2431 	:	val_out <= 16'hc6a8;
             14'h2432 	:	val_out <= 16'hc6ac;
             14'h2433 	:	val_out <= 16'hc6b0;
             14'h2434 	:	val_out <= 16'hc6b4;
             14'h2435 	:	val_out <= 16'hc6b8;
             14'h2436 	:	val_out <= 16'hc6bc;
             14'h2437 	:	val_out <= 16'hc6c0;
             14'h2438 	:	val_out <= 16'hc6c4;
             14'h2439 	:	val_out <= 16'hc6c8;
             14'h243a 	:	val_out <= 16'hc6cc;
             14'h243b 	:	val_out <= 16'hc6d0;
             14'h243c 	:	val_out <= 16'hc6d4;
             14'h243d 	:	val_out <= 16'hc6d8;
             14'h243e 	:	val_out <= 16'hc6dc;
             14'h243f 	:	val_out <= 16'hc6e0;
             14'h2440 	:	val_out <= 16'hc6e4;
             14'h2441 	:	val_out <= 16'hc6e8;
             14'h2442 	:	val_out <= 16'hc6ec;
             14'h2443 	:	val_out <= 16'hc6f0;
             14'h2444 	:	val_out <= 16'hc6f3;
             14'h2445 	:	val_out <= 16'hc6f7;
             14'h2446 	:	val_out <= 16'hc6fb;
             14'h2447 	:	val_out <= 16'hc6ff;
             14'h2448 	:	val_out <= 16'hc703;
             14'h2449 	:	val_out <= 16'hc707;
             14'h244a 	:	val_out <= 16'hc70b;
             14'h244b 	:	val_out <= 16'hc70f;
             14'h244c 	:	val_out <= 16'hc713;
             14'h244d 	:	val_out <= 16'hc717;
             14'h244e 	:	val_out <= 16'hc71b;
             14'h244f 	:	val_out <= 16'hc71f;
             14'h2450 	:	val_out <= 16'hc723;
             14'h2451 	:	val_out <= 16'hc727;
             14'h2452 	:	val_out <= 16'hc72b;
             14'h2453 	:	val_out <= 16'hc72f;
             14'h2454 	:	val_out <= 16'hc733;
             14'h2455 	:	val_out <= 16'hc737;
             14'h2456 	:	val_out <= 16'hc73b;
             14'h2457 	:	val_out <= 16'hc73f;
             14'h2458 	:	val_out <= 16'hc742;
             14'h2459 	:	val_out <= 16'hc746;
             14'h245a 	:	val_out <= 16'hc74a;
             14'h245b 	:	val_out <= 16'hc74e;
             14'h245c 	:	val_out <= 16'hc752;
             14'h245d 	:	val_out <= 16'hc756;
             14'h245e 	:	val_out <= 16'hc75a;
             14'h245f 	:	val_out <= 16'hc75e;
             14'h2460 	:	val_out <= 16'hc762;
             14'h2461 	:	val_out <= 16'hc766;
             14'h2462 	:	val_out <= 16'hc76a;
             14'h2463 	:	val_out <= 16'hc76e;
             14'h2464 	:	val_out <= 16'hc772;
             14'h2465 	:	val_out <= 16'hc776;
             14'h2466 	:	val_out <= 16'hc77a;
             14'h2467 	:	val_out <= 16'hc77e;
             14'h2468 	:	val_out <= 16'hc782;
             14'h2469 	:	val_out <= 16'hc785;
             14'h246a 	:	val_out <= 16'hc789;
             14'h246b 	:	val_out <= 16'hc78d;
             14'h246c 	:	val_out <= 16'hc791;
             14'h246d 	:	val_out <= 16'hc795;
             14'h246e 	:	val_out <= 16'hc799;
             14'h246f 	:	val_out <= 16'hc79d;
             14'h2470 	:	val_out <= 16'hc7a1;
             14'h2471 	:	val_out <= 16'hc7a5;
             14'h2472 	:	val_out <= 16'hc7a9;
             14'h2473 	:	val_out <= 16'hc7ad;
             14'h2474 	:	val_out <= 16'hc7b1;
             14'h2475 	:	val_out <= 16'hc7b5;
             14'h2476 	:	val_out <= 16'hc7b9;
             14'h2477 	:	val_out <= 16'hc7bd;
             14'h2478 	:	val_out <= 16'hc7c0;
             14'h2479 	:	val_out <= 16'hc7c4;
             14'h247a 	:	val_out <= 16'hc7c8;
             14'h247b 	:	val_out <= 16'hc7cc;
             14'h247c 	:	val_out <= 16'hc7d0;
             14'h247d 	:	val_out <= 16'hc7d4;
             14'h247e 	:	val_out <= 16'hc7d8;
             14'h247f 	:	val_out <= 16'hc7dc;
             14'h2480 	:	val_out <= 16'hc7e0;
             14'h2481 	:	val_out <= 16'hc7e4;
             14'h2482 	:	val_out <= 16'hc7e8;
             14'h2483 	:	val_out <= 16'hc7ec;
             14'h2484 	:	val_out <= 16'hc7f0;
             14'h2485 	:	val_out <= 16'hc7f3;
             14'h2486 	:	val_out <= 16'hc7f7;
             14'h2487 	:	val_out <= 16'hc7fb;
             14'h2488 	:	val_out <= 16'hc7ff;
             14'h2489 	:	val_out <= 16'hc803;
             14'h248a 	:	val_out <= 16'hc807;
             14'h248b 	:	val_out <= 16'hc80b;
             14'h248c 	:	val_out <= 16'hc80f;
             14'h248d 	:	val_out <= 16'hc813;
             14'h248e 	:	val_out <= 16'hc817;
             14'h248f 	:	val_out <= 16'hc81b;
             14'h2490 	:	val_out <= 16'hc81f;
             14'h2491 	:	val_out <= 16'hc823;
             14'h2492 	:	val_out <= 16'hc826;
             14'h2493 	:	val_out <= 16'hc82a;
             14'h2494 	:	val_out <= 16'hc82e;
             14'h2495 	:	val_out <= 16'hc832;
             14'h2496 	:	val_out <= 16'hc836;
             14'h2497 	:	val_out <= 16'hc83a;
             14'h2498 	:	val_out <= 16'hc83e;
             14'h2499 	:	val_out <= 16'hc842;
             14'h249a 	:	val_out <= 16'hc846;
             14'h249b 	:	val_out <= 16'hc84a;
             14'h249c 	:	val_out <= 16'hc84e;
             14'h249d 	:	val_out <= 16'hc852;
             14'h249e 	:	val_out <= 16'hc855;
             14'h249f 	:	val_out <= 16'hc859;
             14'h24a0 	:	val_out <= 16'hc85d;
             14'h24a1 	:	val_out <= 16'hc861;
             14'h24a2 	:	val_out <= 16'hc865;
             14'h24a3 	:	val_out <= 16'hc869;
             14'h24a4 	:	val_out <= 16'hc86d;
             14'h24a5 	:	val_out <= 16'hc871;
             14'h24a6 	:	val_out <= 16'hc875;
             14'h24a7 	:	val_out <= 16'hc879;
             14'h24a8 	:	val_out <= 16'hc87d;
             14'h24a9 	:	val_out <= 16'hc880;
             14'h24aa 	:	val_out <= 16'hc884;
             14'h24ab 	:	val_out <= 16'hc888;
             14'h24ac 	:	val_out <= 16'hc88c;
             14'h24ad 	:	val_out <= 16'hc890;
             14'h24ae 	:	val_out <= 16'hc894;
             14'h24af 	:	val_out <= 16'hc898;
             14'h24b0 	:	val_out <= 16'hc89c;
             14'h24b1 	:	val_out <= 16'hc8a0;
             14'h24b2 	:	val_out <= 16'hc8a4;
             14'h24b3 	:	val_out <= 16'hc8a7;
             14'h24b4 	:	val_out <= 16'hc8ab;
             14'h24b5 	:	val_out <= 16'hc8af;
             14'h24b6 	:	val_out <= 16'hc8b3;
             14'h24b7 	:	val_out <= 16'hc8b7;
             14'h24b8 	:	val_out <= 16'hc8bb;
             14'h24b9 	:	val_out <= 16'hc8bf;
             14'h24ba 	:	val_out <= 16'hc8c3;
             14'h24bb 	:	val_out <= 16'hc8c7;
             14'h24bc 	:	val_out <= 16'hc8cb;
             14'h24bd 	:	val_out <= 16'hc8ce;
             14'h24be 	:	val_out <= 16'hc8d2;
             14'h24bf 	:	val_out <= 16'hc8d6;
             14'h24c0 	:	val_out <= 16'hc8da;
             14'h24c1 	:	val_out <= 16'hc8de;
             14'h24c2 	:	val_out <= 16'hc8e2;
             14'h24c3 	:	val_out <= 16'hc8e6;
             14'h24c4 	:	val_out <= 16'hc8ea;
             14'h24c5 	:	val_out <= 16'hc8ee;
             14'h24c6 	:	val_out <= 16'hc8f2;
             14'h24c7 	:	val_out <= 16'hc8f5;
             14'h24c8 	:	val_out <= 16'hc8f9;
             14'h24c9 	:	val_out <= 16'hc8fd;
             14'h24ca 	:	val_out <= 16'hc901;
             14'h24cb 	:	val_out <= 16'hc905;
             14'h24cc 	:	val_out <= 16'hc909;
             14'h24cd 	:	val_out <= 16'hc90d;
             14'h24ce 	:	val_out <= 16'hc911;
             14'h24cf 	:	val_out <= 16'hc915;
             14'h24d0 	:	val_out <= 16'hc918;
             14'h24d1 	:	val_out <= 16'hc91c;
             14'h24d2 	:	val_out <= 16'hc920;
             14'h24d3 	:	val_out <= 16'hc924;
             14'h24d4 	:	val_out <= 16'hc928;
             14'h24d5 	:	val_out <= 16'hc92c;
             14'h24d6 	:	val_out <= 16'hc930;
             14'h24d7 	:	val_out <= 16'hc934;
             14'h24d8 	:	val_out <= 16'hc938;
             14'h24d9 	:	val_out <= 16'hc93b;
             14'h24da 	:	val_out <= 16'hc93f;
             14'h24db 	:	val_out <= 16'hc943;
             14'h24dc 	:	val_out <= 16'hc947;
             14'h24dd 	:	val_out <= 16'hc94b;
             14'h24de 	:	val_out <= 16'hc94f;
             14'h24df 	:	val_out <= 16'hc953;
             14'h24e0 	:	val_out <= 16'hc957;
             14'h24e1 	:	val_out <= 16'hc95a;
             14'h24e2 	:	val_out <= 16'hc95e;
             14'h24e3 	:	val_out <= 16'hc962;
             14'h24e4 	:	val_out <= 16'hc966;
             14'h24e5 	:	val_out <= 16'hc96a;
             14'h24e6 	:	val_out <= 16'hc96e;
             14'h24e7 	:	val_out <= 16'hc972;
             14'h24e8 	:	val_out <= 16'hc976;
             14'h24e9 	:	val_out <= 16'hc979;
             14'h24ea 	:	val_out <= 16'hc97d;
             14'h24eb 	:	val_out <= 16'hc981;
             14'h24ec 	:	val_out <= 16'hc985;
             14'h24ed 	:	val_out <= 16'hc989;
             14'h24ee 	:	val_out <= 16'hc98d;
             14'h24ef 	:	val_out <= 16'hc991;
             14'h24f0 	:	val_out <= 16'hc995;
             14'h24f1 	:	val_out <= 16'hc998;
             14'h24f2 	:	val_out <= 16'hc99c;
             14'h24f3 	:	val_out <= 16'hc9a0;
             14'h24f4 	:	val_out <= 16'hc9a4;
             14'h24f5 	:	val_out <= 16'hc9a8;
             14'h24f6 	:	val_out <= 16'hc9ac;
             14'h24f7 	:	val_out <= 16'hc9b0;
             14'h24f8 	:	val_out <= 16'hc9b4;
             14'h24f9 	:	val_out <= 16'hc9b7;
             14'h24fa 	:	val_out <= 16'hc9bb;
             14'h24fb 	:	val_out <= 16'hc9bf;
             14'h24fc 	:	val_out <= 16'hc9c3;
             14'h24fd 	:	val_out <= 16'hc9c7;
             14'h24fe 	:	val_out <= 16'hc9cb;
             14'h24ff 	:	val_out <= 16'hc9cf;
             14'h2500 	:	val_out <= 16'hc9d3;
             14'h2501 	:	val_out <= 16'hc9d6;
             14'h2502 	:	val_out <= 16'hc9da;
             14'h2503 	:	val_out <= 16'hc9de;
             14'h2504 	:	val_out <= 16'hc9e2;
             14'h2505 	:	val_out <= 16'hc9e6;
             14'h2506 	:	val_out <= 16'hc9ea;
             14'h2507 	:	val_out <= 16'hc9ee;
             14'h2508 	:	val_out <= 16'hc9f1;
             14'h2509 	:	val_out <= 16'hc9f5;
             14'h250a 	:	val_out <= 16'hc9f9;
             14'h250b 	:	val_out <= 16'hc9fd;
             14'h250c 	:	val_out <= 16'hca01;
             14'h250d 	:	val_out <= 16'hca05;
             14'h250e 	:	val_out <= 16'hca09;
             14'h250f 	:	val_out <= 16'hca0c;
             14'h2510 	:	val_out <= 16'hca10;
             14'h2511 	:	val_out <= 16'hca14;
             14'h2512 	:	val_out <= 16'hca18;
             14'h2513 	:	val_out <= 16'hca1c;
             14'h2514 	:	val_out <= 16'hca20;
             14'h2515 	:	val_out <= 16'hca24;
             14'h2516 	:	val_out <= 16'hca27;
             14'h2517 	:	val_out <= 16'hca2b;
             14'h2518 	:	val_out <= 16'hca2f;
             14'h2519 	:	val_out <= 16'hca33;
             14'h251a 	:	val_out <= 16'hca37;
             14'h251b 	:	val_out <= 16'hca3b;
             14'h251c 	:	val_out <= 16'hca3f;
             14'h251d 	:	val_out <= 16'hca42;
             14'h251e 	:	val_out <= 16'hca46;
             14'h251f 	:	val_out <= 16'hca4a;
             14'h2520 	:	val_out <= 16'hca4e;
             14'h2521 	:	val_out <= 16'hca52;
             14'h2522 	:	val_out <= 16'hca56;
             14'h2523 	:	val_out <= 16'hca5a;
             14'h2524 	:	val_out <= 16'hca5d;
             14'h2525 	:	val_out <= 16'hca61;
             14'h2526 	:	val_out <= 16'hca65;
             14'h2527 	:	val_out <= 16'hca69;
             14'h2528 	:	val_out <= 16'hca6d;
             14'h2529 	:	val_out <= 16'hca71;
             14'h252a 	:	val_out <= 16'hca74;
             14'h252b 	:	val_out <= 16'hca78;
             14'h252c 	:	val_out <= 16'hca7c;
             14'h252d 	:	val_out <= 16'hca80;
             14'h252e 	:	val_out <= 16'hca84;
             14'h252f 	:	val_out <= 16'hca88;
             14'h2530 	:	val_out <= 16'hca8b;
             14'h2531 	:	val_out <= 16'hca8f;
             14'h2532 	:	val_out <= 16'hca93;
             14'h2533 	:	val_out <= 16'hca97;
             14'h2534 	:	val_out <= 16'hca9b;
             14'h2535 	:	val_out <= 16'hca9f;
             14'h2536 	:	val_out <= 16'hcaa3;
             14'h2537 	:	val_out <= 16'hcaa6;
             14'h2538 	:	val_out <= 16'hcaaa;
             14'h2539 	:	val_out <= 16'hcaae;
             14'h253a 	:	val_out <= 16'hcab2;
             14'h253b 	:	val_out <= 16'hcab6;
             14'h253c 	:	val_out <= 16'hcaba;
             14'h253d 	:	val_out <= 16'hcabd;
             14'h253e 	:	val_out <= 16'hcac1;
             14'h253f 	:	val_out <= 16'hcac5;
             14'h2540 	:	val_out <= 16'hcac9;
             14'h2541 	:	val_out <= 16'hcacd;
             14'h2542 	:	val_out <= 16'hcad1;
             14'h2543 	:	val_out <= 16'hcad4;
             14'h2544 	:	val_out <= 16'hcad8;
             14'h2545 	:	val_out <= 16'hcadc;
             14'h2546 	:	val_out <= 16'hcae0;
             14'h2547 	:	val_out <= 16'hcae4;
             14'h2548 	:	val_out <= 16'hcae8;
             14'h2549 	:	val_out <= 16'hcaeb;
             14'h254a 	:	val_out <= 16'hcaef;
             14'h254b 	:	val_out <= 16'hcaf3;
             14'h254c 	:	val_out <= 16'hcaf7;
             14'h254d 	:	val_out <= 16'hcafb;
             14'h254e 	:	val_out <= 16'hcaff;
             14'h254f 	:	val_out <= 16'hcb02;
             14'h2550 	:	val_out <= 16'hcb06;
             14'h2551 	:	val_out <= 16'hcb0a;
             14'h2552 	:	val_out <= 16'hcb0e;
             14'h2553 	:	val_out <= 16'hcb12;
             14'h2554 	:	val_out <= 16'hcb16;
             14'h2555 	:	val_out <= 16'hcb19;
             14'h2556 	:	val_out <= 16'hcb1d;
             14'h2557 	:	val_out <= 16'hcb21;
             14'h2558 	:	val_out <= 16'hcb25;
             14'h2559 	:	val_out <= 16'hcb29;
             14'h255a 	:	val_out <= 16'hcb2c;
             14'h255b 	:	val_out <= 16'hcb30;
             14'h255c 	:	val_out <= 16'hcb34;
             14'h255d 	:	val_out <= 16'hcb38;
             14'h255e 	:	val_out <= 16'hcb3c;
             14'h255f 	:	val_out <= 16'hcb40;
             14'h2560 	:	val_out <= 16'hcb43;
             14'h2561 	:	val_out <= 16'hcb47;
             14'h2562 	:	val_out <= 16'hcb4b;
             14'h2563 	:	val_out <= 16'hcb4f;
             14'h2564 	:	val_out <= 16'hcb53;
             14'h2565 	:	val_out <= 16'hcb56;
             14'h2566 	:	val_out <= 16'hcb5a;
             14'h2567 	:	val_out <= 16'hcb5e;
             14'h2568 	:	val_out <= 16'hcb62;
             14'h2569 	:	val_out <= 16'hcb66;
             14'h256a 	:	val_out <= 16'hcb6a;
             14'h256b 	:	val_out <= 16'hcb6d;
             14'h256c 	:	val_out <= 16'hcb71;
             14'h256d 	:	val_out <= 16'hcb75;
             14'h256e 	:	val_out <= 16'hcb79;
             14'h256f 	:	val_out <= 16'hcb7d;
             14'h2570 	:	val_out <= 16'hcb80;
             14'h2571 	:	val_out <= 16'hcb84;
             14'h2572 	:	val_out <= 16'hcb88;
             14'h2573 	:	val_out <= 16'hcb8c;
             14'h2574 	:	val_out <= 16'hcb90;
             14'h2575 	:	val_out <= 16'hcb93;
             14'h2576 	:	val_out <= 16'hcb97;
             14'h2577 	:	val_out <= 16'hcb9b;
             14'h2578 	:	val_out <= 16'hcb9f;
             14'h2579 	:	val_out <= 16'hcba3;
             14'h257a 	:	val_out <= 16'hcba7;
             14'h257b 	:	val_out <= 16'hcbaa;
             14'h257c 	:	val_out <= 16'hcbae;
             14'h257d 	:	val_out <= 16'hcbb2;
             14'h257e 	:	val_out <= 16'hcbb6;
             14'h257f 	:	val_out <= 16'hcbba;
             14'h2580 	:	val_out <= 16'hcbbd;
             14'h2581 	:	val_out <= 16'hcbc1;
             14'h2582 	:	val_out <= 16'hcbc5;
             14'h2583 	:	val_out <= 16'hcbc9;
             14'h2584 	:	val_out <= 16'hcbcd;
             14'h2585 	:	val_out <= 16'hcbd0;
             14'h2586 	:	val_out <= 16'hcbd4;
             14'h2587 	:	val_out <= 16'hcbd8;
             14'h2588 	:	val_out <= 16'hcbdc;
             14'h2589 	:	val_out <= 16'hcbe0;
             14'h258a 	:	val_out <= 16'hcbe3;
             14'h258b 	:	val_out <= 16'hcbe7;
             14'h258c 	:	val_out <= 16'hcbeb;
             14'h258d 	:	val_out <= 16'hcbef;
             14'h258e 	:	val_out <= 16'hcbf3;
             14'h258f 	:	val_out <= 16'hcbf6;
             14'h2590 	:	val_out <= 16'hcbfa;
             14'h2591 	:	val_out <= 16'hcbfe;
             14'h2592 	:	val_out <= 16'hcc02;
             14'h2593 	:	val_out <= 16'hcc06;
             14'h2594 	:	val_out <= 16'hcc09;
             14'h2595 	:	val_out <= 16'hcc0d;
             14'h2596 	:	val_out <= 16'hcc11;
             14'h2597 	:	val_out <= 16'hcc15;
             14'h2598 	:	val_out <= 16'hcc19;
             14'h2599 	:	val_out <= 16'hcc1c;
             14'h259a 	:	val_out <= 16'hcc20;
             14'h259b 	:	val_out <= 16'hcc24;
             14'h259c 	:	val_out <= 16'hcc28;
             14'h259d 	:	val_out <= 16'hcc2b;
             14'h259e 	:	val_out <= 16'hcc2f;
             14'h259f 	:	val_out <= 16'hcc33;
             14'h25a0 	:	val_out <= 16'hcc37;
             14'h25a1 	:	val_out <= 16'hcc3b;
             14'h25a2 	:	val_out <= 16'hcc3e;
             14'h25a3 	:	val_out <= 16'hcc42;
             14'h25a4 	:	val_out <= 16'hcc46;
             14'h25a5 	:	val_out <= 16'hcc4a;
             14'h25a6 	:	val_out <= 16'hcc4e;
             14'h25a7 	:	val_out <= 16'hcc51;
             14'h25a8 	:	val_out <= 16'hcc55;
             14'h25a9 	:	val_out <= 16'hcc59;
             14'h25aa 	:	val_out <= 16'hcc5d;
             14'h25ab 	:	val_out <= 16'hcc61;
             14'h25ac 	:	val_out <= 16'hcc64;
             14'h25ad 	:	val_out <= 16'hcc68;
             14'h25ae 	:	val_out <= 16'hcc6c;
             14'h25af 	:	val_out <= 16'hcc70;
             14'h25b0 	:	val_out <= 16'hcc73;
             14'h25b1 	:	val_out <= 16'hcc77;
             14'h25b2 	:	val_out <= 16'hcc7b;
             14'h25b3 	:	val_out <= 16'hcc7f;
             14'h25b4 	:	val_out <= 16'hcc83;
             14'h25b5 	:	val_out <= 16'hcc86;
             14'h25b6 	:	val_out <= 16'hcc8a;
             14'h25b7 	:	val_out <= 16'hcc8e;
             14'h25b8 	:	val_out <= 16'hcc92;
             14'h25b9 	:	val_out <= 16'hcc95;
             14'h25ba 	:	val_out <= 16'hcc99;
             14'h25bb 	:	val_out <= 16'hcc9d;
             14'h25bc 	:	val_out <= 16'hcca1;
             14'h25bd 	:	val_out <= 16'hcca5;
             14'h25be 	:	val_out <= 16'hcca8;
             14'h25bf 	:	val_out <= 16'hccac;
             14'h25c0 	:	val_out <= 16'hccb0;
             14'h25c1 	:	val_out <= 16'hccb4;
             14'h25c2 	:	val_out <= 16'hccb7;
             14'h25c3 	:	val_out <= 16'hccbb;
             14'h25c4 	:	val_out <= 16'hccbf;
             14'h25c5 	:	val_out <= 16'hccc3;
             14'h25c6 	:	val_out <= 16'hccc6;
             14'h25c7 	:	val_out <= 16'hccca;
             14'h25c8 	:	val_out <= 16'hccce;
             14'h25c9 	:	val_out <= 16'hccd2;
             14'h25ca 	:	val_out <= 16'hccd6;
             14'h25cb 	:	val_out <= 16'hccd9;
             14'h25cc 	:	val_out <= 16'hccdd;
             14'h25cd 	:	val_out <= 16'hcce1;
             14'h25ce 	:	val_out <= 16'hcce5;
             14'h25cf 	:	val_out <= 16'hcce8;
             14'h25d0 	:	val_out <= 16'hccec;
             14'h25d1 	:	val_out <= 16'hccf0;
             14'h25d2 	:	val_out <= 16'hccf4;
             14'h25d3 	:	val_out <= 16'hccf7;
             14'h25d4 	:	val_out <= 16'hccfb;
             14'h25d5 	:	val_out <= 16'hccff;
             14'h25d6 	:	val_out <= 16'hcd03;
             14'h25d7 	:	val_out <= 16'hcd07;
             14'h25d8 	:	val_out <= 16'hcd0a;
             14'h25d9 	:	val_out <= 16'hcd0e;
             14'h25da 	:	val_out <= 16'hcd12;
             14'h25db 	:	val_out <= 16'hcd16;
             14'h25dc 	:	val_out <= 16'hcd19;
             14'h25dd 	:	val_out <= 16'hcd1d;
             14'h25de 	:	val_out <= 16'hcd21;
             14'h25df 	:	val_out <= 16'hcd25;
             14'h25e0 	:	val_out <= 16'hcd28;
             14'h25e1 	:	val_out <= 16'hcd2c;
             14'h25e2 	:	val_out <= 16'hcd30;
             14'h25e3 	:	val_out <= 16'hcd34;
             14'h25e4 	:	val_out <= 16'hcd37;
             14'h25e5 	:	val_out <= 16'hcd3b;
             14'h25e6 	:	val_out <= 16'hcd3f;
             14'h25e7 	:	val_out <= 16'hcd43;
             14'h25e8 	:	val_out <= 16'hcd46;
             14'h25e9 	:	val_out <= 16'hcd4a;
             14'h25ea 	:	val_out <= 16'hcd4e;
             14'h25eb 	:	val_out <= 16'hcd52;
             14'h25ec 	:	val_out <= 16'hcd55;
             14'h25ed 	:	val_out <= 16'hcd59;
             14'h25ee 	:	val_out <= 16'hcd5d;
             14'h25ef 	:	val_out <= 16'hcd61;
             14'h25f0 	:	val_out <= 16'hcd64;
             14'h25f1 	:	val_out <= 16'hcd68;
             14'h25f2 	:	val_out <= 16'hcd6c;
             14'h25f3 	:	val_out <= 16'hcd70;
             14'h25f4 	:	val_out <= 16'hcd73;
             14'h25f5 	:	val_out <= 16'hcd77;
             14'h25f6 	:	val_out <= 16'hcd7b;
             14'h25f7 	:	val_out <= 16'hcd7f;
             14'h25f8 	:	val_out <= 16'hcd82;
             14'h25f9 	:	val_out <= 16'hcd86;
             14'h25fa 	:	val_out <= 16'hcd8a;
             14'h25fb 	:	val_out <= 16'hcd8e;
             14'h25fc 	:	val_out <= 16'hcd91;
             14'h25fd 	:	val_out <= 16'hcd95;
             14'h25fe 	:	val_out <= 16'hcd99;
             14'h25ff 	:	val_out <= 16'hcd9d;
             14'h2600 	:	val_out <= 16'hcda0;
             14'h2601 	:	val_out <= 16'hcda4;
             14'h2602 	:	val_out <= 16'hcda8;
             14'h2603 	:	val_out <= 16'hcdac;
             14'h2604 	:	val_out <= 16'hcdaf;
             14'h2605 	:	val_out <= 16'hcdb3;
             14'h2606 	:	val_out <= 16'hcdb7;
             14'h2607 	:	val_out <= 16'hcdbb;
             14'h2608 	:	val_out <= 16'hcdbe;
             14'h2609 	:	val_out <= 16'hcdc2;
             14'h260a 	:	val_out <= 16'hcdc6;
             14'h260b 	:	val_out <= 16'hcdca;
             14'h260c 	:	val_out <= 16'hcdcd;
             14'h260d 	:	val_out <= 16'hcdd1;
             14'h260e 	:	val_out <= 16'hcdd5;
             14'h260f 	:	val_out <= 16'hcdd8;
             14'h2610 	:	val_out <= 16'hcddc;
             14'h2611 	:	val_out <= 16'hcde0;
             14'h2612 	:	val_out <= 16'hcde4;
             14'h2613 	:	val_out <= 16'hcde7;
             14'h2614 	:	val_out <= 16'hcdeb;
             14'h2615 	:	val_out <= 16'hcdef;
             14'h2616 	:	val_out <= 16'hcdf3;
             14'h2617 	:	val_out <= 16'hcdf6;
             14'h2618 	:	val_out <= 16'hcdfa;
             14'h2619 	:	val_out <= 16'hcdfe;
             14'h261a 	:	val_out <= 16'hce02;
             14'h261b 	:	val_out <= 16'hce05;
             14'h261c 	:	val_out <= 16'hce09;
             14'h261d 	:	val_out <= 16'hce0d;
             14'h261e 	:	val_out <= 16'hce10;
             14'h261f 	:	val_out <= 16'hce14;
             14'h2620 	:	val_out <= 16'hce18;
             14'h2621 	:	val_out <= 16'hce1c;
             14'h2622 	:	val_out <= 16'hce1f;
             14'h2623 	:	val_out <= 16'hce23;
             14'h2624 	:	val_out <= 16'hce27;
             14'h2625 	:	val_out <= 16'hce2b;
             14'h2626 	:	val_out <= 16'hce2e;
             14'h2627 	:	val_out <= 16'hce32;
             14'h2628 	:	val_out <= 16'hce36;
             14'h2629 	:	val_out <= 16'hce39;
             14'h262a 	:	val_out <= 16'hce3d;
             14'h262b 	:	val_out <= 16'hce41;
             14'h262c 	:	val_out <= 16'hce45;
             14'h262d 	:	val_out <= 16'hce48;
             14'h262e 	:	val_out <= 16'hce4c;
             14'h262f 	:	val_out <= 16'hce50;
             14'h2630 	:	val_out <= 16'hce53;
             14'h2631 	:	val_out <= 16'hce57;
             14'h2632 	:	val_out <= 16'hce5b;
             14'h2633 	:	val_out <= 16'hce5f;
             14'h2634 	:	val_out <= 16'hce62;
             14'h2635 	:	val_out <= 16'hce66;
             14'h2636 	:	val_out <= 16'hce6a;
             14'h2637 	:	val_out <= 16'hce6d;
             14'h2638 	:	val_out <= 16'hce71;
             14'h2639 	:	val_out <= 16'hce75;
             14'h263a 	:	val_out <= 16'hce79;
             14'h263b 	:	val_out <= 16'hce7c;
             14'h263c 	:	val_out <= 16'hce80;
             14'h263d 	:	val_out <= 16'hce84;
             14'h263e 	:	val_out <= 16'hce87;
             14'h263f 	:	val_out <= 16'hce8b;
             14'h2640 	:	val_out <= 16'hce8f;
             14'h2641 	:	val_out <= 16'hce93;
             14'h2642 	:	val_out <= 16'hce96;
             14'h2643 	:	val_out <= 16'hce9a;
             14'h2644 	:	val_out <= 16'hce9e;
             14'h2645 	:	val_out <= 16'hcea1;
             14'h2646 	:	val_out <= 16'hcea5;
             14'h2647 	:	val_out <= 16'hcea9;
             14'h2648 	:	val_out <= 16'hcead;
             14'h2649 	:	val_out <= 16'hceb0;
             14'h264a 	:	val_out <= 16'hceb4;
             14'h264b 	:	val_out <= 16'hceb8;
             14'h264c 	:	val_out <= 16'hcebb;
             14'h264d 	:	val_out <= 16'hcebf;
             14'h264e 	:	val_out <= 16'hcec3;
             14'h264f 	:	val_out <= 16'hcec7;
             14'h2650 	:	val_out <= 16'hceca;
             14'h2651 	:	val_out <= 16'hcece;
             14'h2652 	:	val_out <= 16'hced2;
             14'h2653 	:	val_out <= 16'hced5;
             14'h2654 	:	val_out <= 16'hced9;
             14'h2655 	:	val_out <= 16'hcedd;
             14'h2656 	:	val_out <= 16'hcee0;
             14'h2657 	:	val_out <= 16'hcee4;
             14'h2658 	:	val_out <= 16'hcee8;
             14'h2659 	:	val_out <= 16'hceec;
             14'h265a 	:	val_out <= 16'hceef;
             14'h265b 	:	val_out <= 16'hcef3;
             14'h265c 	:	val_out <= 16'hcef7;
             14'h265d 	:	val_out <= 16'hcefa;
             14'h265e 	:	val_out <= 16'hcefe;
             14'h265f 	:	val_out <= 16'hcf02;
             14'h2660 	:	val_out <= 16'hcf05;
             14'h2661 	:	val_out <= 16'hcf09;
             14'h2662 	:	val_out <= 16'hcf0d;
             14'h2663 	:	val_out <= 16'hcf11;
             14'h2664 	:	val_out <= 16'hcf14;
             14'h2665 	:	val_out <= 16'hcf18;
             14'h2666 	:	val_out <= 16'hcf1c;
             14'h2667 	:	val_out <= 16'hcf1f;
             14'h2668 	:	val_out <= 16'hcf23;
             14'h2669 	:	val_out <= 16'hcf27;
             14'h266a 	:	val_out <= 16'hcf2a;
             14'h266b 	:	val_out <= 16'hcf2e;
             14'h266c 	:	val_out <= 16'hcf32;
             14'h266d 	:	val_out <= 16'hcf35;
             14'h266e 	:	val_out <= 16'hcf39;
             14'h266f 	:	val_out <= 16'hcf3d;
             14'h2670 	:	val_out <= 16'hcf41;
             14'h2671 	:	val_out <= 16'hcf44;
             14'h2672 	:	val_out <= 16'hcf48;
             14'h2673 	:	val_out <= 16'hcf4c;
             14'h2674 	:	val_out <= 16'hcf4f;
             14'h2675 	:	val_out <= 16'hcf53;
             14'h2676 	:	val_out <= 16'hcf57;
             14'h2677 	:	val_out <= 16'hcf5a;
             14'h2678 	:	val_out <= 16'hcf5e;
             14'h2679 	:	val_out <= 16'hcf62;
             14'h267a 	:	val_out <= 16'hcf65;
             14'h267b 	:	val_out <= 16'hcf69;
             14'h267c 	:	val_out <= 16'hcf6d;
             14'h267d 	:	val_out <= 16'hcf70;
             14'h267e 	:	val_out <= 16'hcf74;
             14'h267f 	:	val_out <= 16'hcf78;
             14'h2680 	:	val_out <= 16'hcf7b;
             14'h2681 	:	val_out <= 16'hcf7f;
             14'h2682 	:	val_out <= 16'hcf83;
             14'h2683 	:	val_out <= 16'hcf87;
             14'h2684 	:	val_out <= 16'hcf8a;
             14'h2685 	:	val_out <= 16'hcf8e;
             14'h2686 	:	val_out <= 16'hcf92;
             14'h2687 	:	val_out <= 16'hcf95;
             14'h2688 	:	val_out <= 16'hcf99;
             14'h2689 	:	val_out <= 16'hcf9d;
             14'h268a 	:	val_out <= 16'hcfa0;
             14'h268b 	:	val_out <= 16'hcfa4;
             14'h268c 	:	val_out <= 16'hcfa8;
             14'h268d 	:	val_out <= 16'hcfab;
             14'h268e 	:	val_out <= 16'hcfaf;
             14'h268f 	:	val_out <= 16'hcfb3;
             14'h2690 	:	val_out <= 16'hcfb6;
             14'h2691 	:	val_out <= 16'hcfba;
             14'h2692 	:	val_out <= 16'hcfbe;
             14'h2693 	:	val_out <= 16'hcfc1;
             14'h2694 	:	val_out <= 16'hcfc5;
             14'h2695 	:	val_out <= 16'hcfc9;
             14'h2696 	:	val_out <= 16'hcfcc;
             14'h2697 	:	val_out <= 16'hcfd0;
             14'h2698 	:	val_out <= 16'hcfd4;
             14'h2699 	:	val_out <= 16'hcfd7;
             14'h269a 	:	val_out <= 16'hcfdb;
             14'h269b 	:	val_out <= 16'hcfdf;
             14'h269c 	:	val_out <= 16'hcfe2;
             14'h269d 	:	val_out <= 16'hcfe6;
             14'h269e 	:	val_out <= 16'hcfea;
             14'h269f 	:	val_out <= 16'hcfed;
             14'h26a0 	:	val_out <= 16'hcff1;
             14'h26a1 	:	val_out <= 16'hcff5;
             14'h26a2 	:	val_out <= 16'hcff8;
             14'h26a3 	:	val_out <= 16'hcffc;
             14'h26a4 	:	val_out <= 16'hd000;
             14'h26a5 	:	val_out <= 16'hd003;
             14'h26a6 	:	val_out <= 16'hd007;
             14'h26a7 	:	val_out <= 16'hd00b;
             14'h26a8 	:	val_out <= 16'hd00e;
             14'h26a9 	:	val_out <= 16'hd012;
             14'h26aa 	:	val_out <= 16'hd016;
             14'h26ab 	:	val_out <= 16'hd019;
             14'h26ac 	:	val_out <= 16'hd01d;
             14'h26ad 	:	val_out <= 16'hd021;
             14'h26ae 	:	val_out <= 16'hd024;
             14'h26af 	:	val_out <= 16'hd028;
             14'h26b0 	:	val_out <= 16'hd02c;
             14'h26b1 	:	val_out <= 16'hd02f;
             14'h26b2 	:	val_out <= 16'hd033;
             14'h26b3 	:	val_out <= 16'hd037;
             14'h26b4 	:	val_out <= 16'hd03a;
             14'h26b5 	:	val_out <= 16'hd03e;
             14'h26b6 	:	val_out <= 16'hd041;
             14'h26b7 	:	val_out <= 16'hd045;
             14'h26b8 	:	val_out <= 16'hd049;
             14'h26b9 	:	val_out <= 16'hd04c;
             14'h26ba 	:	val_out <= 16'hd050;
             14'h26bb 	:	val_out <= 16'hd054;
             14'h26bc 	:	val_out <= 16'hd057;
             14'h26bd 	:	val_out <= 16'hd05b;
             14'h26be 	:	val_out <= 16'hd05f;
             14'h26bf 	:	val_out <= 16'hd062;
             14'h26c0 	:	val_out <= 16'hd066;
             14'h26c1 	:	val_out <= 16'hd06a;
             14'h26c2 	:	val_out <= 16'hd06d;
             14'h26c3 	:	val_out <= 16'hd071;
             14'h26c4 	:	val_out <= 16'hd075;
             14'h26c5 	:	val_out <= 16'hd078;
             14'h26c6 	:	val_out <= 16'hd07c;
             14'h26c7 	:	val_out <= 16'hd080;
             14'h26c8 	:	val_out <= 16'hd083;
             14'h26c9 	:	val_out <= 16'hd087;
             14'h26ca 	:	val_out <= 16'hd08a;
             14'h26cb 	:	val_out <= 16'hd08e;
             14'h26cc 	:	val_out <= 16'hd092;
             14'h26cd 	:	val_out <= 16'hd095;
             14'h26ce 	:	val_out <= 16'hd099;
             14'h26cf 	:	val_out <= 16'hd09d;
             14'h26d0 	:	val_out <= 16'hd0a0;
             14'h26d1 	:	val_out <= 16'hd0a4;
             14'h26d2 	:	val_out <= 16'hd0a8;
             14'h26d3 	:	val_out <= 16'hd0ab;
             14'h26d4 	:	val_out <= 16'hd0af;
             14'h26d5 	:	val_out <= 16'hd0b3;
             14'h26d6 	:	val_out <= 16'hd0b6;
             14'h26d7 	:	val_out <= 16'hd0ba;
             14'h26d8 	:	val_out <= 16'hd0bd;
             14'h26d9 	:	val_out <= 16'hd0c1;
             14'h26da 	:	val_out <= 16'hd0c5;
             14'h26db 	:	val_out <= 16'hd0c8;
             14'h26dc 	:	val_out <= 16'hd0cc;
             14'h26dd 	:	val_out <= 16'hd0d0;
             14'h26de 	:	val_out <= 16'hd0d3;
             14'h26df 	:	val_out <= 16'hd0d7;
             14'h26e0 	:	val_out <= 16'hd0db;
             14'h26e1 	:	val_out <= 16'hd0de;
             14'h26e2 	:	val_out <= 16'hd0e2;
             14'h26e3 	:	val_out <= 16'hd0e5;
             14'h26e4 	:	val_out <= 16'hd0e9;
             14'h26e5 	:	val_out <= 16'hd0ed;
             14'h26e6 	:	val_out <= 16'hd0f0;
             14'h26e7 	:	val_out <= 16'hd0f4;
             14'h26e8 	:	val_out <= 16'hd0f8;
             14'h26e9 	:	val_out <= 16'hd0fb;
             14'h26ea 	:	val_out <= 16'hd0ff;
             14'h26eb 	:	val_out <= 16'hd102;
             14'h26ec 	:	val_out <= 16'hd106;
             14'h26ed 	:	val_out <= 16'hd10a;
             14'h26ee 	:	val_out <= 16'hd10d;
             14'h26ef 	:	val_out <= 16'hd111;
             14'h26f0 	:	val_out <= 16'hd115;
             14'h26f1 	:	val_out <= 16'hd118;
             14'h26f2 	:	val_out <= 16'hd11c;
             14'h26f3 	:	val_out <= 16'hd11f;
             14'h26f4 	:	val_out <= 16'hd123;
             14'h26f5 	:	val_out <= 16'hd127;
             14'h26f6 	:	val_out <= 16'hd12a;
             14'h26f7 	:	val_out <= 16'hd12e;
             14'h26f8 	:	val_out <= 16'hd132;
             14'h26f9 	:	val_out <= 16'hd135;
             14'h26fa 	:	val_out <= 16'hd139;
             14'h26fb 	:	val_out <= 16'hd13c;
             14'h26fc 	:	val_out <= 16'hd140;
             14'h26fd 	:	val_out <= 16'hd144;
             14'h26fe 	:	val_out <= 16'hd147;
             14'h26ff 	:	val_out <= 16'hd14b;
             14'h2700 	:	val_out <= 16'hd14f;
             14'h2701 	:	val_out <= 16'hd152;
             14'h2702 	:	val_out <= 16'hd156;
             14'h2703 	:	val_out <= 16'hd159;
             14'h2704 	:	val_out <= 16'hd15d;
             14'h2705 	:	val_out <= 16'hd161;
             14'h2706 	:	val_out <= 16'hd164;
             14'h2707 	:	val_out <= 16'hd168;
             14'h2708 	:	val_out <= 16'hd16b;
             14'h2709 	:	val_out <= 16'hd16f;
             14'h270a 	:	val_out <= 16'hd173;
             14'h270b 	:	val_out <= 16'hd176;
             14'h270c 	:	val_out <= 16'hd17a;
             14'h270d 	:	val_out <= 16'hd17e;
             14'h270e 	:	val_out <= 16'hd181;
             14'h270f 	:	val_out <= 16'hd185;
             14'h2710 	:	val_out <= 16'hd188;
             14'h2711 	:	val_out <= 16'hd18c;
             14'h2712 	:	val_out <= 16'hd190;
             14'h2713 	:	val_out <= 16'hd193;
             14'h2714 	:	val_out <= 16'hd197;
             14'h2715 	:	val_out <= 16'hd19a;
             14'h2716 	:	val_out <= 16'hd19e;
             14'h2717 	:	val_out <= 16'hd1a2;
             14'h2718 	:	val_out <= 16'hd1a5;
             14'h2719 	:	val_out <= 16'hd1a9;
             14'h271a 	:	val_out <= 16'hd1ac;
             14'h271b 	:	val_out <= 16'hd1b0;
             14'h271c 	:	val_out <= 16'hd1b4;
             14'h271d 	:	val_out <= 16'hd1b7;
             14'h271e 	:	val_out <= 16'hd1bb;
             14'h271f 	:	val_out <= 16'hd1be;
             14'h2720 	:	val_out <= 16'hd1c2;
             14'h2721 	:	val_out <= 16'hd1c6;
             14'h2722 	:	val_out <= 16'hd1c9;
             14'h2723 	:	val_out <= 16'hd1cd;
             14'h2724 	:	val_out <= 16'hd1d0;
             14'h2725 	:	val_out <= 16'hd1d4;
             14'h2726 	:	val_out <= 16'hd1d8;
             14'h2727 	:	val_out <= 16'hd1db;
             14'h2728 	:	val_out <= 16'hd1df;
             14'h2729 	:	val_out <= 16'hd1e2;
             14'h272a 	:	val_out <= 16'hd1e6;
             14'h272b 	:	val_out <= 16'hd1ea;
             14'h272c 	:	val_out <= 16'hd1ed;
             14'h272d 	:	val_out <= 16'hd1f1;
             14'h272e 	:	val_out <= 16'hd1f4;
             14'h272f 	:	val_out <= 16'hd1f8;
             14'h2730 	:	val_out <= 16'hd1fc;
             14'h2731 	:	val_out <= 16'hd1ff;
             14'h2732 	:	val_out <= 16'hd203;
             14'h2733 	:	val_out <= 16'hd206;
             14'h2734 	:	val_out <= 16'hd20a;
             14'h2735 	:	val_out <= 16'hd20e;
             14'h2736 	:	val_out <= 16'hd211;
             14'h2737 	:	val_out <= 16'hd215;
             14'h2738 	:	val_out <= 16'hd218;
             14'h2739 	:	val_out <= 16'hd21c;
             14'h273a 	:	val_out <= 16'hd220;
             14'h273b 	:	val_out <= 16'hd223;
             14'h273c 	:	val_out <= 16'hd227;
             14'h273d 	:	val_out <= 16'hd22a;
             14'h273e 	:	val_out <= 16'hd22e;
             14'h273f 	:	val_out <= 16'hd231;
             14'h2740 	:	val_out <= 16'hd235;
             14'h2741 	:	val_out <= 16'hd239;
             14'h2742 	:	val_out <= 16'hd23c;
             14'h2743 	:	val_out <= 16'hd240;
             14'h2744 	:	val_out <= 16'hd243;
             14'h2745 	:	val_out <= 16'hd247;
             14'h2746 	:	val_out <= 16'hd24b;
             14'h2747 	:	val_out <= 16'hd24e;
             14'h2748 	:	val_out <= 16'hd252;
             14'h2749 	:	val_out <= 16'hd255;
             14'h274a 	:	val_out <= 16'hd259;
             14'h274b 	:	val_out <= 16'hd25c;
             14'h274c 	:	val_out <= 16'hd260;
             14'h274d 	:	val_out <= 16'hd264;
             14'h274e 	:	val_out <= 16'hd267;
             14'h274f 	:	val_out <= 16'hd26b;
             14'h2750 	:	val_out <= 16'hd26e;
             14'h2751 	:	val_out <= 16'hd272;
             14'h2752 	:	val_out <= 16'hd276;
             14'h2753 	:	val_out <= 16'hd279;
             14'h2754 	:	val_out <= 16'hd27d;
             14'h2755 	:	val_out <= 16'hd280;
             14'h2756 	:	val_out <= 16'hd284;
             14'h2757 	:	val_out <= 16'hd287;
             14'h2758 	:	val_out <= 16'hd28b;
             14'h2759 	:	val_out <= 16'hd28f;
             14'h275a 	:	val_out <= 16'hd292;
             14'h275b 	:	val_out <= 16'hd296;
             14'h275c 	:	val_out <= 16'hd299;
             14'h275d 	:	val_out <= 16'hd29d;
             14'h275e 	:	val_out <= 16'hd2a0;
             14'h275f 	:	val_out <= 16'hd2a4;
             14'h2760 	:	val_out <= 16'hd2a8;
             14'h2761 	:	val_out <= 16'hd2ab;
             14'h2762 	:	val_out <= 16'hd2af;
             14'h2763 	:	val_out <= 16'hd2b2;
             14'h2764 	:	val_out <= 16'hd2b6;
             14'h2765 	:	val_out <= 16'hd2b9;
             14'h2766 	:	val_out <= 16'hd2bd;
             14'h2767 	:	val_out <= 16'hd2c1;
             14'h2768 	:	val_out <= 16'hd2c4;
             14'h2769 	:	val_out <= 16'hd2c8;
             14'h276a 	:	val_out <= 16'hd2cb;
             14'h276b 	:	val_out <= 16'hd2cf;
             14'h276c 	:	val_out <= 16'hd2d2;
             14'h276d 	:	val_out <= 16'hd2d6;
             14'h276e 	:	val_out <= 16'hd2da;
             14'h276f 	:	val_out <= 16'hd2dd;
             14'h2770 	:	val_out <= 16'hd2e1;
             14'h2771 	:	val_out <= 16'hd2e4;
             14'h2772 	:	val_out <= 16'hd2e8;
             14'h2773 	:	val_out <= 16'hd2eb;
             14'h2774 	:	val_out <= 16'hd2ef;
             14'h2775 	:	val_out <= 16'hd2f2;
             14'h2776 	:	val_out <= 16'hd2f6;
             14'h2777 	:	val_out <= 16'hd2fa;
             14'h2778 	:	val_out <= 16'hd2fd;
             14'h2779 	:	val_out <= 16'hd301;
             14'h277a 	:	val_out <= 16'hd304;
             14'h277b 	:	val_out <= 16'hd308;
             14'h277c 	:	val_out <= 16'hd30b;
             14'h277d 	:	val_out <= 16'hd30f;
             14'h277e 	:	val_out <= 16'hd312;
             14'h277f 	:	val_out <= 16'hd316;
             14'h2780 	:	val_out <= 16'hd31a;
             14'h2781 	:	val_out <= 16'hd31d;
             14'h2782 	:	val_out <= 16'hd321;
             14'h2783 	:	val_out <= 16'hd324;
             14'h2784 	:	val_out <= 16'hd328;
             14'h2785 	:	val_out <= 16'hd32b;
             14'h2786 	:	val_out <= 16'hd32f;
             14'h2787 	:	val_out <= 16'hd332;
             14'h2788 	:	val_out <= 16'hd336;
             14'h2789 	:	val_out <= 16'hd33a;
             14'h278a 	:	val_out <= 16'hd33d;
             14'h278b 	:	val_out <= 16'hd341;
             14'h278c 	:	val_out <= 16'hd344;
             14'h278d 	:	val_out <= 16'hd348;
             14'h278e 	:	val_out <= 16'hd34b;
             14'h278f 	:	val_out <= 16'hd34f;
             14'h2790 	:	val_out <= 16'hd352;
             14'h2791 	:	val_out <= 16'hd356;
             14'h2792 	:	val_out <= 16'hd359;
             14'h2793 	:	val_out <= 16'hd35d;
             14'h2794 	:	val_out <= 16'hd361;
             14'h2795 	:	val_out <= 16'hd364;
             14'h2796 	:	val_out <= 16'hd368;
             14'h2797 	:	val_out <= 16'hd36b;
             14'h2798 	:	val_out <= 16'hd36f;
             14'h2799 	:	val_out <= 16'hd372;
             14'h279a 	:	val_out <= 16'hd376;
             14'h279b 	:	val_out <= 16'hd379;
             14'h279c 	:	val_out <= 16'hd37d;
             14'h279d 	:	val_out <= 16'hd380;
             14'h279e 	:	val_out <= 16'hd384;
             14'h279f 	:	val_out <= 16'hd388;
             14'h27a0 	:	val_out <= 16'hd38b;
             14'h27a1 	:	val_out <= 16'hd38f;
             14'h27a2 	:	val_out <= 16'hd392;
             14'h27a3 	:	val_out <= 16'hd396;
             14'h27a4 	:	val_out <= 16'hd399;
             14'h27a5 	:	val_out <= 16'hd39d;
             14'h27a6 	:	val_out <= 16'hd3a0;
             14'h27a7 	:	val_out <= 16'hd3a4;
             14'h27a8 	:	val_out <= 16'hd3a7;
             14'h27a9 	:	val_out <= 16'hd3ab;
             14'h27aa 	:	val_out <= 16'hd3ae;
             14'h27ab 	:	val_out <= 16'hd3b2;
             14'h27ac 	:	val_out <= 16'hd3b5;
             14'h27ad 	:	val_out <= 16'hd3b9;
             14'h27ae 	:	val_out <= 16'hd3bd;
             14'h27af 	:	val_out <= 16'hd3c0;
             14'h27b0 	:	val_out <= 16'hd3c4;
             14'h27b1 	:	val_out <= 16'hd3c7;
             14'h27b2 	:	val_out <= 16'hd3cb;
             14'h27b3 	:	val_out <= 16'hd3ce;
             14'h27b4 	:	val_out <= 16'hd3d2;
             14'h27b5 	:	val_out <= 16'hd3d5;
             14'h27b6 	:	val_out <= 16'hd3d9;
             14'h27b7 	:	val_out <= 16'hd3dc;
             14'h27b8 	:	val_out <= 16'hd3e0;
             14'h27b9 	:	val_out <= 16'hd3e3;
             14'h27ba 	:	val_out <= 16'hd3e7;
             14'h27bb 	:	val_out <= 16'hd3ea;
             14'h27bc 	:	val_out <= 16'hd3ee;
             14'h27bd 	:	val_out <= 16'hd3f1;
             14'h27be 	:	val_out <= 16'hd3f5;
             14'h27bf 	:	val_out <= 16'hd3f8;
             14'h27c0 	:	val_out <= 16'hd3fc;
             14'h27c1 	:	val_out <= 16'hd400;
             14'h27c2 	:	val_out <= 16'hd403;
             14'h27c3 	:	val_out <= 16'hd407;
             14'h27c4 	:	val_out <= 16'hd40a;
             14'h27c5 	:	val_out <= 16'hd40e;
             14'h27c6 	:	val_out <= 16'hd411;
             14'h27c7 	:	val_out <= 16'hd415;
             14'h27c8 	:	val_out <= 16'hd418;
             14'h27c9 	:	val_out <= 16'hd41c;
             14'h27ca 	:	val_out <= 16'hd41f;
             14'h27cb 	:	val_out <= 16'hd423;
             14'h27cc 	:	val_out <= 16'hd426;
             14'h27cd 	:	val_out <= 16'hd42a;
             14'h27ce 	:	val_out <= 16'hd42d;
             14'h27cf 	:	val_out <= 16'hd431;
             14'h27d0 	:	val_out <= 16'hd434;
             14'h27d1 	:	val_out <= 16'hd438;
             14'h27d2 	:	val_out <= 16'hd43b;
             14'h27d3 	:	val_out <= 16'hd43f;
             14'h27d4 	:	val_out <= 16'hd442;
             14'h27d5 	:	val_out <= 16'hd446;
             14'h27d6 	:	val_out <= 16'hd449;
             14'h27d7 	:	val_out <= 16'hd44d;
             14'h27d8 	:	val_out <= 16'hd450;
             14'h27d9 	:	val_out <= 16'hd454;
             14'h27da 	:	val_out <= 16'hd457;
             14'h27db 	:	val_out <= 16'hd45b;
             14'h27dc 	:	val_out <= 16'hd45e;
             14'h27dd 	:	val_out <= 16'hd462;
             14'h27de 	:	val_out <= 16'hd465;
             14'h27df 	:	val_out <= 16'hd469;
             14'h27e0 	:	val_out <= 16'hd46c;
             14'h27e1 	:	val_out <= 16'hd470;
             14'h27e2 	:	val_out <= 16'hd473;
             14'h27e3 	:	val_out <= 16'hd477;
             14'h27e4 	:	val_out <= 16'hd47b;
             14'h27e5 	:	val_out <= 16'hd47e;
             14'h27e6 	:	val_out <= 16'hd482;
             14'h27e7 	:	val_out <= 16'hd485;
             14'h27e8 	:	val_out <= 16'hd489;
             14'h27e9 	:	val_out <= 16'hd48c;
             14'h27ea 	:	val_out <= 16'hd490;
             14'h27eb 	:	val_out <= 16'hd493;
             14'h27ec 	:	val_out <= 16'hd497;
             14'h27ed 	:	val_out <= 16'hd49a;
             14'h27ee 	:	val_out <= 16'hd49e;
             14'h27ef 	:	val_out <= 16'hd4a1;
             14'h27f0 	:	val_out <= 16'hd4a5;
             14'h27f1 	:	val_out <= 16'hd4a8;
             14'h27f2 	:	val_out <= 16'hd4ac;
             14'h27f3 	:	val_out <= 16'hd4af;
             14'h27f4 	:	val_out <= 16'hd4b3;
             14'h27f5 	:	val_out <= 16'hd4b6;
             14'h27f6 	:	val_out <= 16'hd4ba;
             14'h27f7 	:	val_out <= 16'hd4bd;
             14'h27f8 	:	val_out <= 16'hd4c0;
             14'h27f9 	:	val_out <= 16'hd4c4;
             14'h27fa 	:	val_out <= 16'hd4c7;
             14'h27fb 	:	val_out <= 16'hd4cb;
             14'h27fc 	:	val_out <= 16'hd4ce;
             14'h27fd 	:	val_out <= 16'hd4d2;
             14'h27fe 	:	val_out <= 16'hd4d5;
             14'h27ff 	:	val_out <= 16'hd4d9;
             14'h2800 	:	val_out <= 16'hd4dc;
             14'h2801 	:	val_out <= 16'hd4e0;
             14'h2802 	:	val_out <= 16'hd4e3;
             14'h2803 	:	val_out <= 16'hd4e7;
             14'h2804 	:	val_out <= 16'hd4ea;
             14'h2805 	:	val_out <= 16'hd4ee;
             14'h2806 	:	val_out <= 16'hd4f1;
             14'h2807 	:	val_out <= 16'hd4f5;
             14'h2808 	:	val_out <= 16'hd4f8;
             14'h2809 	:	val_out <= 16'hd4fc;
             14'h280a 	:	val_out <= 16'hd4ff;
             14'h280b 	:	val_out <= 16'hd503;
             14'h280c 	:	val_out <= 16'hd506;
             14'h280d 	:	val_out <= 16'hd50a;
             14'h280e 	:	val_out <= 16'hd50d;
             14'h280f 	:	val_out <= 16'hd511;
             14'h2810 	:	val_out <= 16'hd514;
             14'h2811 	:	val_out <= 16'hd518;
             14'h2812 	:	val_out <= 16'hd51b;
             14'h2813 	:	val_out <= 16'hd51f;
             14'h2814 	:	val_out <= 16'hd522;
             14'h2815 	:	val_out <= 16'hd526;
             14'h2816 	:	val_out <= 16'hd529;
             14'h2817 	:	val_out <= 16'hd52d;
             14'h2818 	:	val_out <= 16'hd530;
             14'h2819 	:	val_out <= 16'hd534;
             14'h281a 	:	val_out <= 16'hd537;
             14'h281b 	:	val_out <= 16'hd53a;
             14'h281c 	:	val_out <= 16'hd53e;
             14'h281d 	:	val_out <= 16'hd541;
             14'h281e 	:	val_out <= 16'hd545;
             14'h281f 	:	val_out <= 16'hd548;
             14'h2820 	:	val_out <= 16'hd54c;
             14'h2821 	:	val_out <= 16'hd54f;
             14'h2822 	:	val_out <= 16'hd553;
             14'h2823 	:	val_out <= 16'hd556;
             14'h2824 	:	val_out <= 16'hd55a;
             14'h2825 	:	val_out <= 16'hd55d;
             14'h2826 	:	val_out <= 16'hd561;
             14'h2827 	:	val_out <= 16'hd564;
             14'h2828 	:	val_out <= 16'hd568;
             14'h2829 	:	val_out <= 16'hd56b;
             14'h282a 	:	val_out <= 16'hd56f;
             14'h282b 	:	val_out <= 16'hd572;
             14'h282c 	:	val_out <= 16'hd576;
             14'h282d 	:	val_out <= 16'hd579;
             14'h282e 	:	val_out <= 16'hd57c;
             14'h282f 	:	val_out <= 16'hd580;
             14'h2830 	:	val_out <= 16'hd583;
             14'h2831 	:	val_out <= 16'hd587;
             14'h2832 	:	val_out <= 16'hd58a;
             14'h2833 	:	val_out <= 16'hd58e;
             14'h2834 	:	val_out <= 16'hd591;
             14'h2835 	:	val_out <= 16'hd595;
             14'h2836 	:	val_out <= 16'hd598;
             14'h2837 	:	val_out <= 16'hd59c;
             14'h2838 	:	val_out <= 16'hd59f;
             14'h2839 	:	val_out <= 16'hd5a3;
             14'h283a 	:	val_out <= 16'hd5a6;
             14'h283b 	:	val_out <= 16'hd5aa;
             14'h283c 	:	val_out <= 16'hd5ad;
             14'h283d 	:	val_out <= 16'hd5b0;
             14'h283e 	:	val_out <= 16'hd5b4;
             14'h283f 	:	val_out <= 16'hd5b7;
             14'h2840 	:	val_out <= 16'hd5bb;
             14'h2841 	:	val_out <= 16'hd5be;
             14'h2842 	:	val_out <= 16'hd5c2;
             14'h2843 	:	val_out <= 16'hd5c5;
             14'h2844 	:	val_out <= 16'hd5c9;
             14'h2845 	:	val_out <= 16'hd5cc;
             14'h2846 	:	val_out <= 16'hd5d0;
             14'h2847 	:	val_out <= 16'hd5d3;
             14'h2848 	:	val_out <= 16'hd5d6;
             14'h2849 	:	val_out <= 16'hd5da;
             14'h284a 	:	val_out <= 16'hd5dd;
             14'h284b 	:	val_out <= 16'hd5e1;
             14'h284c 	:	val_out <= 16'hd5e4;
             14'h284d 	:	val_out <= 16'hd5e8;
             14'h284e 	:	val_out <= 16'hd5eb;
             14'h284f 	:	val_out <= 16'hd5ef;
             14'h2850 	:	val_out <= 16'hd5f2;
             14'h2851 	:	val_out <= 16'hd5f6;
             14'h2852 	:	val_out <= 16'hd5f9;
             14'h2853 	:	val_out <= 16'hd5fc;
             14'h2854 	:	val_out <= 16'hd600;
             14'h2855 	:	val_out <= 16'hd603;
             14'h2856 	:	val_out <= 16'hd607;
             14'h2857 	:	val_out <= 16'hd60a;
             14'h2858 	:	val_out <= 16'hd60e;
             14'h2859 	:	val_out <= 16'hd611;
             14'h285a 	:	val_out <= 16'hd615;
             14'h285b 	:	val_out <= 16'hd618;
             14'h285c 	:	val_out <= 16'hd61b;
             14'h285d 	:	val_out <= 16'hd61f;
             14'h285e 	:	val_out <= 16'hd622;
             14'h285f 	:	val_out <= 16'hd626;
             14'h2860 	:	val_out <= 16'hd629;
             14'h2861 	:	val_out <= 16'hd62d;
             14'h2862 	:	val_out <= 16'hd630;
             14'h2863 	:	val_out <= 16'hd634;
             14'h2864 	:	val_out <= 16'hd637;
             14'h2865 	:	val_out <= 16'hd63a;
             14'h2866 	:	val_out <= 16'hd63e;
             14'h2867 	:	val_out <= 16'hd641;
             14'h2868 	:	val_out <= 16'hd645;
             14'h2869 	:	val_out <= 16'hd648;
             14'h286a 	:	val_out <= 16'hd64c;
             14'h286b 	:	val_out <= 16'hd64f;
             14'h286c 	:	val_out <= 16'hd652;
             14'h286d 	:	val_out <= 16'hd656;
             14'h286e 	:	val_out <= 16'hd659;
             14'h286f 	:	val_out <= 16'hd65d;
             14'h2870 	:	val_out <= 16'hd660;
             14'h2871 	:	val_out <= 16'hd664;
             14'h2872 	:	val_out <= 16'hd667;
             14'h2873 	:	val_out <= 16'hd66b;
             14'h2874 	:	val_out <= 16'hd66e;
             14'h2875 	:	val_out <= 16'hd671;
             14'h2876 	:	val_out <= 16'hd675;
             14'h2877 	:	val_out <= 16'hd678;
             14'h2878 	:	val_out <= 16'hd67c;
             14'h2879 	:	val_out <= 16'hd67f;
             14'h287a 	:	val_out <= 16'hd683;
             14'h287b 	:	val_out <= 16'hd686;
             14'h287c 	:	val_out <= 16'hd689;
             14'h287d 	:	val_out <= 16'hd68d;
             14'h287e 	:	val_out <= 16'hd690;
             14'h287f 	:	val_out <= 16'hd694;
             14'h2880 	:	val_out <= 16'hd697;
             14'h2881 	:	val_out <= 16'hd69b;
             14'h2882 	:	val_out <= 16'hd69e;
             14'h2883 	:	val_out <= 16'hd6a1;
             14'h2884 	:	val_out <= 16'hd6a5;
             14'h2885 	:	val_out <= 16'hd6a8;
             14'h2886 	:	val_out <= 16'hd6ac;
             14'h2887 	:	val_out <= 16'hd6af;
             14'h2888 	:	val_out <= 16'hd6b3;
             14'h2889 	:	val_out <= 16'hd6b6;
             14'h288a 	:	val_out <= 16'hd6b9;
             14'h288b 	:	val_out <= 16'hd6bd;
             14'h288c 	:	val_out <= 16'hd6c0;
             14'h288d 	:	val_out <= 16'hd6c4;
             14'h288e 	:	val_out <= 16'hd6c7;
             14'h288f 	:	val_out <= 16'hd6ca;
             14'h2890 	:	val_out <= 16'hd6ce;
             14'h2891 	:	val_out <= 16'hd6d1;
             14'h2892 	:	val_out <= 16'hd6d5;
             14'h2893 	:	val_out <= 16'hd6d8;
             14'h2894 	:	val_out <= 16'hd6dc;
             14'h2895 	:	val_out <= 16'hd6df;
             14'h2896 	:	val_out <= 16'hd6e2;
             14'h2897 	:	val_out <= 16'hd6e6;
             14'h2898 	:	val_out <= 16'hd6e9;
             14'h2899 	:	val_out <= 16'hd6ed;
             14'h289a 	:	val_out <= 16'hd6f0;
             14'h289b 	:	val_out <= 16'hd6f3;
             14'h289c 	:	val_out <= 16'hd6f7;
             14'h289d 	:	val_out <= 16'hd6fa;
             14'h289e 	:	val_out <= 16'hd6fe;
             14'h289f 	:	val_out <= 16'hd701;
             14'h28a0 	:	val_out <= 16'hd704;
             14'h28a1 	:	val_out <= 16'hd708;
             14'h28a2 	:	val_out <= 16'hd70b;
             14'h28a3 	:	val_out <= 16'hd70f;
             14'h28a4 	:	val_out <= 16'hd712;
             14'h28a5 	:	val_out <= 16'hd716;
             14'h28a6 	:	val_out <= 16'hd719;
             14'h28a7 	:	val_out <= 16'hd71c;
             14'h28a8 	:	val_out <= 16'hd720;
             14'h28a9 	:	val_out <= 16'hd723;
             14'h28aa 	:	val_out <= 16'hd727;
             14'h28ab 	:	val_out <= 16'hd72a;
             14'h28ac 	:	val_out <= 16'hd72d;
             14'h28ad 	:	val_out <= 16'hd731;
             14'h28ae 	:	val_out <= 16'hd734;
             14'h28af 	:	val_out <= 16'hd738;
             14'h28b0 	:	val_out <= 16'hd73b;
             14'h28b1 	:	val_out <= 16'hd73e;
             14'h28b2 	:	val_out <= 16'hd742;
             14'h28b3 	:	val_out <= 16'hd745;
             14'h28b4 	:	val_out <= 16'hd749;
             14'h28b5 	:	val_out <= 16'hd74c;
             14'h28b6 	:	val_out <= 16'hd74f;
             14'h28b7 	:	val_out <= 16'hd753;
             14'h28b8 	:	val_out <= 16'hd756;
             14'h28b9 	:	val_out <= 16'hd75a;
             14'h28ba 	:	val_out <= 16'hd75d;
             14'h28bb 	:	val_out <= 16'hd760;
             14'h28bc 	:	val_out <= 16'hd764;
             14'h28bd 	:	val_out <= 16'hd767;
             14'h28be 	:	val_out <= 16'hd76b;
             14'h28bf 	:	val_out <= 16'hd76e;
             14'h28c0 	:	val_out <= 16'hd771;
             14'h28c1 	:	val_out <= 16'hd775;
             14'h28c2 	:	val_out <= 16'hd778;
             14'h28c3 	:	val_out <= 16'hd77c;
             14'h28c4 	:	val_out <= 16'hd77f;
             14'h28c5 	:	val_out <= 16'hd782;
             14'h28c6 	:	val_out <= 16'hd786;
             14'h28c7 	:	val_out <= 16'hd789;
             14'h28c8 	:	val_out <= 16'hd78c;
             14'h28c9 	:	val_out <= 16'hd790;
             14'h28ca 	:	val_out <= 16'hd793;
             14'h28cb 	:	val_out <= 16'hd797;
             14'h28cc 	:	val_out <= 16'hd79a;
             14'h28cd 	:	val_out <= 16'hd79d;
             14'h28ce 	:	val_out <= 16'hd7a1;
             14'h28cf 	:	val_out <= 16'hd7a4;
             14'h28d0 	:	val_out <= 16'hd7a8;
             14'h28d1 	:	val_out <= 16'hd7ab;
             14'h28d2 	:	val_out <= 16'hd7ae;
             14'h28d3 	:	val_out <= 16'hd7b2;
             14'h28d4 	:	val_out <= 16'hd7b5;
             14'h28d5 	:	val_out <= 16'hd7b9;
             14'h28d6 	:	val_out <= 16'hd7bc;
             14'h28d7 	:	val_out <= 16'hd7bf;
             14'h28d8 	:	val_out <= 16'hd7c3;
             14'h28d9 	:	val_out <= 16'hd7c6;
             14'h28da 	:	val_out <= 16'hd7c9;
             14'h28db 	:	val_out <= 16'hd7cd;
             14'h28dc 	:	val_out <= 16'hd7d0;
             14'h28dd 	:	val_out <= 16'hd7d4;
             14'h28de 	:	val_out <= 16'hd7d7;
             14'h28df 	:	val_out <= 16'hd7da;
             14'h28e0 	:	val_out <= 16'hd7de;
             14'h28e1 	:	val_out <= 16'hd7e1;
             14'h28e2 	:	val_out <= 16'hd7e4;
             14'h28e3 	:	val_out <= 16'hd7e8;
             14'h28e4 	:	val_out <= 16'hd7eb;
             14'h28e5 	:	val_out <= 16'hd7ef;
             14'h28e6 	:	val_out <= 16'hd7f2;
             14'h28e7 	:	val_out <= 16'hd7f5;
             14'h28e8 	:	val_out <= 16'hd7f9;
             14'h28e9 	:	val_out <= 16'hd7fc;
             14'h28ea 	:	val_out <= 16'hd7ff;
             14'h28eb 	:	val_out <= 16'hd803;
             14'h28ec 	:	val_out <= 16'hd806;
             14'h28ed 	:	val_out <= 16'hd80a;
             14'h28ee 	:	val_out <= 16'hd80d;
             14'h28ef 	:	val_out <= 16'hd810;
             14'h28f0 	:	val_out <= 16'hd814;
             14'h28f1 	:	val_out <= 16'hd817;
             14'h28f2 	:	val_out <= 16'hd81a;
             14'h28f3 	:	val_out <= 16'hd81e;
             14'h28f4 	:	val_out <= 16'hd821;
             14'h28f5 	:	val_out <= 16'hd824;
             14'h28f6 	:	val_out <= 16'hd828;
             14'h28f7 	:	val_out <= 16'hd82b;
             14'h28f8 	:	val_out <= 16'hd82f;
             14'h28f9 	:	val_out <= 16'hd832;
             14'h28fa 	:	val_out <= 16'hd835;
             14'h28fb 	:	val_out <= 16'hd839;
             14'h28fc 	:	val_out <= 16'hd83c;
             14'h28fd 	:	val_out <= 16'hd83f;
             14'h28fe 	:	val_out <= 16'hd843;
             14'h28ff 	:	val_out <= 16'hd846;
             14'h2900 	:	val_out <= 16'hd84a;
             14'h2901 	:	val_out <= 16'hd84d;
             14'h2902 	:	val_out <= 16'hd850;
             14'h2903 	:	val_out <= 16'hd854;
             14'h2904 	:	val_out <= 16'hd857;
             14'h2905 	:	val_out <= 16'hd85a;
             14'h2906 	:	val_out <= 16'hd85e;
             14'h2907 	:	val_out <= 16'hd861;
             14'h2908 	:	val_out <= 16'hd864;
             14'h2909 	:	val_out <= 16'hd868;
             14'h290a 	:	val_out <= 16'hd86b;
             14'h290b 	:	val_out <= 16'hd86e;
             14'h290c 	:	val_out <= 16'hd872;
             14'h290d 	:	val_out <= 16'hd875;
             14'h290e 	:	val_out <= 16'hd879;
             14'h290f 	:	val_out <= 16'hd87c;
             14'h2910 	:	val_out <= 16'hd87f;
             14'h2911 	:	val_out <= 16'hd883;
             14'h2912 	:	val_out <= 16'hd886;
             14'h2913 	:	val_out <= 16'hd889;
             14'h2914 	:	val_out <= 16'hd88d;
             14'h2915 	:	val_out <= 16'hd890;
             14'h2916 	:	val_out <= 16'hd893;
             14'h2917 	:	val_out <= 16'hd897;
             14'h2918 	:	val_out <= 16'hd89a;
             14'h2919 	:	val_out <= 16'hd89d;
             14'h291a 	:	val_out <= 16'hd8a1;
             14'h291b 	:	val_out <= 16'hd8a4;
             14'h291c 	:	val_out <= 16'hd8a7;
             14'h291d 	:	val_out <= 16'hd8ab;
             14'h291e 	:	val_out <= 16'hd8ae;
             14'h291f 	:	val_out <= 16'hd8b1;
             14'h2920 	:	val_out <= 16'hd8b5;
             14'h2921 	:	val_out <= 16'hd8b8;
             14'h2922 	:	val_out <= 16'hd8bb;
             14'h2923 	:	val_out <= 16'hd8bf;
             14'h2924 	:	val_out <= 16'hd8c2;
             14'h2925 	:	val_out <= 16'hd8c6;
             14'h2926 	:	val_out <= 16'hd8c9;
             14'h2927 	:	val_out <= 16'hd8cc;
             14'h2928 	:	val_out <= 16'hd8d0;
             14'h2929 	:	val_out <= 16'hd8d3;
             14'h292a 	:	val_out <= 16'hd8d6;
             14'h292b 	:	val_out <= 16'hd8da;
             14'h292c 	:	val_out <= 16'hd8dd;
             14'h292d 	:	val_out <= 16'hd8e0;
             14'h292e 	:	val_out <= 16'hd8e4;
             14'h292f 	:	val_out <= 16'hd8e7;
             14'h2930 	:	val_out <= 16'hd8ea;
             14'h2931 	:	val_out <= 16'hd8ee;
             14'h2932 	:	val_out <= 16'hd8f1;
             14'h2933 	:	val_out <= 16'hd8f4;
             14'h2934 	:	val_out <= 16'hd8f8;
             14'h2935 	:	val_out <= 16'hd8fb;
             14'h2936 	:	val_out <= 16'hd8fe;
             14'h2937 	:	val_out <= 16'hd902;
             14'h2938 	:	val_out <= 16'hd905;
             14'h2939 	:	val_out <= 16'hd908;
             14'h293a 	:	val_out <= 16'hd90c;
             14'h293b 	:	val_out <= 16'hd90f;
             14'h293c 	:	val_out <= 16'hd912;
             14'h293d 	:	val_out <= 16'hd916;
             14'h293e 	:	val_out <= 16'hd919;
             14'h293f 	:	val_out <= 16'hd91c;
             14'h2940 	:	val_out <= 16'hd920;
             14'h2941 	:	val_out <= 16'hd923;
             14'h2942 	:	val_out <= 16'hd926;
             14'h2943 	:	val_out <= 16'hd92a;
             14'h2944 	:	val_out <= 16'hd92d;
             14'h2945 	:	val_out <= 16'hd930;
             14'h2946 	:	val_out <= 16'hd934;
             14'h2947 	:	val_out <= 16'hd937;
             14'h2948 	:	val_out <= 16'hd93a;
             14'h2949 	:	val_out <= 16'hd93e;
             14'h294a 	:	val_out <= 16'hd941;
             14'h294b 	:	val_out <= 16'hd944;
             14'h294c 	:	val_out <= 16'hd947;
             14'h294d 	:	val_out <= 16'hd94b;
             14'h294e 	:	val_out <= 16'hd94e;
             14'h294f 	:	val_out <= 16'hd951;
             14'h2950 	:	val_out <= 16'hd955;
             14'h2951 	:	val_out <= 16'hd958;
             14'h2952 	:	val_out <= 16'hd95b;
             14'h2953 	:	val_out <= 16'hd95f;
             14'h2954 	:	val_out <= 16'hd962;
             14'h2955 	:	val_out <= 16'hd965;
             14'h2956 	:	val_out <= 16'hd969;
             14'h2957 	:	val_out <= 16'hd96c;
             14'h2958 	:	val_out <= 16'hd96f;
             14'h2959 	:	val_out <= 16'hd973;
             14'h295a 	:	val_out <= 16'hd976;
             14'h295b 	:	val_out <= 16'hd979;
             14'h295c 	:	val_out <= 16'hd97d;
             14'h295d 	:	val_out <= 16'hd980;
             14'h295e 	:	val_out <= 16'hd983;
             14'h295f 	:	val_out <= 16'hd987;
             14'h2960 	:	val_out <= 16'hd98a;
             14'h2961 	:	val_out <= 16'hd98d;
             14'h2962 	:	val_out <= 16'hd990;
             14'h2963 	:	val_out <= 16'hd994;
             14'h2964 	:	val_out <= 16'hd997;
             14'h2965 	:	val_out <= 16'hd99a;
             14'h2966 	:	val_out <= 16'hd99e;
             14'h2967 	:	val_out <= 16'hd9a1;
             14'h2968 	:	val_out <= 16'hd9a4;
             14'h2969 	:	val_out <= 16'hd9a8;
             14'h296a 	:	val_out <= 16'hd9ab;
             14'h296b 	:	val_out <= 16'hd9ae;
             14'h296c 	:	val_out <= 16'hd9b2;
             14'h296d 	:	val_out <= 16'hd9b5;
             14'h296e 	:	val_out <= 16'hd9b8;
             14'h296f 	:	val_out <= 16'hd9bb;
             14'h2970 	:	val_out <= 16'hd9bf;
             14'h2971 	:	val_out <= 16'hd9c2;
             14'h2972 	:	val_out <= 16'hd9c5;
             14'h2973 	:	val_out <= 16'hd9c9;
             14'h2974 	:	val_out <= 16'hd9cc;
             14'h2975 	:	val_out <= 16'hd9cf;
             14'h2976 	:	val_out <= 16'hd9d3;
             14'h2977 	:	val_out <= 16'hd9d6;
             14'h2978 	:	val_out <= 16'hd9d9;
             14'h2979 	:	val_out <= 16'hd9dc;
             14'h297a 	:	val_out <= 16'hd9e0;
             14'h297b 	:	val_out <= 16'hd9e3;
             14'h297c 	:	val_out <= 16'hd9e6;
             14'h297d 	:	val_out <= 16'hd9ea;
             14'h297e 	:	val_out <= 16'hd9ed;
             14'h297f 	:	val_out <= 16'hd9f0;
             14'h2980 	:	val_out <= 16'hd9f4;
             14'h2981 	:	val_out <= 16'hd9f7;
             14'h2982 	:	val_out <= 16'hd9fa;
             14'h2983 	:	val_out <= 16'hd9fd;
             14'h2984 	:	val_out <= 16'hda01;
             14'h2985 	:	val_out <= 16'hda04;
             14'h2986 	:	val_out <= 16'hda07;
             14'h2987 	:	val_out <= 16'hda0b;
             14'h2988 	:	val_out <= 16'hda0e;
             14'h2989 	:	val_out <= 16'hda11;
             14'h298a 	:	val_out <= 16'hda14;
             14'h298b 	:	val_out <= 16'hda18;
             14'h298c 	:	val_out <= 16'hda1b;
             14'h298d 	:	val_out <= 16'hda1e;
             14'h298e 	:	val_out <= 16'hda22;
             14'h298f 	:	val_out <= 16'hda25;
             14'h2990 	:	val_out <= 16'hda28;
             14'h2991 	:	val_out <= 16'hda2c;
             14'h2992 	:	val_out <= 16'hda2f;
             14'h2993 	:	val_out <= 16'hda32;
             14'h2994 	:	val_out <= 16'hda35;
             14'h2995 	:	val_out <= 16'hda39;
             14'h2996 	:	val_out <= 16'hda3c;
             14'h2997 	:	val_out <= 16'hda3f;
             14'h2998 	:	val_out <= 16'hda43;
             14'h2999 	:	val_out <= 16'hda46;
             14'h299a 	:	val_out <= 16'hda49;
             14'h299b 	:	val_out <= 16'hda4c;
             14'h299c 	:	val_out <= 16'hda50;
             14'h299d 	:	val_out <= 16'hda53;
             14'h299e 	:	val_out <= 16'hda56;
             14'h299f 	:	val_out <= 16'hda59;
             14'h29a0 	:	val_out <= 16'hda5d;
             14'h29a1 	:	val_out <= 16'hda60;
             14'h29a2 	:	val_out <= 16'hda63;
             14'h29a3 	:	val_out <= 16'hda67;
             14'h29a4 	:	val_out <= 16'hda6a;
             14'h29a5 	:	val_out <= 16'hda6d;
             14'h29a6 	:	val_out <= 16'hda70;
             14'h29a7 	:	val_out <= 16'hda74;
             14'h29a8 	:	val_out <= 16'hda77;
             14'h29a9 	:	val_out <= 16'hda7a;
             14'h29aa 	:	val_out <= 16'hda7e;
             14'h29ab 	:	val_out <= 16'hda81;
             14'h29ac 	:	val_out <= 16'hda84;
             14'h29ad 	:	val_out <= 16'hda87;
             14'h29ae 	:	val_out <= 16'hda8b;
             14'h29af 	:	val_out <= 16'hda8e;
             14'h29b0 	:	val_out <= 16'hda91;
             14'h29b1 	:	val_out <= 16'hda94;
             14'h29b2 	:	val_out <= 16'hda98;
             14'h29b3 	:	val_out <= 16'hda9b;
             14'h29b4 	:	val_out <= 16'hda9e;
             14'h29b5 	:	val_out <= 16'hdaa2;
             14'h29b6 	:	val_out <= 16'hdaa5;
             14'h29b7 	:	val_out <= 16'hdaa8;
             14'h29b8 	:	val_out <= 16'hdaab;
             14'h29b9 	:	val_out <= 16'hdaaf;
             14'h29ba 	:	val_out <= 16'hdab2;
             14'h29bb 	:	val_out <= 16'hdab5;
             14'h29bc 	:	val_out <= 16'hdab8;
             14'h29bd 	:	val_out <= 16'hdabc;
             14'h29be 	:	val_out <= 16'hdabf;
             14'h29bf 	:	val_out <= 16'hdac2;
             14'h29c0 	:	val_out <= 16'hdac5;
             14'h29c1 	:	val_out <= 16'hdac9;
             14'h29c2 	:	val_out <= 16'hdacc;
             14'h29c3 	:	val_out <= 16'hdacf;
             14'h29c4 	:	val_out <= 16'hdad2;
             14'h29c5 	:	val_out <= 16'hdad6;
             14'h29c6 	:	val_out <= 16'hdad9;
             14'h29c7 	:	val_out <= 16'hdadc;
             14'h29c8 	:	val_out <= 16'hdae0;
             14'h29c9 	:	val_out <= 16'hdae3;
             14'h29ca 	:	val_out <= 16'hdae6;
             14'h29cb 	:	val_out <= 16'hdae9;
             14'h29cc 	:	val_out <= 16'hdaed;
             14'h29cd 	:	val_out <= 16'hdaf0;
             14'h29ce 	:	val_out <= 16'hdaf3;
             14'h29cf 	:	val_out <= 16'hdaf6;
             14'h29d0 	:	val_out <= 16'hdafa;
             14'h29d1 	:	val_out <= 16'hdafd;
             14'h29d2 	:	val_out <= 16'hdb00;
             14'h29d3 	:	val_out <= 16'hdb03;
             14'h29d4 	:	val_out <= 16'hdb07;
             14'h29d5 	:	val_out <= 16'hdb0a;
             14'h29d6 	:	val_out <= 16'hdb0d;
             14'h29d7 	:	val_out <= 16'hdb10;
             14'h29d8 	:	val_out <= 16'hdb14;
             14'h29d9 	:	val_out <= 16'hdb17;
             14'h29da 	:	val_out <= 16'hdb1a;
             14'h29db 	:	val_out <= 16'hdb1d;
             14'h29dc 	:	val_out <= 16'hdb21;
             14'h29dd 	:	val_out <= 16'hdb24;
             14'h29de 	:	val_out <= 16'hdb27;
             14'h29df 	:	val_out <= 16'hdb2a;
             14'h29e0 	:	val_out <= 16'hdb2e;
             14'h29e1 	:	val_out <= 16'hdb31;
             14'h29e2 	:	val_out <= 16'hdb34;
             14'h29e3 	:	val_out <= 16'hdb37;
             14'h29e4 	:	val_out <= 16'hdb3b;
             14'h29e5 	:	val_out <= 16'hdb3e;
             14'h29e6 	:	val_out <= 16'hdb41;
             14'h29e7 	:	val_out <= 16'hdb44;
             14'h29e8 	:	val_out <= 16'hdb48;
             14'h29e9 	:	val_out <= 16'hdb4b;
             14'h29ea 	:	val_out <= 16'hdb4e;
             14'h29eb 	:	val_out <= 16'hdb51;
             14'h29ec 	:	val_out <= 16'hdb55;
             14'h29ed 	:	val_out <= 16'hdb58;
             14'h29ee 	:	val_out <= 16'hdb5b;
             14'h29ef 	:	val_out <= 16'hdb5e;
             14'h29f0 	:	val_out <= 16'hdb61;
             14'h29f1 	:	val_out <= 16'hdb65;
             14'h29f2 	:	val_out <= 16'hdb68;
             14'h29f3 	:	val_out <= 16'hdb6b;
             14'h29f4 	:	val_out <= 16'hdb6e;
             14'h29f5 	:	val_out <= 16'hdb72;
             14'h29f6 	:	val_out <= 16'hdb75;
             14'h29f7 	:	val_out <= 16'hdb78;
             14'h29f8 	:	val_out <= 16'hdb7b;
             14'h29f9 	:	val_out <= 16'hdb7f;
             14'h29fa 	:	val_out <= 16'hdb82;
             14'h29fb 	:	val_out <= 16'hdb85;
             14'h29fc 	:	val_out <= 16'hdb88;
             14'h29fd 	:	val_out <= 16'hdb8c;
             14'h29fe 	:	val_out <= 16'hdb8f;
             14'h29ff 	:	val_out <= 16'hdb92;
             14'h2a00 	:	val_out <= 16'hdb95;
             14'h2a01 	:	val_out <= 16'hdb98;
             14'h2a02 	:	val_out <= 16'hdb9c;
             14'h2a03 	:	val_out <= 16'hdb9f;
             14'h2a04 	:	val_out <= 16'hdba2;
             14'h2a05 	:	val_out <= 16'hdba5;
             14'h2a06 	:	val_out <= 16'hdba9;
             14'h2a07 	:	val_out <= 16'hdbac;
             14'h2a08 	:	val_out <= 16'hdbaf;
             14'h2a09 	:	val_out <= 16'hdbb2;
             14'h2a0a 	:	val_out <= 16'hdbb5;
             14'h2a0b 	:	val_out <= 16'hdbb9;
             14'h2a0c 	:	val_out <= 16'hdbbc;
             14'h2a0d 	:	val_out <= 16'hdbbf;
             14'h2a0e 	:	val_out <= 16'hdbc2;
             14'h2a0f 	:	val_out <= 16'hdbc6;
             14'h2a10 	:	val_out <= 16'hdbc9;
             14'h2a11 	:	val_out <= 16'hdbcc;
             14'h2a12 	:	val_out <= 16'hdbcf;
             14'h2a13 	:	val_out <= 16'hdbd2;
             14'h2a14 	:	val_out <= 16'hdbd6;
             14'h2a15 	:	val_out <= 16'hdbd9;
             14'h2a16 	:	val_out <= 16'hdbdc;
             14'h2a17 	:	val_out <= 16'hdbdf;
             14'h2a18 	:	val_out <= 16'hdbe3;
             14'h2a19 	:	val_out <= 16'hdbe6;
             14'h2a1a 	:	val_out <= 16'hdbe9;
             14'h2a1b 	:	val_out <= 16'hdbec;
             14'h2a1c 	:	val_out <= 16'hdbef;
             14'h2a1d 	:	val_out <= 16'hdbf3;
             14'h2a1e 	:	val_out <= 16'hdbf6;
             14'h2a1f 	:	val_out <= 16'hdbf9;
             14'h2a20 	:	val_out <= 16'hdbfc;
             14'h2a21 	:	val_out <= 16'hdc00;
             14'h2a22 	:	val_out <= 16'hdc03;
             14'h2a23 	:	val_out <= 16'hdc06;
             14'h2a24 	:	val_out <= 16'hdc09;
             14'h2a25 	:	val_out <= 16'hdc0c;
             14'h2a26 	:	val_out <= 16'hdc10;
             14'h2a27 	:	val_out <= 16'hdc13;
             14'h2a28 	:	val_out <= 16'hdc16;
             14'h2a29 	:	val_out <= 16'hdc19;
             14'h2a2a 	:	val_out <= 16'hdc1c;
             14'h2a2b 	:	val_out <= 16'hdc20;
             14'h2a2c 	:	val_out <= 16'hdc23;
             14'h2a2d 	:	val_out <= 16'hdc26;
             14'h2a2e 	:	val_out <= 16'hdc29;
             14'h2a2f 	:	val_out <= 16'hdc2c;
             14'h2a30 	:	val_out <= 16'hdc30;
             14'h2a31 	:	val_out <= 16'hdc33;
             14'h2a32 	:	val_out <= 16'hdc36;
             14'h2a33 	:	val_out <= 16'hdc39;
             14'h2a34 	:	val_out <= 16'hdc3c;
             14'h2a35 	:	val_out <= 16'hdc40;
             14'h2a36 	:	val_out <= 16'hdc43;
             14'h2a37 	:	val_out <= 16'hdc46;
             14'h2a38 	:	val_out <= 16'hdc49;
             14'h2a39 	:	val_out <= 16'hdc4c;
             14'h2a3a 	:	val_out <= 16'hdc50;
             14'h2a3b 	:	val_out <= 16'hdc53;
             14'h2a3c 	:	val_out <= 16'hdc56;
             14'h2a3d 	:	val_out <= 16'hdc59;
             14'h2a3e 	:	val_out <= 16'hdc5c;
             14'h2a3f 	:	val_out <= 16'hdc60;
             14'h2a40 	:	val_out <= 16'hdc63;
             14'h2a41 	:	val_out <= 16'hdc66;
             14'h2a42 	:	val_out <= 16'hdc69;
             14'h2a43 	:	val_out <= 16'hdc6c;
             14'h2a44 	:	val_out <= 16'hdc70;
             14'h2a45 	:	val_out <= 16'hdc73;
             14'h2a46 	:	val_out <= 16'hdc76;
             14'h2a47 	:	val_out <= 16'hdc79;
             14'h2a48 	:	val_out <= 16'hdc7c;
             14'h2a49 	:	val_out <= 16'hdc80;
             14'h2a4a 	:	val_out <= 16'hdc83;
             14'h2a4b 	:	val_out <= 16'hdc86;
             14'h2a4c 	:	val_out <= 16'hdc89;
             14'h2a4d 	:	val_out <= 16'hdc8c;
             14'h2a4e 	:	val_out <= 16'hdc90;
             14'h2a4f 	:	val_out <= 16'hdc93;
             14'h2a50 	:	val_out <= 16'hdc96;
             14'h2a51 	:	val_out <= 16'hdc99;
             14'h2a52 	:	val_out <= 16'hdc9c;
             14'h2a53 	:	val_out <= 16'hdca0;
             14'h2a54 	:	val_out <= 16'hdca3;
             14'h2a55 	:	val_out <= 16'hdca6;
             14'h2a56 	:	val_out <= 16'hdca9;
             14'h2a57 	:	val_out <= 16'hdcac;
             14'h2a58 	:	val_out <= 16'hdcaf;
             14'h2a59 	:	val_out <= 16'hdcb3;
             14'h2a5a 	:	val_out <= 16'hdcb6;
             14'h2a5b 	:	val_out <= 16'hdcb9;
             14'h2a5c 	:	val_out <= 16'hdcbc;
             14'h2a5d 	:	val_out <= 16'hdcbf;
             14'h2a5e 	:	val_out <= 16'hdcc3;
             14'h2a5f 	:	val_out <= 16'hdcc6;
             14'h2a60 	:	val_out <= 16'hdcc9;
             14'h2a61 	:	val_out <= 16'hdccc;
             14'h2a62 	:	val_out <= 16'hdccf;
             14'h2a63 	:	val_out <= 16'hdcd2;
             14'h2a64 	:	val_out <= 16'hdcd6;
             14'h2a65 	:	val_out <= 16'hdcd9;
             14'h2a66 	:	val_out <= 16'hdcdc;
             14'h2a67 	:	val_out <= 16'hdcdf;
             14'h2a68 	:	val_out <= 16'hdce2;
             14'h2a69 	:	val_out <= 16'hdce6;
             14'h2a6a 	:	val_out <= 16'hdce9;
             14'h2a6b 	:	val_out <= 16'hdcec;
             14'h2a6c 	:	val_out <= 16'hdcef;
             14'h2a6d 	:	val_out <= 16'hdcf2;
             14'h2a6e 	:	val_out <= 16'hdcf5;
             14'h2a6f 	:	val_out <= 16'hdcf9;
             14'h2a70 	:	val_out <= 16'hdcfc;
             14'h2a71 	:	val_out <= 16'hdcff;
             14'h2a72 	:	val_out <= 16'hdd02;
             14'h2a73 	:	val_out <= 16'hdd05;
             14'h2a74 	:	val_out <= 16'hdd08;
             14'h2a75 	:	val_out <= 16'hdd0c;
             14'h2a76 	:	val_out <= 16'hdd0f;
             14'h2a77 	:	val_out <= 16'hdd12;
             14'h2a78 	:	val_out <= 16'hdd15;
             14'h2a79 	:	val_out <= 16'hdd18;
             14'h2a7a 	:	val_out <= 16'hdd1b;
             14'h2a7b 	:	val_out <= 16'hdd1f;
             14'h2a7c 	:	val_out <= 16'hdd22;
             14'h2a7d 	:	val_out <= 16'hdd25;
             14'h2a7e 	:	val_out <= 16'hdd28;
             14'h2a7f 	:	val_out <= 16'hdd2b;
             14'h2a80 	:	val_out <= 16'hdd2e;
             14'h2a81 	:	val_out <= 16'hdd32;
             14'h2a82 	:	val_out <= 16'hdd35;
             14'h2a83 	:	val_out <= 16'hdd38;
             14'h2a84 	:	val_out <= 16'hdd3b;
             14'h2a85 	:	val_out <= 16'hdd3e;
             14'h2a86 	:	val_out <= 16'hdd41;
             14'h2a87 	:	val_out <= 16'hdd45;
             14'h2a88 	:	val_out <= 16'hdd48;
             14'h2a89 	:	val_out <= 16'hdd4b;
             14'h2a8a 	:	val_out <= 16'hdd4e;
             14'h2a8b 	:	val_out <= 16'hdd51;
             14'h2a8c 	:	val_out <= 16'hdd54;
             14'h2a8d 	:	val_out <= 16'hdd57;
             14'h2a8e 	:	val_out <= 16'hdd5b;
             14'h2a8f 	:	val_out <= 16'hdd5e;
             14'h2a90 	:	val_out <= 16'hdd61;
             14'h2a91 	:	val_out <= 16'hdd64;
             14'h2a92 	:	val_out <= 16'hdd67;
             14'h2a93 	:	val_out <= 16'hdd6a;
             14'h2a94 	:	val_out <= 16'hdd6e;
             14'h2a95 	:	val_out <= 16'hdd71;
             14'h2a96 	:	val_out <= 16'hdd74;
             14'h2a97 	:	val_out <= 16'hdd77;
             14'h2a98 	:	val_out <= 16'hdd7a;
             14'h2a99 	:	val_out <= 16'hdd7d;
             14'h2a9a 	:	val_out <= 16'hdd80;
             14'h2a9b 	:	val_out <= 16'hdd84;
             14'h2a9c 	:	val_out <= 16'hdd87;
             14'h2a9d 	:	val_out <= 16'hdd8a;
             14'h2a9e 	:	val_out <= 16'hdd8d;
             14'h2a9f 	:	val_out <= 16'hdd90;
             14'h2aa0 	:	val_out <= 16'hdd93;
             14'h2aa1 	:	val_out <= 16'hdd97;
             14'h2aa2 	:	val_out <= 16'hdd9a;
             14'h2aa3 	:	val_out <= 16'hdd9d;
             14'h2aa4 	:	val_out <= 16'hdda0;
             14'h2aa5 	:	val_out <= 16'hdda3;
             14'h2aa6 	:	val_out <= 16'hdda6;
             14'h2aa7 	:	val_out <= 16'hdda9;
             14'h2aa8 	:	val_out <= 16'hddad;
             14'h2aa9 	:	val_out <= 16'hddb0;
             14'h2aaa 	:	val_out <= 16'hddb3;
             14'h2aab 	:	val_out <= 16'hddb6;
             14'h2aac 	:	val_out <= 16'hddb9;
             14'h2aad 	:	val_out <= 16'hddbc;
             14'h2aae 	:	val_out <= 16'hddbf;
             14'h2aaf 	:	val_out <= 16'hddc3;
             14'h2ab0 	:	val_out <= 16'hddc6;
             14'h2ab1 	:	val_out <= 16'hddc9;
             14'h2ab2 	:	val_out <= 16'hddcc;
             14'h2ab3 	:	val_out <= 16'hddcf;
             14'h2ab4 	:	val_out <= 16'hddd2;
             14'h2ab5 	:	val_out <= 16'hddd5;
             14'h2ab6 	:	val_out <= 16'hddd8;
             14'h2ab7 	:	val_out <= 16'hdddc;
             14'h2ab8 	:	val_out <= 16'hdddf;
             14'h2ab9 	:	val_out <= 16'hdde2;
             14'h2aba 	:	val_out <= 16'hdde5;
             14'h2abb 	:	val_out <= 16'hdde8;
             14'h2abc 	:	val_out <= 16'hddeb;
             14'h2abd 	:	val_out <= 16'hddee;
             14'h2abe 	:	val_out <= 16'hddf2;
             14'h2abf 	:	val_out <= 16'hddf5;
             14'h2ac0 	:	val_out <= 16'hddf8;
             14'h2ac1 	:	val_out <= 16'hddfb;
             14'h2ac2 	:	val_out <= 16'hddfe;
             14'h2ac3 	:	val_out <= 16'hde01;
             14'h2ac4 	:	val_out <= 16'hde04;
             14'h2ac5 	:	val_out <= 16'hde07;
             14'h2ac6 	:	val_out <= 16'hde0b;
             14'h2ac7 	:	val_out <= 16'hde0e;
             14'h2ac8 	:	val_out <= 16'hde11;
             14'h2ac9 	:	val_out <= 16'hde14;
             14'h2aca 	:	val_out <= 16'hde17;
             14'h2acb 	:	val_out <= 16'hde1a;
             14'h2acc 	:	val_out <= 16'hde1d;
             14'h2acd 	:	val_out <= 16'hde20;
             14'h2ace 	:	val_out <= 16'hde24;
             14'h2acf 	:	val_out <= 16'hde27;
             14'h2ad0 	:	val_out <= 16'hde2a;
             14'h2ad1 	:	val_out <= 16'hde2d;
             14'h2ad2 	:	val_out <= 16'hde30;
             14'h2ad3 	:	val_out <= 16'hde33;
             14'h2ad4 	:	val_out <= 16'hde36;
             14'h2ad5 	:	val_out <= 16'hde39;
             14'h2ad6 	:	val_out <= 16'hde3d;
             14'h2ad7 	:	val_out <= 16'hde40;
             14'h2ad8 	:	val_out <= 16'hde43;
             14'h2ad9 	:	val_out <= 16'hde46;
             14'h2ada 	:	val_out <= 16'hde49;
             14'h2adb 	:	val_out <= 16'hde4c;
             14'h2adc 	:	val_out <= 16'hde4f;
             14'h2add 	:	val_out <= 16'hde52;
             14'h2ade 	:	val_out <= 16'hde55;
             14'h2adf 	:	val_out <= 16'hde59;
             14'h2ae0 	:	val_out <= 16'hde5c;
             14'h2ae1 	:	val_out <= 16'hde5f;
             14'h2ae2 	:	val_out <= 16'hde62;
             14'h2ae3 	:	val_out <= 16'hde65;
             14'h2ae4 	:	val_out <= 16'hde68;
             14'h2ae5 	:	val_out <= 16'hde6b;
             14'h2ae6 	:	val_out <= 16'hde6e;
             14'h2ae7 	:	val_out <= 16'hde71;
             14'h2ae8 	:	val_out <= 16'hde75;
             14'h2ae9 	:	val_out <= 16'hde78;
             14'h2aea 	:	val_out <= 16'hde7b;
             14'h2aeb 	:	val_out <= 16'hde7e;
             14'h2aec 	:	val_out <= 16'hde81;
             14'h2aed 	:	val_out <= 16'hde84;
             14'h2aee 	:	val_out <= 16'hde87;
             14'h2aef 	:	val_out <= 16'hde8a;
             14'h2af0 	:	val_out <= 16'hde8d;
             14'h2af1 	:	val_out <= 16'hde91;
             14'h2af2 	:	val_out <= 16'hde94;
             14'h2af3 	:	val_out <= 16'hde97;
             14'h2af4 	:	val_out <= 16'hde9a;
             14'h2af5 	:	val_out <= 16'hde9d;
             14'h2af6 	:	val_out <= 16'hdea0;
             14'h2af7 	:	val_out <= 16'hdea3;
             14'h2af8 	:	val_out <= 16'hdea6;
             14'h2af9 	:	val_out <= 16'hdea9;
             14'h2afa 	:	val_out <= 16'hdeac;
             14'h2afb 	:	val_out <= 16'hdeb0;
             14'h2afc 	:	val_out <= 16'hdeb3;
             14'h2afd 	:	val_out <= 16'hdeb6;
             14'h2afe 	:	val_out <= 16'hdeb9;
             14'h2aff 	:	val_out <= 16'hdebc;
             14'h2b00 	:	val_out <= 16'hdebf;
             14'h2b01 	:	val_out <= 16'hdec2;
             14'h2b02 	:	val_out <= 16'hdec5;
             14'h2b03 	:	val_out <= 16'hdec8;
             14'h2b04 	:	val_out <= 16'hdecb;
             14'h2b05 	:	val_out <= 16'hdecf;
             14'h2b06 	:	val_out <= 16'hded2;
             14'h2b07 	:	val_out <= 16'hded5;
             14'h2b08 	:	val_out <= 16'hded8;
             14'h2b09 	:	val_out <= 16'hdedb;
             14'h2b0a 	:	val_out <= 16'hdede;
             14'h2b0b 	:	val_out <= 16'hdee1;
             14'h2b0c 	:	val_out <= 16'hdee4;
             14'h2b0d 	:	val_out <= 16'hdee7;
             14'h2b0e 	:	val_out <= 16'hdeea;
             14'h2b0f 	:	val_out <= 16'hdeed;
             14'h2b10 	:	val_out <= 16'hdef1;
             14'h2b11 	:	val_out <= 16'hdef4;
             14'h2b12 	:	val_out <= 16'hdef7;
             14'h2b13 	:	val_out <= 16'hdefa;
             14'h2b14 	:	val_out <= 16'hdefd;
             14'h2b15 	:	val_out <= 16'hdf00;
             14'h2b16 	:	val_out <= 16'hdf03;
             14'h2b17 	:	val_out <= 16'hdf06;
             14'h2b18 	:	val_out <= 16'hdf09;
             14'h2b19 	:	val_out <= 16'hdf0c;
             14'h2b1a 	:	val_out <= 16'hdf0f;
             14'h2b1b 	:	val_out <= 16'hdf12;
             14'h2b1c 	:	val_out <= 16'hdf16;
             14'h2b1d 	:	val_out <= 16'hdf19;
             14'h2b1e 	:	val_out <= 16'hdf1c;
             14'h2b1f 	:	val_out <= 16'hdf1f;
             14'h2b20 	:	val_out <= 16'hdf22;
             14'h2b21 	:	val_out <= 16'hdf25;
             14'h2b22 	:	val_out <= 16'hdf28;
             14'h2b23 	:	val_out <= 16'hdf2b;
             14'h2b24 	:	val_out <= 16'hdf2e;
             14'h2b25 	:	val_out <= 16'hdf31;
             14'h2b26 	:	val_out <= 16'hdf34;
             14'h2b27 	:	val_out <= 16'hdf37;
             14'h2b28 	:	val_out <= 16'hdf3b;
             14'h2b29 	:	val_out <= 16'hdf3e;
             14'h2b2a 	:	val_out <= 16'hdf41;
             14'h2b2b 	:	val_out <= 16'hdf44;
             14'h2b2c 	:	val_out <= 16'hdf47;
             14'h2b2d 	:	val_out <= 16'hdf4a;
             14'h2b2e 	:	val_out <= 16'hdf4d;
             14'h2b2f 	:	val_out <= 16'hdf50;
             14'h2b30 	:	val_out <= 16'hdf53;
             14'h2b31 	:	val_out <= 16'hdf56;
             14'h2b32 	:	val_out <= 16'hdf59;
             14'h2b33 	:	val_out <= 16'hdf5c;
             14'h2b34 	:	val_out <= 16'hdf5f;
             14'h2b35 	:	val_out <= 16'hdf62;
             14'h2b36 	:	val_out <= 16'hdf66;
             14'h2b37 	:	val_out <= 16'hdf69;
             14'h2b38 	:	val_out <= 16'hdf6c;
             14'h2b39 	:	val_out <= 16'hdf6f;
             14'h2b3a 	:	val_out <= 16'hdf72;
             14'h2b3b 	:	val_out <= 16'hdf75;
             14'h2b3c 	:	val_out <= 16'hdf78;
             14'h2b3d 	:	val_out <= 16'hdf7b;
             14'h2b3e 	:	val_out <= 16'hdf7e;
             14'h2b3f 	:	val_out <= 16'hdf81;
             14'h2b40 	:	val_out <= 16'hdf84;
             14'h2b41 	:	val_out <= 16'hdf87;
             14'h2b42 	:	val_out <= 16'hdf8a;
             14'h2b43 	:	val_out <= 16'hdf8d;
             14'h2b44 	:	val_out <= 16'hdf90;
             14'h2b45 	:	val_out <= 16'hdf93;
             14'h2b46 	:	val_out <= 16'hdf97;
             14'h2b47 	:	val_out <= 16'hdf9a;
             14'h2b48 	:	val_out <= 16'hdf9d;
             14'h2b49 	:	val_out <= 16'hdfa0;
             14'h2b4a 	:	val_out <= 16'hdfa3;
             14'h2b4b 	:	val_out <= 16'hdfa6;
             14'h2b4c 	:	val_out <= 16'hdfa9;
             14'h2b4d 	:	val_out <= 16'hdfac;
             14'h2b4e 	:	val_out <= 16'hdfaf;
             14'h2b4f 	:	val_out <= 16'hdfb2;
             14'h2b50 	:	val_out <= 16'hdfb5;
             14'h2b51 	:	val_out <= 16'hdfb8;
             14'h2b52 	:	val_out <= 16'hdfbb;
             14'h2b53 	:	val_out <= 16'hdfbe;
             14'h2b54 	:	val_out <= 16'hdfc1;
             14'h2b55 	:	val_out <= 16'hdfc4;
             14'h2b56 	:	val_out <= 16'hdfc7;
             14'h2b57 	:	val_out <= 16'hdfca;
             14'h2b58 	:	val_out <= 16'hdfce;
             14'h2b59 	:	val_out <= 16'hdfd1;
             14'h2b5a 	:	val_out <= 16'hdfd4;
             14'h2b5b 	:	val_out <= 16'hdfd7;
             14'h2b5c 	:	val_out <= 16'hdfda;
             14'h2b5d 	:	val_out <= 16'hdfdd;
             14'h2b5e 	:	val_out <= 16'hdfe0;
             14'h2b5f 	:	val_out <= 16'hdfe3;
             14'h2b60 	:	val_out <= 16'hdfe6;
             14'h2b61 	:	val_out <= 16'hdfe9;
             14'h2b62 	:	val_out <= 16'hdfec;
             14'h2b63 	:	val_out <= 16'hdfef;
             14'h2b64 	:	val_out <= 16'hdff2;
             14'h2b65 	:	val_out <= 16'hdff5;
             14'h2b66 	:	val_out <= 16'hdff8;
             14'h2b67 	:	val_out <= 16'hdffb;
             14'h2b68 	:	val_out <= 16'hdffe;
             14'h2b69 	:	val_out <= 16'he001;
             14'h2b6a 	:	val_out <= 16'he004;
             14'h2b6b 	:	val_out <= 16'he007;
             14'h2b6c 	:	val_out <= 16'he00a;
             14'h2b6d 	:	val_out <= 16'he00d;
             14'h2b6e 	:	val_out <= 16'he011;
             14'h2b6f 	:	val_out <= 16'he014;
             14'h2b70 	:	val_out <= 16'he017;
             14'h2b71 	:	val_out <= 16'he01a;
             14'h2b72 	:	val_out <= 16'he01d;
             14'h2b73 	:	val_out <= 16'he020;
             14'h2b74 	:	val_out <= 16'he023;
             14'h2b75 	:	val_out <= 16'he026;
             14'h2b76 	:	val_out <= 16'he029;
             14'h2b77 	:	val_out <= 16'he02c;
             14'h2b78 	:	val_out <= 16'he02f;
             14'h2b79 	:	val_out <= 16'he032;
             14'h2b7a 	:	val_out <= 16'he035;
             14'h2b7b 	:	val_out <= 16'he038;
             14'h2b7c 	:	val_out <= 16'he03b;
             14'h2b7d 	:	val_out <= 16'he03e;
             14'h2b7e 	:	val_out <= 16'he041;
             14'h2b7f 	:	val_out <= 16'he044;
             14'h2b80 	:	val_out <= 16'he047;
             14'h2b81 	:	val_out <= 16'he04a;
             14'h2b82 	:	val_out <= 16'he04d;
             14'h2b83 	:	val_out <= 16'he050;
             14'h2b84 	:	val_out <= 16'he053;
             14'h2b85 	:	val_out <= 16'he056;
             14'h2b86 	:	val_out <= 16'he059;
             14'h2b87 	:	val_out <= 16'he05c;
             14'h2b88 	:	val_out <= 16'he05f;
             14'h2b89 	:	val_out <= 16'he062;
             14'h2b8a 	:	val_out <= 16'he065;
             14'h2b8b 	:	val_out <= 16'he068;
             14'h2b8c 	:	val_out <= 16'he06b;
             14'h2b8d 	:	val_out <= 16'he06e;
             14'h2b8e 	:	val_out <= 16'he072;
             14'h2b8f 	:	val_out <= 16'he075;
             14'h2b90 	:	val_out <= 16'he078;
             14'h2b91 	:	val_out <= 16'he07b;
             14'h2b92 	:	val_out <= 16'he07e;
             14'h2b93 	:	val_out <= 16'he081;
             14'h2b94 	:	val_out <= 16'he084;
             14'h2b95 	:	val_out <= 16'he087;
             14'h2b96 	:	val_out <= 16'he08a;
             14'h2b97 	:	val_out <= 16'he08d;
             14'h2b98 	:	val_out <= 16'he090;
             14'h2b99 	:	val_out <= 16'he093;
             14'h2b9a 	:	val_out <= 16'he096;
             14'h2b9b 	:	val_out <= 16'he099;
             14'h2b9c 	:	val_out <= 16'he09c;
             14'h2b9d 	:	val_out <= 16'he09f;
             14'h2b9e 	:	val_out <= 16'he0a2;
             14'h2b9f 	:	val_out <= 16'he0a5;
             14'h2ba0 	:	val_out <= 16'he0a8;
             14'h2ba1 	:	val_out <= 16'he0ab;
             14'h2ba2 	:	val_out <= 16'he0ae;
             14'h2ba3 	:	val_out <= 16'he0b1;
             14'h2ba4 	:	val_out <= 16'he0b4;
             14'h2ba5 	:	val_out <= 16'he0b7;
             14'h2ba6 	:	val_out <= 16'he0ba;
             14'h2ba7 	:	val_out <= 16'he0bd;
             14'h2ba8 	:	val_out <= 16'he0c0;
             14'h2ba9 	:	val_out <= 16'he0c3;
             14'h2baa 	:	val_out <= 16'he0c6;
             14'h2bab 	:	val_out <= 16'he0c9;
             14'h2bac 	:	val_out <= 16'he0cc;
             14'h2bad 	:	val_out <= 16'he0cf;
             14'h2bae 	:	val_out <= 16'he0d2;
             14'h2baf 	:	val_out <= 16'he0d5;
             14'h2bb0 	:	val_out <= 16'he0d8;
             14'h2bb1 	:	val_out <= 16'he0db;
             14'h2bb2 	:	val_out <= 16'he0de;
             14'h2bb3 	:	val_out <= 16'he0e1;
             14'h2bb4 	:	val_out <= 16'he0e4;
             14'h2bb5 	:	val_out <= 16'he0e7;
             14'h2bb6 	:	val_out <= 16'he0ea;
             14'h2bb7 	:	val_out <= 16'he0ed;
             14'h2bb8 	:	val_out <= 16'he0f0;
             14'h2bb9 	:	val_out <= 16'he0f3;
             14'h2bba 	:	val_out <= 16'he0f6;
             14'h2bbb 	:	val_out <= 16'he0f9;
             14'h2bbc 	:	val_out <= 16'he0fc;
             14'h2bbd 	:	val_out <= 16'he0ff;
             14'h2bbe 	:	val_out <= 16'he102;
             14'h2bbf 	:	val_out <= 16'he105;
             14'h2bc0 	:	val_out <= 16'he108;
             14'h2bc1 	:	val_out <= 16'he10b;
             14'h2bc2 	:	val_out <= 16'he10e;
             14'h2bc3 	:	val_out <= 16'he111;
             14'h2bc4 	:	val_out <= 16'he114;
             14'h2bc5 	:	val_out <= 16'he117;
             14'h2bc6 	:	val_out <= 16'he11a;
             14'h2bc7 	:	val_out <= 16'he11d;
             14'h2bc8 	:	val_out <= 16'he120;
             14'h2bc9 	:	val_out <= 16'he123;
             14'h2bca 	:	val_out <= 16'he126;
             14'h2bcb 	:	val_out <= 16'he129;
             14'h2bcc 	:	val_out <= 16'he12c;
             14'h2bcd 	:	val_out <= 16'he12f;
             14'h2bce 	:	val_out <= 16'he132;
             14'h2bcf 	:	val_out <= 16'he135;
             14'h2bd0 	:	val_out <= 16'he138;
             14'h2bd1 	:	val_out <= 16'he13b;
             14'h2bd2 	:	val_out <= 16'he13e;
             14'h2bd3 	:	val_out <= 16'he141;
             14'h2bd4 	:	val_out <= 16'he144;
             14'h2bd5 	:	val_out <= 16'he147;
             14'h2bd6 	:	val_out <= 16'he14a;
             14'h2bd7 	:	val_out <= 16'he14d;
             14'h2bd8 	:	val_out <= 16'he150;
             14'h2bd9 	:	val_out <= 16'he153;
             14'h2bda 	:	val_out <= 16'he156;
             14'h2bdb 	:	val_out <= 16'he159;
             14'h2bdc 	:	val_out <= 16'he15c;
             14'h2bdd 	:	val_out <= 16'he15f;
             14'h2bde 	:	val_out <= 16'he162;
             14'h2bdf 	:	val_out <= 16'he165;
             14'h2be0 	:	val_out <= 16'he168;
             14'h2be1 	:	val_out <= 16'he16b;
             14'h2be2 	:	val_out <= 16'he16d;
             14'h2be3 	:	val_out <= 16'he170;
             14'h2be4 	:	val_out <= 16'he173;
             14'h2be5 	:	val_out <= 16'he176;
             14'h2be6 	:	val_out <= 16'he179;
             14'h2be7 	:	val_out <= 16'he17c;
             14'h2be8 	:	val_out <= 16'he17f;
             14'h2be9 	:	val_out <= 16'he182;
             14'h2bea 	:	val_out <= 16'he185;
             14'h2beb 	:	val_out <= 16'he188;
             14'h2bec 	:	val_out <= 16'he18b;
             14'h2bed 	:	val_out <= 16'he18e;
             14'h2bee 	:	val_out <= 16'he191;
             14'h2bef 	:	val_out <= 16'he194;
             14'h2bf0 	:	val_out <= 16'he197;
             14'h2bf1 	:	val_out <= 16'he19a;
             14'h2bf2 	:	val_out <= 16'he19d;
             14'h2bf3 	:	val_out <= 16'he1a0;
             14'h2bf4 	:	val_out <= 16'he1a3;
             14'h2bf5 	:	val_out <= 16'he1a6;
             14'h2bf6 	:	val_out <= 16'he1a9;
             14'h2bf7 	:	val_out <= 16'he1ac;
             14'h2bf8 	:	val_out <= 16'he1af;
             14'h2bf9 	:	val_out <= 16'he1b2;
             14'h2bfa 	:	val_out <= 16'he1b5;
             14'h2bfb 	:	val_out <= 16'he1b8;
             14'h2bfc 	:	val_out <= 16'he1bb;
             14'h2bfd 	:	val_out <= 16'he1be;
             14'h2bfe 	:	val_out <= 16'he1c1;
             14'h2bff 	:	val_out <= 16'he1c4;
             14'h2c00 	:	val_out <= 16'he1c7;
             14'h2c01 	:	val_out <= 16'he1ca;
             14'h2c02 	:	val_out <= 16'he1cc;
             14'h2c03 	:	val_out <= 16'he1cf;
             14'h2c04 	:	val_out <= 16'he1d2;
             14'h2c05 	:	val_out <= 16'he1d5;
             14'h2c06 	:	val_out <= 16'he1d8;
             14'h2c07 	:	val_out <= 16'he1db;
             14'h2c08 	:	val_out <= 16'he1de;
             14'h2c09 	:	val_out <= 16'he1e1;
             14'h2c0a 	:	val_out <= 16'he1e4;
             14'h2c0b 	:	val_out <= 16'he1e7;
             14'h2c0c 	:	val_out <= 16'he1ea;
             14'h2c0d 	:	val_out <= 16'he1ed;
             14'h2c0e 	:	val_out <= 16'he1f0;
             14'h2c0f 	:	val_out <= 16'he1f3;
             14'h2c10 	:	val_out <= 16'he1f6;
             14'h2c11 	:	val_out <= 16'he1f9;
             14'h2c12 	:	val_out <= 16'he1fc;
             14'h2c13 	:	val_out <= 16'he1ff;
             14'h2c14 	:	val_out <= 16'he202;
             14'h2c15 	:	val_out <= 16'he205;
             14'h2c16 	:	val_out <= 16'he208;
             14'h2c17 	:	val_out <= 16'he20b;
             14'h2c18 	:	val_out <= 16'he20d;
             14'h2c19 	:	val_out <= 16'he210;
             14'h2c1a 	:	val_out <= 16'he213;
             14'h2c1b 	:	val_out <= 16'he216;
             14'h2c1c 	:	val_out <= 16'he219;
             14'h2c1d 	:	val_out <= 16'he21c;
             14'h2c1e 	:	val_out <= 16'he21f;
             14'h2c1f 	:	val_out <= 16'he222;
             14'h2c20 	:	val_out <= 16'he225;
             14'h2c21 	:	val_out <= 16'he228;
             14'h2c22 	:	val_out <= 16'he22b;
             14'h2c23 	:	val_out <= 16'he22e;
             14'h2c24 	:	val_out <= 16'he231;
             14'h2c25 	:	val_out <= 16'he234;
             14'h2c26 	:	val_out <= 16'he237;
             14'h2c27 	:	val_out <= 16'he23a;
             14'h2c28 	:	val_out <= 16'he23d;
             14'h2c29 	:	val_out <= 16'he240;
             14'h2c2a 	:	val_out <= 16'he242;
             14'h2c2b 	:	val_out <= 16'he245;
             14'h2c2c 	:	val_out <= 16'he248;
             14'h2c2d 	:	val_out <= 16'he24b;
             14'h2c2e 	:	val_out <= 16'he24e;
             14'h2c2f 	:	val_out <= 16'he251;
             14'h2c30 	:	val_out <= 16'he254;
             14'h2c31 	:	val_out <= 16'he257;
             14'h2c32 	:	val_out <= 16'he25a;
             14'h2c33 	:	val_out <= 16'he25d;
             14'h2c34 	:	val_out <= 16'he260;
             14'h2c35 	:	val_out <= 16'he263;
             14'h2c36 	:	val_out <= 16'he266;
             14'h2c37 	:	val_out <= 16'he269;
             14'h2c38 	:	val_out <= 16'he26c;
             14'h2c39 	:	val_out <= 16'he26f;
             14'h2c3a 	:	val_out <= 16'he271;
             14'h2c3b 	:	val_out <= 16'he274;
             14'h2c3c 	:	val_out <= 16'he277;
             14'h2c3d 	:	val_out <= 16'he27a;
             14'h2c3e 	:	val_out <= 16'he27d;
             14'h2c3f 	:	val_out <= 16'he280;
             14'h2c40 	:	val_out <= 16'he283;
             14'h2c41 	:	val_out <= 16'he286;
             14'h2c42 	:	val_out <= 16'he289;
             14'h2c43 	:	val_out <= 16'he28c;
             14'h2c44 	:	val_out <= 16'he28f;
             14'h2c45 	:	val_out <= 16'he292;
             14'h2c46 	:	val_out <= 16'he295;
             14'h2c47 	:	val_out <= 16'he298;
             14'h2c48 	:	val_out <= 16'he29a;
             14'h2c49 	:	val_out <= 16'he29d;
             14'h2c4a 	:	val_out <= 16'he2a0;
             14'h2c4b 	:	val_out <= 16'he2a3;
             14'h2c4c 	:	val_out <= 16'he2a6;
             14'h2c4d 	:	val_out <= 16'he2a9;
             14'h2c4e 	:	val_out <= 16'he2ac;
             14'h2c4f 	:	val_out <= 16'he2af;
             14'h2c50 	:	val_out <= 16'he2b2;
             14'h2c51 	:	val_out <= 16'he2b5;
             14'h2c52 	:	val_out <= 16'he2b8;
             14'h2c53 	:	val_out <= 16'he2bb;
             14'h2c54 	:	val_out <= 16'he2bd;
             14'h2c55 	:	val_out <= 16'he2c0;
             14'h2c56 	:	val_out <= 16'he2c3;
             14'h2c57 	:	val_out <= 16'he2c6;
             14'h2c58 	:	val_out <= 16'he2c9;
             14'h2c59 	:	val_out <= 16'he2cc;
             14'h2c5a 	:	val_out <= 16'he2cf;
             14'h2c5b 	:	val_out <= 16'he2d2;
             14'h2c5c 	:	val_out <= 16'he2d5;
             14'h2c5d 	:	val_out <= 16'he2d8;
             14'h2c5e 	:	val_out <= 16'he2db;
             14'h2c5f 	:	val_out <= 16'he2de;
             14'h2c60 	:	val_out <= 16'he2e0;
             14'h2c61 	:	val_out <= 16'he2e3;
             14'h2c62 	:	val_out <= 16'he2e6;
             14'h2c63 	:	val_out <= 16'he2e9;
             14'h2c64 	:	val_out <= 16'he2ec;
             14'h2c65 	:	val_out <= 16'he2ef;
             14'h2c66 	:	val_out <= 16'he2f2;
             14'h2c67 	:	val_out <= 16'he2f5;
             14'h2c68 	:	val_out <= 16'he2f8;
             14'h2c69 	:	val_out <= 16'he2fb;
             14'h2c6a 	:	val_out <= 16'he2fe;
             14'h2c6b 	:	val_out <= 16'he300;
             14'h2c6c 	:	val_out <= 16'he303;
             14'h2c6d 	:	val_out <= 16'he306;
             14'h2c6e 	:	val_out <= 16'he309;
             14'h2c6f 	:	val_out <= 16'he30c;
             14'h2c70 	:	val_out <= 16'he30f;
             14'h2c71 	:	val_out <= 16'he312;
             14'h2c72 	:	val_out <= 16'he315;
             14'h2c73 	:	val_out <= 16'he318;
             14'h2c74 	:	val_out <= 16'he31b;
             14'h2c75 	:	val_out <= 16'he31d;
             14'h2c76 	:	val_out <= 16'he320;
             14'h2c77 	:	val_out <= 16'he323;
             14'h2c78 	:	val_out <= 16'he326;
             14'h2c79 	:	val_out <= 16'he329;
             14'h2c7a 	:	val_out <= 16'he32c;
             14'h2c7b 	:	val_out <= 16'he32f;
             14'h2c7c 	:	val_out <= 16'he332;
             14'h2c7d 	:	val_out <= 16'he335;
             14'h2c7e 	:	val_out <= 16'he338;
             14'h2c7f 	:	val_out <= 16'he33a;
             14'h2c80 	:	val_out <= 16'he33d;
             14'h2c81 	:	val_out <= 16'he340;
             14'h2c82 	:	val_out <= 16'he343;
             14'h2c83 	:	val_out <= 16'he346;
             14'h2c84 	:	val_out <= 16'he349;
             14'h2c85 	:	val_out <= 16'he34c;
             14'h2c86 	:	val_out <= 16'he34f;
             14'h2c87 	:	val_out <= 16'he352;
             14'h2c88 	:	val_out <= 16'he354;
             14'h2c89 	:	val_out <= 16'he357;
             14'h2c8a 	:	val_out <= 16'he35a;
             14'h2c8b 	:	val_out <= 16'he35d;
             14'h2c8c 	:	val_out <= 16'he360;
             14'h2c8d 	:	val_out <= 16'he363;
             14'h2c8e 	:	val_out <= 16'he366;
             14'h2c8f 	:	val_out <= 16'he369;
             14'h2c90 	:	val_out <= 16'he36c;
             14'h2c91 	:	val_out <= 16'he36e;
             14'h2c92 	:	val_out <= 16'he371;
             14'h2c93 	:	val_out <= 16'he374;
             14'h2c94 	:	val_out <= 16'he377;
             14'h2c95 	:	val_out <= 16'he37a;
             14'h2c96 	:	val_out <= 16'he37d;
             14'h2c97 	:	val_out <= 16'he380;
             14'h2c98 	:	val_out <= 16'he383;
             14'h2c99 	:	val_out <= 16'he385;
             14'h2c9a 	:	val_out <= 16'he388;
             14'h2c9b 	:	val_out <= 16'he38b;
             14'h2c9c 	:	val_out <= 16'he38e;
             14'h2c9d 	:	val_out <= 16'he391;
             14'h2c9e 	:	val_out <= 16'he394;
             14'h2c9f 	:	val_out <= 16'he397;
             14'h2ca0 	:	val_out <= 16'he39a;
             14'h2ca1 	:	val_out <= 16'he39c;
             14'h2ca2 	:	val_out <= 16'he39f;
             14'h2ca3 	:	val_out <= 16'he3a2;
             14'h2ca4 	:	val_out <= 16'he3a5;
             14'h2ca5 	:	val_out <= 16'he3a8;
             14'h2ca6 	:	val_out <= 16'he3ab;
             14'h2ca7 	:	val_out <= 16'he3ae;
             14'h2ca8 	:	val_out <= 16'he3b1;
             14'h2ca9 	:	val_out <= 16'he3b3;
             14'h2caa 	:	val_out <= 16'he3b6;
             14'h2cab 	:	val_out <= 16'he3b9;
             14'h2cac 	:	val_out <= 16'he3bc;
             14'h2cad 	:	val_out <= 16'he3bf;
             14'h2cae 	:	val_out <= 16'he3c2;
             14'h2caf 	:	val_out <= 16'he3c5;
             14'h2cb0 	:	val_out <= 16'he3c8;
             14'h2cb1 	:	val_out <= 16'he3ca;
             14'h2cb2 	:	val_out <= 16'he3cd;
             14'h2cb3 	:	val_out <= 16'he3d0;
             14'h2cb4 	:	val_out <= 16'he3d3;
             14'h2cb5 	:	val_out <= 16'he3d6;
             14'h2cb6 	:	val_out <= 16'he3d9;
             14'h2cb7 	:	val_out <= 16'he3dc;
             14'h2cb8 	:	val_out <= 16'he3de;
             14'h2cb9 	:	val_out <= 16'he3e1;
             14'h2cba 	:	val_out <= 16'he3e4;
             14'h2cbb 	:	val_out <= 16'he3e7;
             14'h2cbc 	:	val_out <= 16'he3ea;
             14'h2cbd 	:	val_out <= 16'he3ed;
             14'h2cbe 	:	val_out <= 16'he3f0;
             14'h2cbf 	:	val_out <= 16'he3f3;
             14'h2cc0 	:	val_out <= 16'he3f5;
             14'h2cc1 	:	val_out <= 16'he3f8;
             14'h2cc2 	:	val_out <= 16'he3fb;
             14'h2cc3 	:	val_out <= 16'he3fe;
             14'h2cc4 	:	val_out <= 16'he401;
             14'h2cc5 	:	val_out <= 16'he404;
             14'h2cc6 	:	val_out <= 16'he407;
             14'h2cc7 	:	val_out <= 16'he409;
             14'h2cc8 	:	val_out <= 16'he40c;
             14'h2cc9 	:	val_out <= 16'he40f;
             14'h2cca 	:	val_out <= 16'he412;
             14'h2ccb 	:	val_out <= 16'he415;
             14'h2ccc 	:	val_out <= 16'he418;
             14'h2ccd 	:	val_out <= 16'he41b;
             14'h2cce 	:	val_out <= 16'he41d;
             14'h2ccf 	:	val_out <= 16'he420;
             14'h2cd0 	:	val_out <= 16'he423;
             14'h2cd1 	:	val_out <= 16'he426;
             14'h2cd2 	:	val_out <= 16'he429;
             14'h2cd3 	:	val_out <= 16'he42c;
             14'h2cd4 	:	val_out <= 16'he42e;
             14'h2cd5 	:	val_out <= 16'he431;
             14'h2cd6 	:	val_out <= 16'he434;
             14'h2cd7 	:	val_out <= 16'he437;
             14'h2cd8 	:	val_out <= 16'he43a;
             14'h2cd9 	:	val_out <= 16'he43d;
             14'h2cda 	:	val_out <= 16'he440;
             14'h2cdb 	:	val_out <= 16'he442;
             14'h2cdc 	:	val_out <= 16'he445;
             14'h2cdd 	:	val_out <= 16'he448;
             14'h2cde 	:	val_out <= 16'he44b;
             14'h2cdf 	:	val_out <= 16'he44e;
             14'h2ce0 	:	val_out <= 16'he451;
             14'h2ce1 	:	val_out <= 16'he453;
             14'h2ce2 	:	val_out <= 16'he456;
             14'h2ce3 	:	val_out <= 16'he459;
             14'h2ce4 	:	val_out <= 16'he45c;
             14'h2ce5 	:	val_out <= 16'he45f;
             14'h2ce6 	:	val_out <= 16'he462;
             14'h2ce7 	:	val_out <= 16'he464;
             14'h2ce8 	:	val_out <= 16'he467;
             14'h2ce9 	:	val_out <= 16'he46a;
             14'h2cea 	:	val_out <= 16'he46d;
             14'h2ceb 	:	val_out <= 16'he470;
             14'h2cec 	:	val_out <= 16'he473;
             14'h2ced 	:	val_out <= 16'he475;
             14'h2cee 	:	val_out <= 16'he478;
             14'h2cef 	:	val_out <= 16'he47b;
             14'h2cf0 	:	val_out <= 16'he47e;
             14'h2cf1 	:	val_out <= 16'he481;
             14'h2cf2 	:	val_out <= 16'he484;
             14'h2cf3 	:	val_out <= 16'he486;
             14'h2cf4 	:	val_out <= 16'he489;
             14'h2cf5 	:	val_out <= 16'he48c;
             14'h2cf6 	:	val_out <= 16'he48f;
             14'h2cf7 	:	val_out <= 16'he492;
             14'h2cf8 	:	val_out <= 16'he495;
             14'h2cf9 	:	val_out <= 16'he497;
             14'h2cfa 	:	val_out <= 16'he49a;
             14'h2cfb 	:	val_out <= 16'he49d;
             14'h2cfc 	:	val_out <= 16'he4a0;
             14'h2cfd 	:	val_out <= 16'he4a3;
             14'h2cfe 	:	val_out <= 16'he4a6;
             14'h2cff 	:	val_out <= 16'he4a8;
             14'h2d00 	:	val_out <= 16'he4ab;
             14'h2d01 	:	val_out <= 16'he4ae;
             14'h2d02 	:	val_out <= 16'he4b1;
             14'h2d03 	:	val_out <= 16'he4b4;
             14'h2d04 	:	val_out <= 16'he4b7;
             14'h2d05 	:	val_out <= 16'he4b9;
             14'h2d06 	:	val_out <= 16'he4bc;
             14'h2d07 	:	val_out <= 16'he4bf;
             14'h2d08 	:	val_out <= 16'he4c2;
             14'h2d09 	:	val_out <= 16'he4c5;
             14'h2d0a 	:	val_out <= 16'he4c7;
             14'h2d0b 	:	val_out <= 16'he4ca;
             14'h2d0c 	:	val_out <= 16'he4cd;
             14'h2d0d 	:	val_out <= 16'he4d0;
             14'h2d0e 	:	val_out <= 16'he4d3;
             14'h2d0f 	:	val_out <= 16'he4d6;
             14'h2d10 	:	val_out <= 16'he4d8;
             14'h2d11 	:	val_out <= 16'he4db;
             14'h2d12 	:	val_out <= 16'he4de;
             14'h2d13 	:	val_out <= 16'he4e1;
             14'h2d14 	:	val_out <= 16'he4e4;
             14'h2d15 	:	val_out <= 16'he4e6;
             14'h2d16 	:	val_out <= 16'he4e9;
             14'h2d17 	:	val_out <= 16'he4ec;
             14'h2d18 	:	val_out <= 16'he4ef;
             14'h2d19 	:	val_out <= 16'he4f2;
             14'h2d1a 	:	val_out <= 16'he4f5;
             14'h2d1b 	:	val_out <= 16'he4f7;
             14'h2d1c 	:	val_out <= 16'he4fa;
             14'h2d1d 	:	val_out <= 16'he4fd;
             14'h2d1e 	:	val_out <= 16'he500;
             14'h2d1f 	:	val_out <= 16'he503;
             14'h2d20 	:	val_out <= 16'he505;
             14'h2d21 	:	val_out <= 16'he508;
             14'h2d22 	:	val_out <= 16'he50b;
             14'h2d23 	:	val_out <= 16'he50e;
             14'h2d24 	:	val_out <= 16'he511;
             14'h2d25 	:	val_out <= 16'he513;
             14'h2d26 	:	val_out <= 16'he516;
             14'h2d27 	:	val_out <= 16'he519;
             14'h2d28 	:	val_out <= 16'he51c;
             14'h2d29 	:	val_out <= 16'he51f;
             14'h2d2a 	:	val_out <= 16'he521;
             14'h2d2b 	:	val_out <= 16'he524;
             14'h2d2c 	:	val_out <= 16'he527;
             14'h2d2d 	:	val_out <= 16'he52a;
             14'h2d2e 	:	val_out <= 16'he52d;
             14'h2d2f 	:	val_out <= 16'he52f;
             14'h2d30 	:	val_out <= 16'he532;
             14'h2d31 	:	val_out <= 16'he535;
             14'h2d32 	:	val_out <= 16'he538;
             14'h2d33 	:	val_out <= 16'he53b;
             14'h2d34 	:	val_out <= 16'he53d;
             14'h2d35 	:	val_out <= 16'he540;
             14'h2d36 	:	val_out <= 16'he543;
             14'h2d37 	:	val_out <= 16'he546;
             14'h2d38 	:	val_out <= 16'he549;
             14'h2d39 	:	val_out <= 16'he54b;
             14'h2d3a 	:	val_out <= 16'he54e;
             14'h2d3b 	:	val_out <= 16'he551;
             14'h2d3c 	:	val_out <= 16'he554;
             14'h2d3d 	:	val_out <= 16'he557;
             14'h2d3e 	:	val_out <= 16'he559;
             14'h2d3f 	:	val_out <= 16'he55c;
             14'h2d40 	:	val_out <= 16'he55f;
             14'h2d41 	:	val_out <= 16'he562;
             14'h2d42 	:	val_out <= 16'he565;
             14'h2d43 	:	val_out <= 16'he567;
             14'h2d44 	:	val_out <= 16'he56a;
             14'h2d45 	:	val_out <= 16'he56d;
             14'h2d46 	:	val_out <= 16'he570;
             14'h2d47 	:	val_out <= 16'he572;
             14'h2d48 	:	val_out <= 16'he575;
             14'h2d49 	:	val_out <= 16'he578;
             14'h2d4a 	:	val_out <= 16'he57b;
             14'h2d4b 	:	val_out <= 16'he57e;
             14'h2d4c 	:	val_out <= 16'he580;
             14'h2d4d 	:	val_out <= 16'he583;
             14'h2d4e 	:	val_out <= 16'he586;
             14'h2d4f 	:	val_out <= 16'he589;
             14'h2d50 	:	val_out <= 16'he58c;
             14'h2d51 	:	val_out <= 16'he58e;
             14'h2d52 	:	val_out <= 16'he591;
             14'h2d53 	:	val_out <= 16'he594;
             14'h2d54 	:	val_out <= 16'he597;
             14'h2d55 	:	val_out <= 16'he599;
             14'h2d56 	:	val_out <= 16'he59c;
             14'h2d57 	:	val_out <= 16'he59f;
             14'h2d58 	:	val_out <= 16'he5a2;
             14'h2d59 	:	val_out <= 16'he5a5;
             14'h2d5a 	:	val_out <= 16'he5a7;
             14'h2d5b 	:	val_out <= 16'he5aa;
             14'h2d5c 	:	val_out <= 16'he5ad;
             14'h2d5d 	:	val_out <= 16'he5b0;
             14'h2d5e 	:	val_out <= 16'he5b2;
             14'h2d5f 	:	val_out <= 16'he5b5;
             14'h2d60 	:	val_out <= 16'he5b8;
             14'h2d61 	:	val_out <= 16'he5bb;
             14'h2d62 	:	val_out <= 16'he5bd;
             14'h2d63 	:	val_out <= 16'he5c0;
             14'h2d64 	:	val_out <= 16'he5c3;
             14'h2d65 	:	val_out <= 16'he5c6;
             14'h2d66 	:	val_out <= 16'he5c9;
             14'h2d67 	:	val_out <= 16'he5cb;
             14'h2d68 	:	val_out <= 16'he5ce;
             14'h2d69 	:	val_out <= 16'he5d1;
             14'h2d6a 	:	val_out <= 16'he5d4;
             14'h2d6b 	:	val_out <= 16'he5d6;
             14'h2d6c 	:	val_out <= 16'he5d9;
             14'h2d6d 	:	val_out <= 16'he5dc;
             14'h2d6e 	:	val_out <= 16'he5df;
             14'h2d6f 	:	val_out <= 16'he5e1;
             14'h2d70 	:	val_out <= 16'he5e4;
             14'h2d71 	:	val_out <= 16'he5e7;
             14'h2d72 	:	val_out <= 16'he5ea;
             14'h2d73 	:	val_out <= 16'he5ed;
             14'h2d74 	:	val_out <= 16'he5ef;
             14'h2d75 	:	val_out <= 16'he5f2;
             14'h2d76 	:	val_out <= 16'he5f5;
             14'h2d77 	:	val_out <= 16'he5f8;
             14'h2d78 	:	val_out <= 16'he5fa;
             14'h2d79 	:	val_out <= 16'he5fd;
             14'h2d7a 	:	val_out <= 16'he600;
             14'h2d7b 	:	val_out <= 16'he603;
             14'h2d7c 	:	val_out <= 16'he605;
             14'h2d7d 	:	val_out <= 16'he608;
             14'h2d7e 	:	val_out <= 16'he60b;
             14'h2d7f 	:	val_out <= 16'he60e;
             14'h2d80 	:	val_out <= 16'he610;
             14'h2d81 	:	val_out <= 16'he613;
             14'h2d82 	:	val_out <= 16'he616;
             14'h2d83 	:	val_out <= 16'he619;
             14'h2d84 	:	val_out <= 16'he61b;
             14'h2d85 	:	val_out <= 16'he61e;
             14'h2d86 	:	val_out <= 16'he621;
             14'h2d87 	:	val_out <= 16'he624;
             14'h2d88 	:	val_out <= 16'he626;
             14'h2d89 	:	val_out <= 16'he629;
             14'h2d8a 	:	val_out <= 16'he62c;
             14'h2d8b 	:	val_out <= 16'he62f;
             14'h2d8c 	:	val_out <= 16'he631;
             14'h2d8d 	:	val_out <= 16'he634;
             14'h2d8e 	:	val_out <= 16'he637;
             14'h2d8f 	:	val_out <= 16'he63a;
             14'h2d90 	:	val_out <= 16'he63c;
             14'h2d91 	:	val_out <= 16'he63f;
             14'h2d92 	:	val_out <= 16'he642;
             14'h2d93 	:	val_out <= 16'he645;
             14'h2d94 	:	val_out <= 16'he647;
             14'h2d95 	:	val_out <= 16'he64a;
             14'h2d96 	:	val_out <= 16'he64d;
             14'h2d97 	:	val_out <= 16'he650;
             14'h2d98 	:	val_out <= 16'he652;
             14'h2d99 	:	val_out <= 16'he655;
             14'h2d9a 	:	val_out <= 16'he658;
             14'h2d9b 	:	val_out <= 16'he65b;
             14'h2d9c 	:	val_out <= 16'he65d;
             14'h2d9d 	:	val_out <= 16'he660;
             14'h2d9e 	:	val_out <= 16'he663;
             14'h2d9f 	:	val_out <= 16'he666;
             14'h2da0 	:	val_out <= 16'he668;
             14'h2da1 	:	val_out <= 16'he66b;
             14'h2da2 	:	val_out <= 16'he66e;
             14'h2da3 	:	val_out <= 16'he671;
             14'h2da4 	:	val_out <= 16'he673;
             14'h2da5 	:	val_out <= 16'he676;
             14'h2da6 	:	val_out <= 16'he679;
             14'h2da7 	:	val_out <= 16'he67b;
             14'h2da8 	:	val_out <= 16'he67e;
             14'h2da9 	:	val_out <= 16'he681;
             14'h2daa 	:	val_out <= 16'he684;
             14'h2dab 	:	val_out <= 16'he686;
             14'h2dac 	:	val_out <= 16'he689;
             14'h2dad 	:	val_out <= 16'he68c;
             14'h2dae 	:	val_out <= 16'he68f;
             14'h2daf 	:	val_out <= 16'he691;
             14'h2db0 	:	val_out <= 16'he694;
             14'h2db1 	:	val_out <= 16'he697;
             14'h2db2 	:	val_out <= 16'he69a;
             14'h2db3 	:	val_out <= 16'he69c;
             14'h2db4 	:	val_out <= 16'he69f;
             14'h2db5 	:	val_out <= 16'he6a2;
             14'h2db6 	:	val_out <= 16'he6a4;
             14'h2db7 	:	val_out <= 16'he6a7;
             14'h2db8 	:	val_out <= 16'he6aa;
             14'h2db9 	:	val_out <= 16'he6ad;
             14'h2dba 	:	val_out <= 16'he6af;
             14'h2dbb 	:	val_out <= 16'he6b2;
             14'h2dbc 	:	val_out <= 16'he6b5;
             14'h2dbd 	:	val_out <= 16'he6b7;
             14'h2dbe 	:	val_out <= 16'he6ba;
             14'h2dbf 	:	val_out <= 16'he6bd;
             14'h2dc0 	:	val_out <= 16'he6c0;
             14'h2dc1 	:	val_out <= 16'he6c2;
             14'h2dc2 	:	val_out <= 16'he6c5;
             14'h2dc3 	:	val_out <= 16'he6c8;
             14'h2dc4 	:	val_out <= 16'he6cb;
             14'h2dc5 	:	val_out <= 16'he6cd;
             14'h2dc6 	:	val_out <= 16'he6d0;
             14'h2dc7 	:	val_out <= 16'he6d3;
             14'h2dc8 	:	val_out <= 16'he6d5;
             14'h2dc9 	:	val_out <= 16'he6d8;
             14'h2dca 	:	val_out <= 16'he6db;
             14'h2dcb 	:	val_out <= 16'he6de;
             14'h2dcc 	:	val_out <= 16'he6e0;
             14'h2dcd 	:	val_out <= 16'he6e3;
             14'h2dce 	:	val_out <= 16'he6e6;
             14'h2dcf 	:	val_out <= 16'he6e8;
             14'h2dd0 	:	val_out <= 16'he6eb;
             14'h2dd1 	:	val_out <= 16'he6ee;
             14'h2dd2 	:	val_out <= 16'he6f1;
             14'h2dd3 	:	val_out <= 16'he6f3;
             14'h2dd4 	:	val_out <= 16'he6f6;
             14'h2dd5 	:	val_out <= 16'he6f9;
             14'h2dd6 	:	val_out <= 16'he6fb;
             14'h2dd7 	:	val_out <= 16'he6fe;
             14'h2dd8 	:	val_out <= 16'he701;
             14'h2dd9 	:	val_out <= 16'he704;
             14'h2dda 	:	val_out <= 16'he706;
             14'h2ddb 	:	val_out <= 16'he709;
             14'h2ddc 	:	val_out <= 16'he70c;
             14'h2ddd 	:	val_out <= 16'he70e;
             14'h2dde 	:	val_out <= 16'he711;
             14'h2ddf 	:	val_out <= 16'he714;
             14'h2de0 	:	val_out <= 16'he716;
             14'h2de1 	:	val_out <= 16'he719;
             14'h2de2 	:	val_out <= 16'he71c;
             14'h2de3 	:	val_out <= 16'he71f;
             14'h2de4 	:	val_out <= 16'he721;
             14'h2de5 	:	val_out <= 16'he724;
             14'h2de6 	:	val_out <= 16'he727;
             14'h2de7 	:	val_out <= 16'he729;
             14'h2de8 	:	val_out <= 16'he72c;
             14'h2de9 	:	val_out <= 16'he72f;
             14'h2dea 	:	val_out <= 16'he731;
             14'h2deb 	:	val_out <= 16'he734;
             14'h2dec 	:	val_out <= 16'he737;
             14'h2ded 	:	val_out <= 16'he73a;
             14'h2dee 	:	val_out <= 16'he73c;
             14'h2def 	:	val_out <= 16'he73f;
             14'h2df0 	:	val_out <= 16'he742;
             14'h2df1 	:	val_out <= 16'he744;
             14'h2df2 	:	val_out <= 16'he747;
             14'h2df3 	:	val_out <= 16'he74a;
             14'h2df4 	:	val_out <= 16'he74c;
             14'h2df5 	:	val_out <= 16'he74f;
             14'h2df6 	:	val_out <= 16'he752;
             14'h2df7 	:	val_out <= 16'he754;
             14'h2df8 	:	val_out <= 16'he757;
             14'h2df9 	:	val_out <= 16'he75a;
             14'h2dfa 	:	val_out <= 16'he75d;
             14'h2dfb 	:	val_out <= 16'he75f;
             14'h2dfc 	:	val_out <= 16'he762;
             14'h2dfd 	:	val_out <= 16'he765;
             14'h2dfe 	:	val_out <= 16'he767;
             14'h2dff 	:	val_out <= 16'he76a;
             14'h2e00 	:	val_out <= 16'he76d;
             14'h2e01 	:	val_out <= 16'he76f;
             14'h2e02 	:	val_out <= 16'he772;
             14'h2e03 	:	val_out <= 16'he775;
             14'h2e04 	:	val_out <= 16'he777;
             14'h2e05 	:	val_out <= 16'he77a;
             14'h2e06 	:	val_out <= 16'he77d;
             14'h2e07 	:	val_out <= 16'he77f;
             14'h2e08 	:	val_out <= 16'he782;
             14'h2e09 	:	val_out <= 16'he785;
             14'h2e0a 	:	val_out <= 16'he788;
             14'h2e0b 	:	val_out <= 16'he78a;
             14'h2e0c 	:	val_out <= 16'he78d;
             14'h2e0d 	:	val_out <= 16'he790;
             14'h2e0e 	:	val_out <= 16'he792;
             14'h2e0f 	:	val_out <= 16'he795;
             14'h2e10 	:	val_out <= 16'he798;
             14'h2e11 	:	val_out <= 16'he79a;
             14'h2e12 	:	val_out <= 16'he79d;
             14'h2e13 	:	val_out <= 16'he7a0;
             14'h2e14 	:	val_out <= 16'he7a2;
             14'h2e15 	:	val_out <= 16'he7a5;
             14'h2e16 	:	val_out <= 16'he7a8;
             14'h2e17 	:	val_out <= 16'he7aa;
             14'h2e18 	:	val_out <= 16'he7ad;
             14'h2e19 	:	val_out <= 16'he7b0;
             14'h2e1a 	:	val_out <= 16'he7b2;
             14'h2e1b 	:	val_out <= 16'he7b5;
             14'h2e1c 	:	val_out <= 16'he7b8;
             14'h2e1d 	:	val_out <= 16'he7ba;
             14'h2e1e 	:	val_out <= 16'he7bd;
             14'h2e1f 	:	val_out <= 16'he7c0;
             14'h2e20 	:	val_out <= 16'he7c2;
             14'h2e21 	:	val_out <= 16'he7c5;
             14'h2e22 	:	val_out <= 16'he7c8;
             14'h2e23 	:	val_out <= 16'he7ca;
             14'h2e24 	:	val_out <= 16'he7cd;
             14'h2e25 	:	val_out <= 16'he7d0;
             14'h2e26 	:	val_out <= 16'he7d2;
             14'h2e27 	:	val_out <= 16'he7d5;
             14'h2e28 	:	val_out <= 16'he7d8;
             14'h2e29 	:	val_out <= 16'he7da;
             14'h2e2a 	:	val_out <= 16'he7dd;
             14'h2e2b 	:	val_out <= 16'he7e0;
             14'h2e2c 	:	val_out <= 16'he7e2;
             14'h2e2d 	:	val_out <= 16'he7e5;
             14'h2e2e 	:	val_out <= 16'he7e8;
             14'h2e2f 	:	val_out <= 16'he7ea;
             14'h2e30 	:	val_out <= 16'he7ed;
             14'h2e31 	:	val_out <= 16'he7f0;
             14'h2e32 	:	val_out <= 16'he7f2;
             14'h2e33 	:	val_out <= 16'he7f5;
             14'h2e34 	:	val_out <= 16'he7f8;
             14'h2e35 	:	val_out <= 16'he7fa;
             14'h2e36 	:	val_out <= 16'he7fd;
             14'h2e37 	:	val_out <= 16'he800;
             14'h2e38 	:	val_out <= 16'he802;
             14'h2e39 	:	val_out <= 16'he805;
             14'h2e3a 	:	val_out <= 16'he808;
             14'h2e3b 	:	val_out <= 16'he80a;
             14'h2e3c 	:	val_out <= 16'he80d;
             14'h2e3d 	:	val_out <= 16'he810;
             14'h2e3e 	:	val_out <= 16'he812;
             14'h2e3f 	:	val_out <= 16'he815;
             14'h2e40 	:	val_out <= 16'he817;
             14'h2e41 	:	val_out <= 16'he81a;
             14'h2e42 	:	val_out <= 16'he81d;
             14'h2e43 	:	val_out <= 16'he81f;
             14'h2e44 	:	val_out <= 16'he822;
             14'h2e45 	:	val_out <= 16'he825;
             14'h2e46 	:	val_out <= 16'he827;
             14'h2e47 	:	val_out <= 16'he82a;
             14'h2e48 	:	val_out <= 16'he82d;
             14'h2e49 	:	val_out <= 16'he82f;
             14'h2e4a 	:	val_out <= 16'he832;
             14'h2e4b 	:	val_out <= 16'he835;
             14'h2e4c 	:	val_out <= 16'he837;
             14'h2e4d 	:	val_out <= 16'he83a;
             14'h2e4e 	:	val_out <= 16'he83d;
             14'h2e4f 	:	val_out <= 16'he83f;
             14'h2e50 	:	val_out <= 16'he842;
             14'h2e51 	:	val_out <= 16'he844;
             14'h2e52 	:	val_out <= 16'he847;
             14'h2e53 	:	val_out <= 16'he84a;
             14'h2e54 	:	val_out <= 16'he84c;
             14'h2e55 	:	val_out <= 16'he84f;
             14'h2e56 	:	val_out <= 16'he852;
             14'h2e57 	:	val_out <= 16'he854;
             14'h2e58 	:	val_out <= 16'he857;
             14'h2e59 	:	val_out <= 16'he85a;
             14'h2e5a 	:	val_out <= 16'he85c;
             14'h2e5b 	:	val_out <= 16'he85f;
             14'h2e5c 	:	val_out <= 16'he862;
             14'h2e5d 	:	val_out <= 16'he864;
             14'h2e5e 	:	val_out <= 16'he867;
             14'h2e5f 	:	val_out <= 16'he869;
             14'h2e60 	:	val_out <= 16'he86c;
             14'h2e61 	:	val_out <= 16'he86f;
             14'h2e62 	:	val_out <= 16'he871;
             14'h2e63 	:	val_out <= 16'he874;
             14'h2e64 	:	val_out <= 16'he877;
             14'h2e65 	:	val_out <= 16'he879;
             14'h2e66 	:	val_out <= 16'he87c;
             14'h2e67 	:	val_out <= 16'he87e;
             14'h2e68 	:	val_out <= 16'he881;
             14'h2e69 	:	val_out <= 16'he884;
             14'h2e6a 	:	val_out <= 16'he886;
             14'h2e6b 	:	val_out <= 16'he889;
             14'h2e6c 	:	val_out <= 16'he88c;
             14'h2e6d 	:	val_out <= 16'he88e;
             14'h2e6e 	:	val_out <= 16'he891;
             14'h2e6f 	:	val_out <= 16'he893;
             14'h2e70 	:	val_out <= 16'he896;
             14'h2e71 	:	val_out <= 16'he899;
             14'h2e72 	:	val_out <= 16'he89b;
             14'h2e73 	:	val_out <= 16'he89e;
             14'h2e74 	:	val_out <= 16'he8a1;
             14'h2e75 	:	val_out <= 16'he8a3;
             14'h2e76 	:	val_out <= 16'he8a6;
             14'h2e77 	:	val_out <= 16'he8a8;
             14'h2e78 	:	val_out <= 16'he8ab;
             14'h2e79 	:	val_out <= 16'he8ae;
             14'h2e7a 	:	val_out <= 16'he8b0;
             14'h2e7b 	:	val_out <= 16'he8b3;
             14'h2e7c 	:	val_out <= 16'he8b6;
             14'h2e7d 	:	val_out <= 16'he8b8;
             14'h2e7e 	:	val_out <= 16'he8bb;
             14'h2e7f 	:	val_out <= 16'he8bd;
             14'h2e80 	:	val_out <= 16'he8c0;
             14'h2e81 	:	val_out <= 16'he8c3;
             14'h2e82 	:	val_out <= 16'he8c5;
             14'h2e83 	:	val_out <= 16'he8c8;
             14'h2e84 	:	val_out <= 16'he8cb;
             14'h2e85 	:	val_out <= 16'he8cd;
             14'h2e86 	:	val_out <= 16'he8d0;
             14'h2e87 	:	val_out <= 16'he8d2;
             14'h2e88 	:	val_out <= 16'he8d5;
             14'h2e89 	:	val_out <= 16'he8d8;
             14'h2e8a 	:	val_out <= 16'he8da;
             14'h2e8b 	:	val_out <= 16'he8dd;
             14'h2e8c 	:	val_out <= 16'he8df;
             14'h2e8d 	:	val_out <= 16'he8e2;
             14'h2e8e 	:	val_out <= 16'he8e5;
             14'h2e8f 	:	val_out <= 16'he8e7;
             14'h2e90 	:	val_out <= 16'he8ea;
             14'h2e91 	:	val_out <= 16'he8ec;
             14'h2e92 	:	val_out <= 16'he8ef;
             14'h2e93 	:	val_out <= 16'he8f2;
             14'h2e94 	:	val_out <= 16'he8f4;
             14'h2e95 	:	val_out <= 16'he8f7;
             14'h2e96 	:	val_out <= 16'he8f9;
             14'h2e97 	:	val_out <= 16'he8fc;
             14'h2e98 	:	val_out <= 16'he8ff;
             14'h2e99 	:	val_out <= 16'he901;
             14'h2e9a 	:	val_out <= 16'he904;
             14'h2e9b 	:	val_out <= 16'he906;
             14'h2e9c 	:	val_out <= 16'he909;
             14'h2e9d 	:	val_out <= 16'he90c;
             14'h2e9e 	:	val_out <= 16'he90e;
             14'h2e9f 	:	val_out <= 16'he911;
             14'h2ea0 	:	val_out <= 16'he913;
             14'h2ea1 	:	val_out <= 16'he916;
             14'h2ea2 	:	val_out <= 16'he919;
             14'h2ea3 	:	val_out <= 16'he91b;
             14'h2ea4 	:	val_out <= 16'he91e;
             14'h2ea5 	:	val_out <= 16'he920;
             14'h2ea6 	:	val_out <= 16'he923;
             14'h2ea7 	:	val_out <= 16'he926;
             14'h2ea8 	:	val_out <= 16'he928;
             14'h2ea9 	:	val_out <= 16'he92b;
             14'h2eaa 	:	val_out <= 16'he92d;
             14'h2eab 	:	val_out <= 16'he930;
             14'h2eac 	:	val_out <= 16'he933;
             14'h2ead 	:	val_out <= 16'he935;
             14'h2eae 	:	val_out <= 16'he938;
             14'h2eaf 	:	val_out <= 16'he93a;
             14'h2eb0 	:	val_out <= 16'he93d;
             14'h2eb1 	:	val_out <= 16'he940;
             14'h2eb2 	:	val_out <= 16'he942;
             14'h2eb3 	:	val_out <= 16'he945;
             14'h2eb4 	:	val_out <= 16'he947;
             14'h2eb5 	:	val_out <= 16'he94a;
             14'h2eb6 	:	val_out <= 16'he94d;
             14'h2eb7 	:	val_out <= 16'he94f;
             14'h2eb8 	:	val_out <= 16'he952;
             14'h2eb9 	:	val_out <= 16'he954;
             14'h2eba 	:	val_out <= 16'he957;
             14'h2ebb 	:	val_out <= 16'he959;
             14'h2ebc 	:	val_out <= 16'he95c;
             14'h2ebd 	:	val_out <= 16'he95f;
             14'h2ebe 	:	val_out <= 16'he961;
             14'h2ebf 	:	val_out <= 16'he964;
             14'h2ec0 	:	val_out <= 16'he966;
             14'h2ec1 	:	val_out <= 16'he969;
             14'h2ec2 	:	val_out <= 16'he96c;
             14'h2ec3 	:	val_out <= 16'he96e;
             14'h2ec4 	:	val_out <= 16'he971;
             14'h2ec5 	:	val_out <= 16'he973;
             14'h2ec6 	:	val_out <= 16'he976;
             14'h2ec7 	:	val_out <= 16'he978;
             14'h2ec8 	:	val_out <= 16'he97b;
             14'h2ec9 	:	val_out <= 16'he97e;
             14'h2eca 	:	val_out <= 16'he980;
             14'h2ecb 	:	val_out <= 16'he983;
             14'h2ecc 	:	val_out <= 16'he985;
             14'h2ecd 	:	val_out <= 16'he988;
             14'h2ece 	:	val_out <= 16'he98a;
             14'h2ecf 	:	val_out <= 16'he98d;
             14'h2ed0 	:	val_out <= 16'he990;
             14'h2ed1 	:	val_out <= 16'he992;
             14'h2ed2 	:	val_out <= 16'he995;
             14'h2ed3 	:	val_out <= 16'he997;
             14'h2ed4 	:	val_out <= 16'he99a;
             14'h2ed5 	:	val_out <= 16'he99c;
             14'h2ed6 	:	val_out <= 16'he99f;
             14'h2ed7 	:	val_out <= 16'he9a2;
             14'h2ed8 	:	val_out <= 16'he9a4;
             14'h2ed9 	:	val_out <= 16'he9a7;
             14'h2eda 	:	val_out <= 16'he9a9;
             14'h2edb 	:	val_out <= 16'he9ac;
             14'h2edc 	:	val_out <= 16'he9ae;
             14'h2edd 	:	val_out <= 16'he9b1;
             14'h2ede 	:	val_out <= 16'he9b4;
             14'h2edf 	:	val_out <= 16'he9b6;
             14'h2ee0 	:	val_out <= 16'he9b9;
             14'h2ee1 	:	val_out <= 16'he9bb;
             14'h2ee2 	:	val_out <= 16'he9be;
             14'h2ee3 	:	val_out <= 16'he9c0;
             14'h2ee4 	:	val_out <= 16'he9c3;
             14'h2ee5 	:	val_out <= 16'he9c5;
             14'h2ee6 	:	val_out <= 16'he9c8;
             14'h2ee7 	:	val_out <= 16'he9cb;
             14'h2ee8 	:	val_out <= 16'he9cd;
             14'h2ee9 	:	val_out <= 16'he9d0;
             14'h2eea 	:	val_out <= 16'he9d2;
             14'h2eeb 	:	val_out <= 16'he9d5;
             14'h2eec 	:	val_out <= 16'he9d7;
             14'h2eed 	:	val_out <= 16'he9da;
             14'h2eee 	:	val_out <= 16'he9dd;
             14'h2eef 	:	val_out <= 16'he9df;
             14'h2ef0 	:	val_out <= 16'he9e2;
             14'h2ef1 	:	val_out <= 16'he9e4;
             14'h2ef2 	:	val_out <= 16'he9e7;
             14'h2ef3 	:	val_out <= 16'he9e9;
             14'h2ef4 	:	val_out <= 16'he9ec;
             14'h2ef5 	:	val_out <= 16'he9ee;
             14'h2ef6 	:	val_out <= 16'he9f1;
             14'h2ef7 	:	val_out <= 16'he9f3;
             14'h2ef8 	:	val_out <= 16'he9f6;
             14'h2ef9 	:	val_out <= 16'he9f9;
             14'h2efa 	:	val_out <= 16'he9fb;
             14'h2efb 	:	val_out <= 16'he9fe;
             14'h2efc 	:	val_out <= 16'hea00;
             14'h2efd 	:	val_out <= 16'hea03;
             14'h2efe 	:	val_out <= 16'hea05;
             14'h2eff 	:	val_out <= 16'hea08;
             14'h2f00 	:	val_out <= 16'hea0a;
             14'h2f01 	:	val_out <= 16'hea0d;
             14'h2f02 	:	val_out <= 16'hea10;
             14'h2f03 	:	val_out <= 16'hea12;
             14'h2f04 	:	val_out <= 16'hea15;
             14'h2f05 	:	val_out <= 16'hea17;
             14'h2f06 	:	val_out <= 16'hea1a;
             14'h2f07 	:	val_out <= 16'hea1c;
             14'h2f08 	:	val_out <= 16'hea1f;
             14'h2f09 	:	val_out <= 16'hea21;
             14'h2f0a 	:	val_out <= 16'hea24;
             14'h2f0b 	:	val_out <= 16'hea26;
             14'h2f0c 	:	val_out <= 16'hea29;
             14'h2f0d 	:	val_out <= 16'hea2b;
             14'h2f0e 	:	val_out <= 16'hea2e;
             14'h2f0f 	:	val_out <= 16'hea31;
             14'h2f10 	:	val_out <= 16'hea33;
             14'h2f11 	:	val_out <= 16'hea36;
             14'h2f12 	:	val_out <= 16'hea38;
             14'h2f13 	:	val_out <= 16'hea3b;
             14'h2f14 	:	val_out <= 16'hea3d;
             14'h2f15 	:	val_out <= 16'hea40;
             14'h2f16 	:	val_out <= 16'hea42;
             14'h2f17 	:	val_out <= 16'hea45;
             14'h2f18 	:	val_out <= 16'hea47;
             14'h2f19 	:	val_out <= 16'hea4a;
             14'h2f1a 	:	val_out <= 16'hea4c;
             14'h2f1b 	:	val_out <= 16'hea4f;
             14'h2f1c 	:	val_out <= 16'hea51;
             14'h2f1d 	:	val_out <= 16'hea54;
             14'h2f1e 	:	val_out <= 16'hea57;
             14'h2f1f 	:	val_out <= 16'hea59;
             14'h2f20 	:	val_out <= 16'hea5c;
             14'h2f21 	:	val_out <= 16'hea5e;
             14'h2f22 	:	val_out <= 16'hea61;
             14'h2f23 	:	val_out <= 16'hea63;
             14'h2f24 	:	val_out <= 16'hea66;
             14'h2f25 	:	val_out <= 16'hea68;
             14'h2f26 	:	val_out <= 16'hea6b;
             14'h2f27 	:	val_out <= 16'hea6d;
             14'h2f28 	:	val_out <= 16'hea70;
             14'h2f29 	:	val_out <= 16'hea72;
             14'h2f2a 	:	val_out <= 16'hea75;
             14'h2f2b 	:	val_out <= 16'hea77;
             14'h2f2c 	:	val_out <= 16'hea7a;
             14'h2f2d 	:	val_out <= 16'hea7c;
             14'h2f2e 	:	val_out <= 16'hea7f;
             14'h2f2f 	:	val_out <= 16'hea81;
             14'h2f30 	:	val_out <= 16'hea84;
             14'h2f31 	:	val_out <= 16'hea87;
             14'h2f32 	:	val_out <= 16'hea89;
             14'h2f33 	:	val_out <= 16'hea8c;
             14'h2f34 	:	val_out <= 16'hea8e;
             14'h2f35 	:	val_out <= 16'hea91;
             14'h2f36 	:	val_out <= 16'hea93;
             14'h2f37 	:	val_out <= 16'hea96;
             14'h2f38 	:	val_out <= 16'hea98;
             14'h2f39 	:	val_out <= 16'hea9b;
             14'h2f3a 	:	val_out <= 16'hea9d;
             14'h2f3b 	:	val_out <= 16'heaa0;
             14'h2f3c 	:	val_out <= 16'heaa2;
             14'h2f3d 	:	val_out <= 16'heaa5;
             14'h2f3e 	:	val_out <= 16'heaa7;
             14'h2f3f 	:	val_out <= 16'heaaa;
             14'h2f40 	:	val_out <= 16'heaac;
             14'h2f41 	:	val_out <= 16'heaaf;
             14'h2f42 	:	val_out <= 16'heab1;
             14'h2f43 	:	val_out <= 16'heab4;
             14'h2f44 	:	val_out <= 16'heab6;
             14'h2f45 	:	val_out <= 16'heab9;
             14'h2f46 	:	val_out <= 16'heabb;
             14'h2f47 	:	val_out <= 16'heabe;
             14'h2f48 	:	val_out <= 16'heac0;
             14'h2f49 	:	val_out <= 16'heac3;
             14'h2f4a 	:	val_out <= 16'heac5;
             14'h2f4b 	:	val_out <= 16'heac8;
             14'h2f4c 	:	val_out <= 16'heaca;
             14'h2f4d 	:	val_out <= 16'heacd;
             14'h2f4e 	:	val_out <= 16'heacf;
             14'h2f4f 	:	val_out <= 16'head2;
             14'h2f50 	:	val_out <= 16'head4;
             14'h2f51 	:	val_out <= 16'head7;
             14'h2f52 	:	val_out <= 16'head9;
             14'h2f53 	:	val_out <= 16'headc;
             14'h2f54 	:	val_out <= 16'heade;
             14'h2f55 	:	val_out <= 16'heae1;
             14'h2f56 	:	val_out <= 16'heae3;
             14'h2f57 	:	val_out <= 16'heae6;
             14'h2f58 	:	val_out <= 16'heae8;
             14'h2f59 	:	val_out <= 16'heaeb;
             14'h2f5a 	:	val_out <= 16'heaed;
             14'h2f5b 	:	val_out <= 16'heaf0;
             14'h2f5c 	:	val_out <= 16'heaf2;
             14'h2f5d 	:	val_out <= 16'heaf5;
             14'h2f5e 	:	val_out <= 16'heaf7;
             14'h2f5f 	:	val_out <= 16'heafa;
             14'h2f60 	:	val_out <= 16'heafc;
             14'h2f61 	:	val_out <= 16'heaff;
             14'h2f62 	:	val_out <= 16'heb01;
             14'h2f63 	:	val_out <= 16'heb04;
             14'h2f64 	:	val_out <= 16'heb06;
             14'h2f65 	:	val_out <= 16'heb09;
             14'h2f66 	:	val_out <= 16'heb0b;
             14'h2f67 	:	val_out <= 16'heb0e;
             14'h2f68 	:	val_out <= 16'heb10;
             14'h2f69 	:	val_out <= 16'heb13;
             14'h2f6a 	:	val_out <= 16'heb15;
             14'h2f6b 	:	val_out <= 16'heb18;
             14'h2f6c 	:	val_out <= 16'heb1a;
             14'h2f6d 	:	val_out <= 16'heb1d;
             14'h2f6e 	:	val_out <= 16'heb1f;
             14'h2f6f 	:	val_out <= 16'heb22;
             14'h2f70 	:	val_out <= 16'heb24;
             14'h2f71 	:	val_out <= 16'heb27;
             14'h2f72 	:	val_out <= 16'heb29;
             14'h2f73 	:	val_out <= 16'heb2c;
             14'h2f74 	:	val_out <= 16'heb2e;
             14'h2f75 	:	val_out <= 16'heb31;
             14'h2f76 	:	val_out <= 16'heb33;
             14'h2f77 	:	val_out <= 16'heb35;
             14'h2f78 	:	val_out <= 16'heb38;
             14'h2f79 	:	val_out <= 16'heb3a;
             14'h2f7a 	:	val_out <= 16'heb3d;
             14'h2f7b 	:	val_out <= 16'heb3f;
             14'h2f7c 	:	val_out <= 16'heb42;
             14'h2f7d 	:	val_out <= 16'heb44;
             14'h2f7e 	:	val_out <= 16'heb47;
             14'h2f7f 	:	val_out <= 16'heb49;
             14'h2f80 	:	val_out <= 16'heb4c;
             14'h2f81 	:	val_out <= 16'heb4e;
             14'h2f82 	:	val_out <= 16'heb51;
             14'h2f83 	:	val_out <= 16'heb53;
             14'h2f84 	:	val_out <= 16'heb56;
             14'h2f85 	:	val_out <= 16'heb58;
             14'h2f86 	:	val_out <= 16'heb5b;
             14'h2f87 	:	val_out <= 16'heb5d;
             14'h2f88 	:	val_out <= 16'heb60;
             14'h2f89 	:	val_out <= 16'heb62;
             14'h2f8a 	:	val_out <= 16'heb65;
             14'h2f8b 	:	val_out <= 16'heb67;
             14'h2f8c 	:	val_out <= 16'heb69;
             14'h2f8d 	:	val_out <= 16'heb6c;
             14'h2f8e 	:	val_out <= 16'heb6e;
             14'h2f8f 	:	val_out <= 16'heb71;
             14'h2f90 	:	val_out <= 16'heb73;
             14'h2f91 	:	val_out <= 16'heb76;
             14'h2f92 	:	val_out <= 16'heb78;
             14'h2f93 	:	val_out <= 16'heb7b;
             14'h2f94 	:	val_out <= 16'heb7d;
             14'h2f95 	:	val_out <= 16'heb80;
             14'h2f96 	:	val_out <= 16'heb82;
             14'h2f97 	:	val_out <= 16'heb85;
             14'h2f98 	:	val_out <= 16'heb87;
             14'h2f99 	:	val_out <= 16'heb89;
             14'h2f9a 	:	val_out <= 16'heb8c;
             14'h2f9b 	:	val_out <= 16'heb8e;
             14'h2f9c 	:	val_out <= 16'heb91;
             14'h2f9d 	:	val_out <= 16'heb93;
             14'h2f9e 	:	val_out <= 16'heb96;
             14'h2f9f 	:	val_out <= 16'heb98;
             14'h2fa0 	:	val_out <= 16'heb9b;
             14'h2fa1 	:	val_out <= 16'heb9d;
             14'h2fa2 	:	val_out <= 16'heba0;
             14'h2fa3 	:	val_out <= 16'heba2;
             14'h2fa4 	:	val_out <= 16'heba5;
             14'h2fa5 	:	val_out <= 16'heba7;
             14'h2fa6 	:	val_out <= 16'heba9;
             14'h2fa7 	:	val_out <= 16'hebac;
             14'h2fa8 	:	val_out <= 16'hebae;
             14'h2fa9 	:	val_out <= 16'hebb1;
             14'h2faa 	:	val_out <= 16'hebb3;
             14'h2fab 	:	val_out <= 16'hebb6;
             14'h2fac 	:	val_out <= 16'hebb8;
             14'h2fad 	:	val_out <= 16'hebbb;
             14'h2fae 	:	val_out <= 16'hebbd;
             14'h2faf 	:	val_out <= 16'hebc0;
             14'h2fb0 	:	val_out <= 16'hebc2;
             14'h2fb1 	:	val_out <= 16'hebc4;
             14'h2fb2 	:	val_out <= 16'hebc7;
             14'h2fb3 	:	val_out <= 16'hebc9;
             14'h2fb4 	:	val_out <= 16'hebcc;
             14'h2fb5 	:	val_out <= 16'hebce;
             14'h2fb6 	:	val_out <= 16'hebd1;
             14'h2fb7 	:	val_out <= 16'hebd3;
             14'h2fb8 	:	val_out <= 16'hebd6;
             14'h2fb9 	:	val_out <= 16'hebd8;
             14'h2fba 	:	val_out <= 16'hebda;
             14'h2fbb 	:	val_out <= 16'hebdd;
             14'h2fbc 	:	val_out <= 16'hebdf;
             14'h2fbd 	:	val_out <= 16'hebe2;
             14'h2fbe 	:	val_out <= 16'hebe4;
             14'h2fbf 	:	val_out <= 16'hebe7;
             14'h2fc0 	:	val_out <= 16'hebe9;
             14'h2fc1 	:	val_out <= 16'hebec;
             14'h2fc2 	:	val_out <= 16'hebee;
             14'h2fc3 	:	val_out <= 16'hebf0;
             14'h2fc4 	:	val_out <= 16'hebf3;
             14'h2fc5 	:	val_out <= 16'hebf5;
             14'h2fc6 	:	val_out <= 16'hebf8;
             14'h2fc7 	:	val_out <= 16'hebfa;
             14'h2fc8 	:	val_out <= 16'hebfd;
             14'h2fc9 	:	val_out <= 16'hebff;
             14'h2fca 	:	val_out <= 16'hec01;
             14'h2fcb 	:	val_out <= 16'hec04;
             14'h2fcc 	:	val_out <= 16'hec06;
             14'h2fcd 	:	val_out <= 16'hec09;
             14'h2fce 	:	val_out <= 16'hec0b;
             14'h2fcf 	:	val_out <= 16'hec0e;
             14'h2fd0 	:	val_out <= 16'hec10;
             14'h2fd1 	:	val_out <= 16'hec12;
             14'h2fd2 	:	val_out <= 16'hec15;
             14'h2fd3 	:	val_out <= 16'hec17;
             14'h2fd4 	:	val_out <= 16'hec1a;
             14'h2fd5 	:	val_out <= 16'hec1c;
             14'h2fd6 	:	val_out <= 16'hec1f;
             14'h2fd7 	:	val_out <= 16'hec21;
             14'h2fd8 	:	val_out <= 16'hec23;
             14'h2fd9 	:	val_out <= 16'hec26;
             14'h2fda 	:	val_out <= 16'hec28;
             14'h2fdb 	:	val_out <= 16'hec2b;
             14'h2fdc 	:	val_out <= 16'hec2d;
             14'h2fdd 	:	val_out <= 16'hec30;
             14'h2fde 	:	val_out <= 16'hec32;
             14'h2fdf 	:	val_out <= 16'hec34;
             14'h2fe0 	:	val_out <= 16'hec37;
             14'h2fe1 	:	val_out <= 16'hec39;
             14'h2fe2 	:	val_out <= 16'hec3c;
             14'h2fe3 	:	val_out <= 16'hec3e;
             14'h2fe4 	:	val_out <= 16'hec41;
             14'h2fe5 	:	val_out <= 16'hec43;
             14'h2fe6 	:	val_out <= 16'hec45;
             14'h2fe7 	:	val_out <= 16'hec48;
             14'h2fe8 	:	val_out <= 16'hec4a;
             14'h2fe9 	:	val_out <= 16'hec4d;
             14'h2fea 	:	val_out <= 16'hec4f;
             14'h2feb 	:	val_out <= 16'hec51;
             14'h2fec 	:	val_out <= 16'hec54;
             14'h2fed 	:	val_out <= 16'hec56;
             14'h2fee 	:	val_out <= 16'hec59;
             14'h2fef 	:	val_out <= 16'hec5b;
             14'h2ff0 	:	val_out <= 16'hec5e;
             14'h2ff1 	:	val_out <= 16'hec60;
             14'h2ff2 	:	val_out <= 16'hec62;
             14'h2ff3 	:	val_out <= 16'hec65;
             14'h2ff4 	:	val_out <= 16'hec67;
             14'h2ff5 	:	val_out <= 16'hec6a;
             14'h2ff6 	:	val_out <= 16'hec6c;
             14'h2ff7 	:	val_out <= 16'hec6e;
             14'h2ff8 	:	val_out <= 16'hec71;
             14'h2ff9 	:	val_out <= 16'hec73;
             14'h2ffa 	:	val_out <= 16'hec76;
             14'h2ffb 	:	val_out <= 16'hec78;
             14'h2ffc 	:	val_out <= 16'hec7a;
             14'h2ffd 	:	val_out <= 16'hec7d;
             14'h2ffe 	:	val_out <= 16'hec7f;
             14'h2fff 	:	val_out <= 16'hec82;
             14'h3000 	:	val_out <= 16'hec84;
             14'h3001 	:	val_out <= 16'hec86;
             14'h3002 	:	val_out <= 16'hec89;
             14'h3003 	:	val_out <= 16'hec8b;
             14'h3004 	:	val_out <= 16'hec8e;
             14'h3005 	:	val_out <= 16'hec90;
             14'h3006 	:	val_out <= 16'hec92;
             14'h3007 	:	val_out <= 16'hec95;
             14'h3008 	:	val_out <= 16'hec97;
             14'h3009 	:	val_out <= 16'hec9a;
             14'h300a 	:	val_out <= 16'hec9c;
             14'h300b 	:	val_out <= 16'hec9e;
             14'h300c 	:	val_out <= 16'heca1;
             14'h300d 	:	val_out <= 16'heca3;
             14'h300e 	:	val_out <= 16'heca6;
             14'h300f 	:	val_out <= 16'heca8;
             14'h3010 	:	val_out <= 16'hecaa;
             14'h3011 	:	val_out <= 16'hecad;
             14'h3012 	:	val_out <= 16'hecaf;
             14'h3013 	:	val_out <= 16'hecb2;
             14'h3014 	:	val_out <= 16'hecb4;
             14'h3015 	:	val_out <= 16'hecb6;
             14'h3016 	:	val_out <= 16'hecb9;
             14'h3017 	:	val_out <= 16'hecbb;
             14'h3018 	:	val_out <= 16'hecbe;
             14'h3019 	:	val_out <= 16'hecc0;
             14'h301a 	:	val_out <= 16'hecc2;
             14'h301b 	:	val_out <= 16'hecc5;
             14'h301c 	:	val_out <= 16'hecc7;
             14'h301d 	:	val_out <= 16'hecca;
             14'h301e 	:	val_out <= 16'heccc;
             14'h301f 	:	val_out <= 16'hecce;
             14'h3020 	:	val_out <= 16'hecd1;
             14'h3021 	:	val_out <= 16'hecd3;
             14'h3022 	:	val_out <= 16'hecd5;
             14'h3023 	:	val_out <= 16'hecd8;
             14'h3024 	:	val_out <= 16'hecda;
             14'h3025 	:	val_out <= 16'hecdd;
             14'h3026 	:	val_out <= 16'hecdf;
             14'h3027 	:	val_out <= 16'hece1;
             14'h3028 	:	val_out <= 16'hece4;
             14'h3029 	:	val_out <= 16'hece6;
             14'h302a 	:	val_out <= 16'hece9;
             14'h302b 	:	val_out <= 16'heceb;
             14'h302c 	:	val_out <= 16'heced;
             14'h302d 	:	val_out <= 16'hecf0;
             14'h302e 	:	val_out <= 16'hecf2;
             14'h302f 	:	val_out <= 16'hecf4;
             14'h3030 	:	val_out <= 16'hecf7;
             14'h3031 	:	val_out <= 16'hecf9;
             14'h3032 	:	val_out <= 16'hecfc;
             14'h3033 	:	val_out <= 16'hecfe;
             14'h3034 	:	val_out <= 16'hed00;
             14'h3035 	:	val_out <= 16'hed03;
             14'h3036 	:	val_out <= 16'hed05;
             14'h3037 	:	val_out <= 16'hed07;
             14'h3038 	:	val_out <= 16'hed0a;
             14'h3039 	:	val_out <= 16'hed0c;
             14'h303a 	:	val_out <= 16'hed0f;
             14'h303b 	:	val_out <= 16'hed11;
             14'h303c 	:	val_out <= 16'hed13;
             14'h303d 	:	val_out <= 16'hed16;
             14'h303e 	:	val_out <= 16'hed18;
             14'h303f 	:	val_out <= 16'hed1a;
             14'h3040 	:	val_out <= 16'hed1d;
             14'h3041 	:	val_out <= 16'hed1f;
             14'h3042 	:	val_out <= 16'hed22;
             14'h3043 	:	val_out <= 16'hed24;
             14'h3044 	:	val_out <= 16'hed26;
             14'h3045 	:	val_out <= 16'hed29;
             14'h3046 	:	val_out <= 16'hed2b;
             14'h3047 	:	val_out <= 16'hed2d;
             14'h3048 	:	val_out <= 16'hed30;
             14'h3049 	:	val_out <= 16'hed32;
             14'h304a 	:	val_out <= 16'hed34;
             14'h304b 	:	val_out <= 16'hed37;
             14'h304c 	:	val_out <= 16'hed39;
             14'h304d 	:	val_out <= 16'hed3c;
             14'h304e 	:	val_out <= 16'hed3e;
             14'h304f 	:	val_out <= 16'hed40;
             14'h3050 	:	val_out <= 16'hed43;
             14'h3051 	:	val_out <= 16'hed45;
             14'h3052 	:	val_out <= 16'hed47;
             14'h3053 	:	val_out <= 16'hed4a;
             14'h3054 	:	val_out <= 16'hed4c;
             14'h3055 	:	val_out <= 16'hed4e;
             14'h3056 	:	val_out <= 16'hed51;
             14'h3057 	:	val_out <= 16'hed53;
             14'h3058 	:	val_out <= 16'hed55;
             14'h3059 	:	val_out <= 16'hed58;
             14'h305a 	:	val_out <= 16'hed5a;
             14'h305b 	:	val_out <= 16'hed5d;
             14'h305c 	:	val_out <= 16'hed5f;
             14'h305d 	:	val_out <= 16'hed61;
             14'h305e 	:	val_out <= 16'hed64;
             14'h305f 	:	val_out <= 16'hed66;
             14'h3060 	:	val_out <= 16'hed68;
             14'h3061 	:	val_out <= 16'hed6b;
             14'h3062 	:	val_out <= 16'hed6d;
             14'h3063 	:	val_out <= 16'hed6f;
             14'h3064 	:	val_out <= 16'hed72;
             14'h3065 	:	val_out <= 16'hed74;
             14'h3066 	:	val_out <= 16'hed76;
             14'h3067 	:	val_out <= 16'hed79;
             14'h3068 	:	val_out <= 16'hed7b;
             14'h3069 	:	val_out <= 16'hed7d;
             14'h306a 	:	val_out <= 16'hed80;
             14'h306b 	:	val_out <= 16'hed82;
             14'h306c 	:	val_out <= 16'hed84;
             14'h306d 	:	val_out <= 16'hed87;
             14'h306e 	:	val_out <= 16'hed89;
             14'h306f 	:	val_out <= 16'hed8c;
             14'h3070 	:	val_out <= 16'hed8e;
             14'h3071 	:	val_out <= 16'hed90;
             14'h3072 	:	val_out <= 16'hed93;
             14'h3073 	:	val_out <= 16'hed95;
             14'h3074 	:	val_out <= 16'hed97;
             14'h3075 	:	val_out <= 16'hed9a;
             14'h3076 	:	val_out <= 16'hed9c;
             14'h3077 	:	val_out <= 16'hed9e;
             14'h3078 	:	val_out <= 16'heda1;
             14'h3079 	:	val_out <= 16'heda3;
             14'h307a 	:	val_out <= 16'heda5;
             14'h307b 	:	val_out <= 16'heda8;
             14'h307c 	:	val_out <= 16'hedaa;
             14'h307d 	:	val_out <= 16'hedac;
             14'h307e 	:	val_out <= 16'hedaf;
             14'h307f 	:	val_out <= 16'hedb1;
             14'h3080 	:	val_out <= 16'hedb3;
             14'h3081 	:	val_out <= 16'hedb6;
             14'h3082 	:	val_out <= 16'hedb8;
             14'h3083 	:	val_out <= 16'hedba;
             14'h3084 	:	val_out <= 16'hedbd;
             14'h3085 	:	val_out <= 16'hedbf;
             14'h3086 	:	val_out <= 16'hedc1;
             14'h3087 	:	val_out <= 16'hedc4;
             14'h3088 	:	val_out <= 16'hedc6;
             14'h3089 	:	val_out <= 16'hedc8;
             14'h308a 	:	val_out <= 16'hedcb;
             14'h308b 	:	val_out <= 16'hedcd;
             14'h308c 	:	val_out <= 16'hedcf;
             14'h308d 	:	val_out <= 16'hedd2;
             14'h308e 	:	val_out <= 16'hedd4;
             14'h308f 	:	val_out <= 16'hedd6;
             14'h3090 	:	val_out <= 16'hedd8;
             14'h3091 	:	val_out <= 16'heddb;
             14'h3092 	:	val_out <= 16'heddd;
             14'h3093 	:	val_out <= 16'heddf;
             14'h3094 	:	val_out <= 16'hede2;
             14'h3095 	:	val_out <= 16'hede4;
             14'h3096 	:	val_out <= 16'hede6;
             14'h3097 	:	val_out <= 16'hede9;
             14'h3098 	:	val_out <= 16'hedeb;
             14'h3099 	:	val_out <= 16'heded;
             14'h309a 	:	val_out <= 16'hedf0;
             14'h309b 	:	val_out <= 16'hedf2;
             14'h309c 	:	val_out <= 16'hedf4;
             14'h309d 	:	val_out <= 16'hedf7;
             14'h309e 	:	val_out <= 16'hedf9;
             14'h309f 	:	val_out <= 16'hedfb;
             14'h30a0 	:	val_out <= 16'hedfe;
             14'h30a1 	:	val_out <= 16'hee00;
             14'h30a2 	:	val_out <= 16'hee02;
             14'h30a3 	:	val_out <= 16'hee05;
             14'h30a4 	:	val_out <= 16'hee07;
             14'h30a5 	:	val_out <= 16'hee09;
             14'h30a6 	:	val_out <= 16'hee0b;
             14'h30a7 	:	val_out <= 16'hee0e;
             14'h30a8 	:	val_out <= 16'hee10;
             14'h30a9 	:	val_out <= 16'hee12;
             14'h30aa 	:	val_out <= 16'hee15;
             14'h30ab 	:	val_out <= 16'hee17;
             14'h30ac 	:	val_out <= 16'hee19;
             14'h30ad 	:	val_out <= 16'hee1c;
             14'h30ae 	:	val_out <= 16'hee1e;
             14'h30af 	:	val_out <= 16'hee20;
             14'h30b0 	:	val_out <= 16'hee23;
             14'h30b1 	:	val_out <= 16'hee25;
             14'h30b2 	:	val_out <= 16'hee27;
             14'h30b3 	:	val_out <= 16'hee29;
             14'h30b4 	:	val_out <= 16'hee2c;
             14'h30b5 	:	val_out <= 16'hee2e;
             14'h30b6 	:	val_out <= 16'hee30;
             14'h30b7 	:	val_out <= 16'hee33;
             14'h30b8 	:	val_out <= 16'hee35;
             14'h30b9 	:	val_out <= 16'hee37;
             14'h30ba 	:	val_out <= 16'hee3a;
             14'h30bb 	:	val_out <= 16'hee3c;
             14'h30bc 	:	val_out <= 16'hee3e;
             14'h30bd 	:	val_out <= 16'hee40;
             14'h30be 	:	val_out <= 16'hee43;
             14'h30bf 	:	val_out <= 16'hee45;
             14'h30c0 	:	val_out <= 16'hee47;
             14'h30c1 	:	val_out <= 16'hee4a;
             14'h30c2 	:	val_out <= 16'hee4c;
             14'h30c3 	:	val_out <= 16'hee4e;
             14'h30c4 	:	val_out <= 16'hee51;
             14'h30c5 	:	val_out <= 16'hee53;
             14'h30c6 	:	val_out <= 16'hee55;
             14'h30c7 	:	val_out <= 16'hee57;
             14'h30c8 	:	val_out <= 16'hee5a;
             14'h30c9 	:	val_out <= 16'hee5c;
             14'h30ca 	:	val_out <= 16'hee5e;
             14'h30cb 	:	val_out <= 16'hee61;
             14'h30cc 	:	val_out <= 16'hee63;
             14'h30cd 	:	val_out <= 16'hee65;
             14'h30ce 	:	val_out <= 16'hee67;
             14'h30cf 	:	val_out <= 16'hee6a;
             14'h30d0 	:	val_out <= 16'hee6c;
             14'h30d1 	:	val_out <= 16'hee6e;
             14'h30d2 	:	val_out <= 16'hee71;
             14'h30d3 	:	val_out <= 16'hee73;
             14'h30d4 	:	val_out <= 16'hee75;
             14'h30d5 	:	val_out <= 16'hee78;
             14'h30d6 	:	val_out <= 16'hee7a;
             14'h30d7 	:	val_out <= 16'hee7c;
             14'h30d8 	:	val_out <= 16'hee7e;
             14'h30d9 	:	val_out <= 16'hee81;
             14'h30da 	:	val_out <= 16'hee83;
             14'h30db 	:	val_out <= 16'hee85;
             14'h30dc 	:	val_out <= 16'hee87;
             14'h30dd 	:	val_out <= 16'hee8a;
             14'h30de 	:	val_out <= 16'hee8c;
             14'h30df 	:	val_out <= 16'hee8e;
             14'h30e0 	:	val_out <= 16'hee91;
             14'h30e1 	:	val_out <= 16'hee93;
             14'h30e2 	:	val_out <= 16'hee95;
             14'h30e3 	:	val_out <= 16'hee97;
             14'h30e4 	:	val_out <= 16'hee9a;
             14'h30e5 	:	val_out <= 16'hee9c;
             14'h30e6 	:	val_out <= 16'hee9e;
             14'h30e7 	:	val_out <= 16'heea1;
             14'h30e8 	:	val_out <= 16'heea3;
             14'h30e9 	:	val_out <= 16'heea5;
             14'h30ea 	:	val_out <= 16'heea7;
             14'h30eb 	:	val_out <= 16'heeaa;
             14'h30ec 	:	val_out <= 16'heeac;
             14'h30ed 	:	val_out <= 16'heeae;
             14'h30ee 	:	val_out <= 16'heeb0;
             14'h30ef 	:	val_out <= 16'heeb3;
             14'h30f0 	:	val_out <= 16'heeb5;
             14'h30f1 	:	val_out <= 16'heeb7;
             14'h30f2 	:	val_out <= 16'heeba;
             14'h30f3 	:	val_out <= 16'heebc;
             14'h30f4 	:	val_out <= 16'heebe;
             14'h30f5 	:	val_out <= 16'heec0;
             14'h30f6 	:	val_out <= 16'heec3;
             14'h30f7 	:	val_out <= 16'heec5;
             14'h30f8 	:	val_out <= 16'heec7;
             14'h30f9 	:	val_out <= 16'heec9;
             14'h30fa 	:	val_out <= 16'heecc;
             14'h30fb 	:	val_out <= 16'heece;
             14'h30fc 	:	val_out <= 16'heed0;
             14'h30fd 	:	val_out <= 16'heed2;
             14'h30fe 	:	val_out <= 16'heed5;
             14'h30ff 	:	val_out <= 16'heed7;
             14'h3100 	:	val_out <= 16'heed9;
             14'h3101 	:	val_out <= 16'heedc;
             14'h3102 	:	val_out <= 16'heede;
             14'h3103 	:	val_out <= 16'heee0;
             14'h3104 	:	val_out <= 16'heee2;
             14'h3105 	:	val_out <= 16'heee5;
             14'h3106 	:	val_out <= 16'heee7;
             14'h3107 	:	val_out <= 16'heee9;
             14'h3108 	:	val_out <= 16'heeeb;
             14'h3109 	:	val_out <= 16'heeee;
             14'h310a 	:	val_out <= 16'heef0;
             14'h310b 	:	val_out <= 16'heef2;
             14'h310c 	:	val_out <= 16'heef4;
             14'h310d 	:	val_out <= 16'heef7;
             14'h310e 	:	val_out <= 16'heef9;
             14'h310f 	:	val_out <= 16'heefb;
             14'h3110 	:	val_out <= 16'heefd;
             14'h3111 	:	val_out <= 16'hef00;
             14'h3112 	:	val_out <= 16'hef02;
             14'h3113 	:	val_out <= 16'hef04;
             14'h3114 	:	val_out <= 16'hef06;
             14'h3115 	:	val_out <= 16'hef09;
             14'h3116 	:	val_out <= 16'hef0b;
             14'h3117 	:	val_out <= 16'hef0d;
             14'h3118 	:	val_out <= 16'hef0f;
             14'h3119 	:	val_out <= 16'hef12;
             14'h311a 	:	val_out <= 16'hef14;
             14'h311b 	:	val_out <= 16'hef16;
             14'h311c 	:	val_out <= 16'hef18;
             14'h311d 	:	val_out <= 16'hef1b;
             14'h311e 	:	val_out <= 16'hef1d;
             14'h311f 	:	val_out <= 16'hef1f;
             14'h3120 	:	val_out <= 16'hef21;
             14'h3121 	:	val_out <= 16'hef24;
             14'h3122 	:	val_out <= 16'hef26;
             14'h3123 	:	val_out <= 16'hef28;
             14'h3124 	:	val_out <= 16'hef2a;
             14'h3125 	:	val_out <= 16'hef2d;
             14'h3126 	:	val_out <= 16'hef2f;
             14'h3127 	:	val_out <= 16'hef31;
             14'h3128 	:	val_out <= 16'hef33;
             14'h3129 	:	val_out <= 16'hef35;
             14'h312a 	:	val_out <= 16'hef38;
             14'h312b 	:	val_out <= 16'hef3a;
             14'h312c 	:	val_out <= 16'hef3c;
             14'h312d 	:	val_out <= 16'hef3e;
             14'h312e 	:	val_out <= 16'hef41;
             14'h312f 	:	val_out <= 16'hef43;
             14'h3130 	:	val_out <= 16'hef45;
             14'h3131 	:	val_out <= 16'hef47;
             14'h3132 	:	val_out <= 16'hef4a;
             14'h3133 	:	val_out <= 16'hef4c;
             14'h3134 	:	val_out <= 16'hef4e;
             14'h3135 	:	val_out <= 16'hef50;
             14'h3136 	:	val_out <= 16'hef53;
             14'h3137 	:	val_out <= 16'hef55;
             14'h3138 	:	val_out <= 16'hef57;
             14'h3139 	:	val_out <= 16'hef59;
             14'h313a 	:	val_out <= 16'hef5b;
             14'h313b 	:	val_out <= 16'hef5e;
             14'h313c 	:	val_out <= 16'hef60;
             14'h313d 	:	val_out <= 16'hef62;
             14'h313e 	:	val_out <= 16'hef64;
             14'h313f 	:	val_out <= 16'hef67;
             14'h3140 	:	val_out <= 16'hef69;
             14'h3141 	:	val_out <= 16'hef6b;
             14'h3142 	:	val_out <= 16'hef6d;
             14'h3143 	:	val_out <= 16'hef6f;
             14'h3144 	:	val_out <= 16'hef72;
             14'h3145 	:	val_out <= 16'hef74;
             14'h3146 	:	val_out <= 16'hef76;
             14'h3147 	:	val_out <= 16'hef78;
             14'h3148 	:	val_out <= 16'hef7b;
             14'h3149 	:	val_out <= 16'hef7d;
             14'h314a 	:	val_out <= 16'hef7f;
             14'h314b 	:	val_out <= 16'hef81;
             14'h314c 	:	val_out <= 16'hef83;
             14'h314d 	:	val_out <= 16'hef86;
             14'h314e 	:	val_out <= 16'hef88;
             14'h314f 	:	val_out <= 16'hef8a;
             14'h3150 	:	val_out <= 16'hef8c;
             14'h3151 	:	val_out <= 16'hef8f;
             14'h3152 	:	val_out <= 16'hef91;
             14'h3153 	:	val_out <= 16'hef93;
             14'h3154 	:	val_out <= 16'hef95;
             14'h3155 	:	val_out <= 16'hef97;
             14'h3156 	:	val_out <= 16'hef9a;
             14'h3157 	:	val_out <= 16'hef9c;
             14'h3158 	:	val_out <= 16'hef9e;
             14'h3159 	:	val_out <= 16'hefa0;
             14'h315a 	:	val_out <= 16'hefa2;
             14'h315b 	:	val_out <= 16'hefa5;
             14'h315c 	:	val_out <= 16'hefa7;
             14'h315d 	:	val_out <= 16'hefa9;
             14'h315e 	:	val_out <= 16'hefab;
             14'h315f 	:	val_out <= 16'hefae;
             14'h3160 	:	val_out <= 16'hefb0;
             14'h3161 	:	val_out <= 16'hefb2;
             14'h3162 	:	val_out <= 16'hefb4;
             14'h3163 	:	val_out <= 16'hefb6;
             14'h3164 	:	val_out <= 16'hefb9;
             14'h3165 	:	val_out <= 16'hefbb;
             14'h3166 	:	val_out <= 16'hefbd;
             14'h3167 	:	val_out <= 16'hefbf;
             14'h3168 	:	val_out <= 16'hefc1;
             14'h3169 	:	val_out <= 16'hefc4;
             14'h316a 	:	val_out <= 16'hefc6;
             14'h316b 	:	val_out <= 16'hefc8;
             14'h316c 	:	val_out <= 16'hefca;
             14'h316d 	:	val_out <= 16'hefcc;
             14'h316e 	:	val_out <= 16'hefcf;
             14'h316f 	:	val_out <= 16'hefd1;
             14'h3170 	:	val_out <= 16'hefd3;
             14'h3171 	:	val_out <= 16'hefd5;
             14'h3172 	:	val_out <= 16'hefd7;
             14'h3173 	:	val_out <= 16'hefda;
             14'h3174 	:	val_out <= 16'hefdc;
             14'h3175 	:	val_out <= 16'hefde;
             14'h3176 	:	val_out <= 16'hefe0;
             14'h3177 	:	val_out <= 16'hefe2;
             14'h3178 	:	val_out <= 16'hefe5;
             14'h3179 	:	val_out <= 16'hefe7;
             14'h317a 	:	val_out <= 16'hefe9;
             14'h317b 	:	val_out <= 16'hefeb;
             14'h317c 	:	val_out <= 16'hefed;
             14'h317d 	:	val_out <= 16'hefef;
             14'h317e 	:	val_out <= 16'heff2;
             14'h317f 	:	val_out <= 16'heff4;
             14'h3180 	:	val_out <= 16'heff6;
             14'h3181 	:	val_out <= 16'heff8;
             14'h3182 	:	val_out <= 16'heffa;
             14'h3183 	:	val_out <= 16'heffd;
             14'h3184 	:	val_out <= 16'hefff;
             14'h3185 	:	val_out <= 16'hf001;
             14'h3186 	:	val_out <= 16'hf003;
             14'h3187 	:	val_out <= 16'hf005;
             14'h3188 	:	val_out <= 16'hf008;
             14'h3189 	:	val_out <= 16'hf00a;
             14'h318a 	:	val_out <= 16'hf00c;
             14'h318b 	:	val_out <= 16'hf00e;
             14'h318c 	:	val_out <= 16'hf010;
             14'h318d 	:	val_out <= 16'hf012;
             14'h318e 	:	val_out <= 16'hf015;
             14'h318f 	:	val_out <= 16'hf017;
             14'h3190 	:	val_out <= 16'hf019;
             14'h3191 	:	val_out <= 16'hf01b;
             14'h3192 	:	val_out <= 16'hf01d;
             14'h3193 	:	val_out <= 16'hf020;
             14'h3194 	:	val_out <= 16'hf022;
             14'h3195 	:	val_out <= 16'hf024;
             14'h3196 	:	val_out <= 16'hf026;
             14'h3197 	:	val_out <= 16'hf028;
             14'h3198 	:	val_out <= 16'hf02a;
             14'h3199 	:	val_out <= 16'hf02d;
             14'h319a 	:	val_out <= 16'hf02f;
             14'h319b 	:	val_out <= 16'hf031;
             14'h319c 	:	val_out <= 16'hf033;
             14'h319d 	:	val_out <= 16'hf035;
             14'h319e 	:	val_out <= 16'hf037;
             14'h319f 	:	val_out <= 16'hf03a;
             14'h31a0 	:	val_out <= 16'hf03c;
             14'h31a1 	:	val_out <= 16'hf03e;
             14'h31a2 	:	val_out <= 16'hf040;
             14'h31a3 	:	val_out <= 16'hf042;
             14'h31a4 	:	val_out <= 16'hf044;
             14'h31a5 	:	val_out <= 16'hf047;
             14'h31a6 	:	val_out <= 16'hf049;
             14'h31a7 	:	val_out <= 16'hf04b;
             14'h31a8 	:	val_out <= 16'hf04d;
             14'h31a9 	:	val_out <= 16'hf04f;
             14'h31aa 	:	val_out <= 16'hf051;
             14'h31ab 	:	val_out <= 16'hf054;
             14'h31ac 	:	val_out <= 16'hf056;
             14'h31ad 	:	val_out <= 16'hf058;
             14'h31ae 	:	val_out <= 16'hf05a;
             14'h31af 	:	val_out <= 16'hf05c;
             14'h31b0 	:	val_out <= 16'hf05e;
             14'h31b1 	:	val_out <= 16'hf061;
             14'h31b2 	:	val_out <= 16'hf063;
             14'h31b3 	:	val_out <= 16'hf065;
             14'h31b4 	:	val_out <= 16'hf067;
             14'h31b5 	:	val_out <= 16'hf069;
             14'h31b6 	:	val_out <= 16'hf06b;
             14'h31b7 	:	val_out <= 16'hf06e;
             14'h31b8 	:	val_out <= 16'hf070;
             14'h31b9 	:	val_out <= 16'hf072;
             14'h31ba 	:	val_out <= 16'hf074;
             14'h31bb 	:	val_out <= 16'hf076;
             14'h31bc 	:	val_out <= 16'hf078;
             14'h31bd 	:	val_out <= 16'hf07b;
             14'h31be 	:	val_out <= 16'hf07d;
             14'h31bf 	:	val_out <= 16'hf07f;
             14'h31c0 	:	val_out <= 16'hf081;
             14'h31c1 	:	val_out <= 16'hf083;
             14'h31c2 	:	val_out <= 16'hf085;
             14'h31c3 	:	val_out <= 16'hf087;
             14'h31c4 	:	val_out <= 16'hf08a;
             14'h31c5 	:	val_out <= 16'hf08c;
             14'h31c6 	:	val_out <= 16'hf08e;
             14'h31c7 	:	val_out <= 16'hf090;
             14'h31c8 	:	val_out <= 16'hf092;
             14'h31c9 	:	val_out <= 16'hf094;
             14'h31ca 	:	val_out <= 16'hf096;
             14'h31cb 	:	val_out <= 16'hf099;
             14'h31cc 	:	val_out <= 16'hf09b;
             14'h31cd 	:	val_out <= 16'hf09d;
             14'h31ce 	:	val_out <= 16'hf09f;
             14'h31cf 	:	val_out <= 16'hf0a1;
             14'h31d0 	:	val_out <= 16'hf0a3;
             14'h31d1 	:	val_out <= 16'hf0a5;
             14'h31d2 	:	val_out <= 16'hf0a8;
             14'h31d3 	:	val_out <= 16'hf0aa;
             14'h31d4 	:	val_out <= 16'hf0ac;
             14'h31d5 	:	val_out <= 16'hf0ae;
             14'h31d6 	:	val_out <= 16'hf0b0;
             14'h31d7 	:	val_out <= 16'hf0b2;
             14'h31d8 	:	val_out <= 16'hf0b4;
             14'h31d9 	:	val_out <= 16'hf0b7;
             14'h31da 	:	val_out <= 16'hf0b9;
             14'h31db 	:	val_out <= 16'hf0bb;
             14'h31dc 	:	val_out <= 16'hf0bd;
             14'h31dd 	:	val_out <= 16'hf0bf;
             14'h31de 	:	val_out <= 16'hf0c1;
             14'h31df 	:	val_out <= 16'hf0c3;
             14'h31e0 	:	val_out <= 16'hf0c6;
             14'h31e1 	:	val_out <= 16'hf0c8;
             14'h31e2 	:	val_out <= 16'hf0ca;
             14'h31e3 	:	val_out <= 16'hf0cc;
             14'h31e4 	:	val_out <= 16'hf0ce;
             14'h31e5 	:	val_out <= 16'hf0d0;
             14'h31e6 	:	val_out <= 16'hf0d2;
             14'h31e7 	:	val_out <= 16'hf0d5;
             14'h31e8 	:	val_out <= 16'hf0d7;
             14'h31e9 	:	val_out <= 16'hf0d9;
             14'h31ea 	:	val_out <= 16'hf0db;
             14'h31eb 	:	val_out <= 16'hf0dd;
             14'h31ec 	:	val_out <= 16'hf0df;
             14'h31ed 	:	val_out <= 16'hf0e1;
             14'h31ee 	:	val_out <= 16'hf0e3;
             14'h31ef 	:	val_out <= 16'hf0e6;
             14'h31f0 	:	val_out <= 16'hf0e8;
             14'h31f1 	:	val_out <= 16'hf0ea;
             14'h31f2 	:	val_out <= 16'hf0ec;
             14'h31f3 	:	val_out <= 16'hf0ee;
             14'h31f4 	:	val_out <= 16'hf0f0;
             14'h31f5 	:	val_out <= 16'hf0f2;
             14'h31f6 	:	val_out <= 16'hf0f4;
             14'h31f7 	:	val_out <= 16'hf0f7;
             14'h31f8 	:	val_out <= 16'hf0f9;
             14'h31f9 	:	val_out <= 16'hf0fb;
             14'h31fa 	:	val_out <= 16'hf0fd;
             14'h31fb 	:	val_out <= 16'hf0ff;
             14'h31fc 	:	val_out <= 16'hf101;
             14'h31fd 	:	val_out <= 16'hf103;
             14'h31fe 	:	val_out <= 16'hf105;
             14'h31ff 	:	val_out <= 16'hf107;
             14'h3200 	:	val_out <= 16'hf10a;
             14'h3201 	:	val_out <= 16'hf10c;
             14'h3202 	:	val_out <= 16'hf10e;
             14'h3203 	:	val_out <= 16'hf110;
             14'h3204 	:	val_out <= 16'hf112;
             14'h3205 	:	val_out <= 16'hf114;
             14'h3206 	:	val_out <= 16'hf116;
             14'h3207 	:	val_out <= 16'hf118;
             14'h3208 	:	val_out <= 16'hf11b;
             14'h3209 	:	val_out <= 16'hf11d;
             14'h320a 	:	val_out <= 16'hf11f;
             14'h320b 	:	val_out <= 16'hf121;
             14'h320c 	:	val_out <= 16'hf123;
             14'h320d 	:	val_out <= 16'hf125;
             14'h320e 	:	val_out <= 16'hf127;
             14'h320f 	:	val_out <= 16'hf129;
             14'h3210 	:	val_out <= 16'hf12b;
             14'h3211 	:	val_out <= 16'hf12d;
             14'h3212 	:	val_out <= 16'hf130;
             14'h3213 	:	val_out <= 16'hf132;
             14'h3214 	:	val_out <= 16'hf134;
             14'h3215 	:	val_out <= 16'hf136;
             14'h3216 	:	val_out <= 16'hf138;
             14'h3217 	:	val_out <= 16'hf13a;
             14'h3218 	:	val_out <= 16'hf13c;
             14'h3219 	:	val_out <= 16'hf13e;
             14'h321a 	:	val_out <= 16'hf140;
             14'h321b 	:	val_out <= 16'hf143;
             14'h321c 	:	val_out <= 16'hf145;
             14'h321d 	:	val_out <= 16'hf147;
             14'h321e 	:	val_out <= 16'hf149;
             14'h321f 	:	val_out <= 16'hf14b;
             14'h3220 	:	val_out <= 16'hf14d;
             14'h3221 	:	val_out <= 16'hf14f;
             14'h3222 	:	val_out <= 16'hf151;
             14'h3223 	:	val_out <= 16'hf153;
             14'h3224 	:	val_out <= 16'hf155;
             14'h3225 	:	val_out <= 16'hf158;
             14'h3226 	:	val_out <= 16'hf15a;
             14'h3227 	:	val_out <= 16'hf15c;
             14'h3228 	:	val_out <= 16'hf15e;
             14'h3229 	:	val_out <= 16'hf160;
             14'h322a 	:	val_out <= 16'hf162;
             14'h322b 	:	val_out <= 16'hf164;
             14'h322c 	:	val_out <= 16'hf166;
             14'h322d 	:	val_out <= 16'hf168;
             14'h322e 	:	val_out <= 16'hf16a;
             14'h322f 	:	val_out <= 16'hf16c;
             14'h3230 	:	val_out <= 16'hf16f;
             14'h3231 	:	val_out <= 16'hf171;
             14'h3232 	:	val_out <= 16'hf173;
             14'h3233 	:	val_out <= 16'hf175;
             14'h3234 	:	val_out <= 16'hf177;
             14'h3235 	:	val_out <= 16'hf179;
             14'h3236 	:	val_out <= 16'hf17b;
             14'h3237 	:	val_out <= 16'hf17d;
             14'h3238 	:	val_out <= 16'hf17f;
             14'h3239 	:	val_out <= 16'hf181;
             14'h323a 	:	val_out <= 16'hf183;
             14'h323b 	:	val_out <= 16'hf185;
             14'h323c 	:	val_out <= 16'hf188;
             14'h323d 	:	val_out <= 16'hf18a;
             14'h323e 	:	val_out <= 16'hf18c;
             14'h323f 	:	val_out <= 16'hf18e;
             14'h3240 	:	val_out <= 16'hf190;
             14'h3241 	:	val_out <= 16'hf192;
             14'h3242 	:	val_out <= 16'hf194;
             14'h3243 	:	val_out <= 16'hf196;
             14'h3244 	:	val_out <= 16'hf198;
             14'h3245 	:	val_out <= 16'hf19a;
             14'h3246 	:	val_out <= 16'hf19c;
             14'h3247 	:	val_out <= 16'hf19e;
             14'h3248 	:	val_out <= 16'hf1a1;
             14'h3249 	:	val_out <= 16'hf1a3;
             14'h324a 	:	val_out <= 16'hf1a5;
             14'h324b 	:	val_out <= 16'hf1a7;
             14'h324c 	:	val_out <= 16'hf1a9;
             14'h324d 	:	val_out <= 16'hf1ab;
             14'h324e 	:	val_out <= 16'hf1ad;
             14'h324f 	:	val_out <= 16'hf1af;
             14'h3250 	:	val_out <= 16'hf1b1;
             14'h3251 	:	val_out <= 16'hf1b3;
             14'h3252 	:	val_out <= 16'hf1b5;
             14'h3253 	:	val_out <= 16'hf1b7;
             14'h3254 	:	val_out <= 16'hf1b9;
             14'h3255 	:	val_out <= 16'hf1bb;
             14'h3256 	:	val_out <= 16'hf1be;
             14'h3257 	:	val_out <= 16'hf1c0;
             14'h3258 	:	val_out <= 16'hf1c2;
             14'h3259 	:	val_out <= 16'hf1c4;
             14'h325a 	:	val_out <= 16'hf1c6;
             14'h325b 	:	val_out <= 16'hf1c8;
             14'h325c 	:	val_out <= 16'hf1ca;
             14'h325d 	:	val_out <= 16'hf1cc;
             14'h325e 	:	val_out <= 16'hf1ce;
             14'h325f 	:	val_out <= 16'hf1d0;
             14'h3260 	:	val_out <= 16'hf1d2;
             14'h3261 	:	val_out <= 16'hf1d4;
             14'h3262 	:	val_out <= 16'hf1d6;
             14'h3263 	:	val_out <= 16'hf1d8;
             14'h3264 	:	val_out <= 16'hf1da;
             14'h3265 	:	val_out <= 16'hf1dc;
             14'h3266 	:	val_out <= 16'hf1df;
             14'h3267 	:	val_out <= 16'hf1e1;
             14'h3268 	:	val_out <= 16'hf1e3;
             14'h3269 	:	val_out <= 16'hf1e5;
             14'h326a 	:	val_out <= 16'hf1e7;
             14'h326b 	:	val_out <= 16'hf1e9;
             14'h326c 	:	val_out <= 16'hf1eb;
             14'h326d 	:	val_out <= 16'hf1ed;
             14'h326e 	:	val_out <= 16'hf1ef;
             14'h326f 	:	val_out <= 16'hf1f1;
             14'h3270 	:	val_out <= 16'hf1f3;
             14'h3271 	:	val_out <= 16'hf1f5;
             14'h3272 	:	val_out <= 16'hf1f7;
             14'h3273 	:	val_out <= 16'hf1f9;
             14'h3274 	:	val_out <= 16'hf1fb;
             14'h3275 	:	val_out <= 16'hf1fd;
             14'h3276 	:	val_out <= 16'hf1ff;
             14'h3277 	:	val_out <= 16'hf201;
             14'h3278 	:	val_out <= 16'hf203;
             14'h3279 	:	val_out <= 16'hf206;
             14'h327a 	:	val_out <= 16'hf208;
             14'h327b 	:	val_out <= 16'hf20a;
             14'h327c 	:	val_out <= 16'hf20c;
             14'h327d 	:	val_out <= 16'hf20e;
             14'h327e 	:	val_out <= 16'hf210;
             14'h327f 	:	val_out <= 16'hf212;
             14'h3280 	:	val_out <= 16'hf214;
             14'h3281 	:	val_out <= 16'hf216;
             14'h3282 	:	val_out <= 16'hf218;
             14'h3283 	:	val_out <= 16'hf21a;
             14'h3284 	:	val_out <= 16'hf21c;
             14'h3285 	:	val_out <= 16'hf21e;
             14'h3286 	:	val_out <= 16'hf220;
             14'h3287 	:	val_out <= 16'hf222;
             14'h3288 	:	val_out <= 16'hf224;
             14'h3289 	:	val_out <= 16'hf226;
             14'h328a 	:	val_out <= 16'hf228;
             14'h328b 	:	val_out <= 16'hf22a;
             14'h328c 	:	val_out <= 16'hf22c;
             14'h328d 	:	val_out <= 16'hf22e;
             14'h328e 	:	val_out <= 16'hf230;
             14'h328f 	:	val_out <= 16'hf232;
             14'h3290 	:	val_out <= 16'hf234;
             14'h3291 	:	val_out <= 16'hf237;
             14'h3292 	:	val_out <= 16'hf239;
             14'h3293 	:	val_out <= 16'hf23b;
             14'h3294 	:	val_out <= 16'hf23d;
             14'h3295 	:	val_out <= 16'hf23f;
             14'h3296 	:	val_out <= 16'hf241;
             14'h3297 	:	val_out <= 16'hf243;
             14'h3298 	:	val_out <= 16'hf245;
             14'h3299 	:	val_out <= 16'hf247;
             14'h329a 	:	val_out <= 16'hf249;
             14'h329b 	:	val_out <= 16'hf24b;
             14'h329c 	:	val_out <= 16'hf24d;
             14'h329d 	:	val_out <= 16'hf24f;
             14'h329e 	:	val_out <= 16'hf251;
             14'h329f 	:	val_out <= 16'hf253;
             14'h32a0 	:	val_out <= 16'hf255;
             14'h32a1 	:	val_out <= 16'hf257;
             14'h32a2 	:	val_out <= 16'hf259;
             14'h32a3 	:	val_out <= 16'hf25b;
             14'h32a4 	:	val_out <= 16'hf25d;
             14'h32a5 	:	val_out <= 16'hf25f;
             14'h32a6 	:	val_out <= 16'hf261;
             14'h32a7 	:	val_out <= 16'hf263;
             14'h32a8 	:	val_out <= 16'hf265;
             14'h32a9 	:	val_out <= 16'hf267;
             14'h32aa 	:	val_out <= 16'hf269;
             14'h32ab 	:	val_out <= 16'hf26b;
             14'h32ac 	:	val_out <= 16'hf26d;
             14'h32ad 	:	val_out <= 16'hf26f;
             14'h32ae 	:	val_out <= 16'hf271;
             14'h32af 	:	val_out <= 16'hf273;
             14'h32b0 	:	val_out <= 16'hf275;
             14'h32b1 	:	val_out <= 16'hf277;
             14'h32b2 	:	val_out <= 16'hf279;
             14'h32b3 	:	val_out <= 16'hf27b;
             14'h32b4 	:	val_out <= 16'hf27d;
             14'h32b5 	:	val_out <= 16'hf27f;
             14'h32b6 	:	val_out <= 16'hf281;
             14'h32b7 	:	val_out <= 16'hf283;
             14'h32b8 	:	val_out <= 16'hf285;
             14'h32b9 	:	val_out <= 16'hf287;
             14'h32ba 	:	val_out <= 16'hf289;
             14'h32bb 	:	val_out <= 16'hf28b;
             14'h32bc 	:	val_out <= 16'hf28d;
             14'h32bd 	:	val_out <= 16'hf28f;
             14'h32be 	:	val_out <= 16'hf291;
             14'h32bf 	:	val_out <= 16'hf293;
             14'h32c0 	:	val_out <= 16'hf295;
             14'h32c1 	:	val_out <= 16'hf297;
             14'h32c2 	:	val_out <= 16'hf299;
             14'h32c3 	:	val_out <= 16'hf29b;
             14'h32c4 	:	val_out <= 16'hf29d;
             14'h32c5 	:	val_out <= 16'hf2a0;
             14'h32c6 	:	val_out <= 16'hf2a2;
             14'h32c7 	:	val_out <= 16'hf2a4;
             14'h32c8 	:	val_out <= 16'hf2a6;
             14'h32c9 	:	val_out <= 16'hf2a8;
             14'h32ca 	:	val_out <= 16'hf2aa;
             14'h32cb 	:	val_out <= 16'hf2ac;
             14'h32cc 	:	val_out <= 16'hf2ae;
             14'h32cd 	:	val_out <= 16'hf2b0;
             14'h32ce 	:	val_out <= 16'hf2b2;
             14'h32cf 	:	val_out <= 16'hf2b4;
             14'h32d0 	:	val_out <= 16'hf2b6;
             14'h32d1 	:	val_out <= 16'hf2b8;
             14'h32d2 	:	val_out <= 16'hf2ba;
             14'h32d3 	:	val_out <= 16'hf2bc;
             14'h32d4 	:	val_out <= 16'hf2be;
             14'h32d5 	:	val_out <= 16'hf2bf;
             14'h32d6 	:	val_out <= 16'hf2c1;
             14'h32d7 	:	val_out <= 16'hf2c3;
             14'h32d8 	:	val_out <= 16'hf2c5;
             14'h32d9 	:	val_out <= 16'hf2c7;
             14'h32da 	:	val_out <= 16'hf2c9;
             14'h32db 	:	val_out <= 16'hf2cb;
             14'h32dc 	:	val_out <= 16'hf2cd;
             14'h32dd 	:	val_out <= 16'hf2cf;
             14'h32de 	:	val_out <= 16'hf2d1;
             14'h32df 	:	val_out <= 16'hf2d3;
             14'h32e0 	:	val_out <= 16'hf2d5;
             14'h32e1 	:	val_out <= 16'hf2d7;
             14'h32e2 	:	val_out <= 16'hf2d9;
             14'h32e3 	:	val_out <= 16'hf2db;
             14'h32e4 	:	val_out <= 16'hf2dd;
             14'h32e5 	:	val_out <= 16'hf2df;
             14'h32e6 	:	val_out <= 16'hf2e1;
             14'h32e7 	:	val_out <= 16'hf2e3;
             14'h32e8 	:	val_out <= 16'hf2e5;
             14'h32e9 	:	val_out <= 16'hf2e7;
             14'h32ea 	:	val_out <= 16'hf2e9;
             14'h32eb 	:	val_out <= 16'hf2eb;
             14'h32ec 	:	val_out <= 16'hf2ed;
             14'h32ed 	:	val_out <= 16'hf2ef;
             14'h32ee 	:	val_out <= 16'hf2f1;
             14'h32ef 	:	val_out <= 16'hf2f3;
             14'h32f0 	:	val_out <= 16'hf2f5;
             14'h32f1 	:	val_out <= 16'hf2f7;
             14'h32f2 	:	val_out <= 16'hf2f9;
             14'h32f3 	:	val_out <= 16'hf2fb;
             14'h32f4 	:	val_out <= 16'hf2fd;
             14'h32f5 	:	val_out <= 16'hf2ff;
             14'h32f6 	:	val_out <= 16'hf301;
             14'h32f7 	:	val_out <= 16'hf303;
             14'h32f8 	:	val_out <= 16'hf305;
             14'h32f9 	:	val_out <= 16'hf307;
             14'h32fa 	:	val_out <= 16'hf309;
             14'h32fb 	:	val_out <= 16'hf30b;
             14'h32fc 	:	val_out <= 16'hf30d;
             14'h32fd 	:	val_out <= 16'hf30f;
             14'h32fe 	:	val_out <= 16'hf311;
             14'h32ff 	:	val_out <= 16'hf313;
             14'h3300 	:	val_out <= 16'hf315;
             14'h3301 	:	val_out <= 16'hf317;
             14'h3302 	:	val_out <= 16'hf319;
             14'h3303 	:	val_out <= 16'hf31b;
             14'h3304 	:	val_out <= 16'hf31d;
             14'h3305 	:	val_out <= 16'hf31f;
             14'h3306 	:	val_out <= 16'hf321;
             14'h3307 	:	val_out <= 16'hf323;
             14'h3308 	:	val_out <= 16'hf325;
             14'h3309 	:	val_out <= 16'hf326;
             14'h330a 	:	val_out <= 16'hf328;
             14'h330b 	:	val_out <= 16'hf32a;
             14'h330c 	:	val_out <= 16'hf32c;
             14'h330d 	:	val_out <= 16'hf32e;
             14'h330e 	:	val_out <= 16'hf330;
             14'h330f 	:	val_out <= 16'hf332;
             14'h3310 	:	val_out <= 16'hf334;
             14'h3311 	:	val_out <= 16'hf336;
             14'h3312 	:	val_out <= 16'hf338;
             14'h3313 	:	val_out <= 16'hf33a;
             14'h3314 	:	val_out <= 16'hf33c;
             14'h3315 	:	val_out <= 16'hf33e;
             14'h3316 	:	val_out <= 16'hf340;
             14'h3317 	:	val_out <= 16'hf342;
             14'h3318 	:	val_out <= 16'hf344;
             14'h3319 	:	val_out <= 16'hf346;
             14'h331a 	:	val_out <= 16'hf348;
             14'h331b 	:	val_out <= 16'hf34a;
             14'h331c 	:	val_out <= 16'hf34c;
             14'h331d 	:	val_out <= 16'hf34e;
             14'h331e 	:	val_out <= 16'hf350;
             14'h331f 	:	val_out <= 16'hf352;
             14'h3320 	:	val_out <= 16'hf354;
             14'h3321 	:	val_out <= 16'hf355;
             14'h3322 	:	val_out <= 16'hf357;
             14'h3323 	:	val_out <= 16'hf359;
             14'h3324 	:	val_out <= 16'hf35b;
             14'h3325 	:	val_out <= 16'hf35d;
             14'h3326 	:	val_out <= 16'hf35f;
             14'h3327 	:	val_out <= 16'hf361;
             14'h3328 	:	val_out <= 16'hf363;
             14'h3329 	:	val_out <= 16'hf365;
             14'h332a 	:	val_out <= 16'hf367;
             14'h332b 	:	val_out <= 16'hf369;
             14'h332c 	:	val_out <= 16'hf36b;
             14'h332d 	:	val_out <= 16'hf36d;
             14'h332e 	:	val_out <= 16'hf36f;
             14'h332f 	:	val_out <= 16'hf371;
             14'h3330 	:	val_out <= 16'hf373;
             14'h3331 	:	val_out <= 16'hf375;
             14'h3332 	:	val_out <= 16'hf377;
             14'h3333 	:	val_out <= 16'hf379;
             14'h3334 	:	val_out <= 16'hf37a;
             14'h3335 	:	val_out <= 16'hf37c;
             14'h3336 	:	val_out <= 16'hf37e;
             14'h3337 	:	val_out <= 16'hf380;
             14'h3338 	:	val_out <= 16'hf382;
             14'h3339 	:	val_out <= 16'hf384;
             14'h333a 	:	val_out <= 16'hf386;
             14'h333b 	:	val_out <= 16'hf388;
             14'h333c 	:	val_out <= 16'hf38a;
             14'h333d 	:	val_out <= 16'hf38c;
             14'h333e 	:	val_out <= 16'hf38e;
             14'h333f 	:	val_out <= 16'hf390;
             14'h3340 	:	val_out <= 16'hf392;
             14'h3341 	:	val_out <= 16'hf394;
             14'h3342 	:	val_out <= 16'hf396;
             14'h3343 	:	val_out <= 16'hf398;
             14'h3344 	:	val_out <= 16'hf399;
             14'h3345 	:	val_out <= 16'hf39b;
             14'h3346 	:	val_out <= 16'hf39d;
             14'h3347 	:	val_out <= 16'hf39f;
             14'h3348 	:	val_out <= 16'hf3a1;
             14'h3349 	:	val_out <= 16'hf3a3;
             14'h334a 	:	val_out <= 16'hf3a5;
             14'h334b 	:	val_out <= 16'hf3a7;
             14'h334c 	:	val_out <= 16'hf3a9;
             14'h334d 	:	val_out <= 16'hf3ab;
             14'h334e 	:	val_out <= 16'hf3ad;
             14'h334f 	:	val_out <= 16'hf3af;
             14'h3350 	:	val_out <= 16'hf3b1;
             14'h3351 	:	val_out <= 16'hf3b3;
             14'h3352 	:	val_out <= 16'hf3b4;
             14'h3353 	:	val_out <= 16'hf3b6;
             14'h3354 	:	val_out <= 16'hf3b8;
             14'h3355 	:	val_out <= 16'hf3ba;
             14'h3356 	:	val_out <= 16'hf3bc;
             14'h3357 	:	val_out <= 16'hf3be;
             14'h3358 	:	val_out <= 16'hf3c0;
             14'h3359 	:	val_out <= 16'hf3c2;
             14'h335a 	:	val_out <= 16'hf3c4;
             14'h335b 	:	val_out <= 16'hf3c6;
             14'h335c 	:	val_out <= 16'hf3c8;
             14'h335d 	:	val_out <= 16'hf3ca;
             14'h335e 	:	val_out <= 16'hf3cb;
             14'h335f 	:	val_out <= 16'hf3cd;
             14'h3360 	:	val_out <= 16'hf3cf;
             14'h3361 	:	val_out <= 16'hf3d1;
             14'h3362 	:	val_out <= 16'hf3d3;
             14'h3363 	:	val_out <= 16'hf3d5;
             14'h3364 	:	val_out <= 16'hf3d7;
             14'h3365 	:	val_out <= 16'hf3d9;
             14'h3366 	:	val_out <= 16'hf3db;
             14'h3367 	:	val_out <= 16'hf3dd;
             14'h3368 	:	val_out <= 16'hf3df;
             14'h3369 	:	val_out <= 16'hf3e1;
             14'h336a 	:	val_out <= 16'hf3e2;
             14'h336b 	:	val_out <= 16'hf3e4;
             14'h336c 	:	val_out <= 16'hf3e6;
             14'h336d 	:	val_out <= 16'hf3e8;
             14'h336e 	:	val_out <= 16'hf3ea;
             14'h336f 	:	val_out <= 16'hf3ec;
             14'h3370 	:	val_out <= 16'hf3ee;
             14'h3371 	:	val_out <= 16'hf3f0;
             14'h3372 	:	val_out <= 16'hf3f2;
             14'h3373 	:	val_out <= 16'hf3f4;
             14'h3374 	:	val_out <= 16'hf3f6;
             14'h3375 	:	val_out <= 16'hf3f7;
             14'h3376 	:	val_out <= 16'hf3f9;
             14'h3377 	:	val_out <= 16'hf3fb;
             14'h3378 	:	val_out <= 16'hf3fd;
             14'h3379 	:	val_out <= 16'hf3ff;
             14'h337a 	:	val_out <= 16'hf401;
             14'h337b 	:	val_out <= 16'hf403;
             14'h337c 	:	val_out <= 16'hf405;
             14'h337d 	:	val_out <= 16'hf407;
             14'h337e 	:	val_out <= 16'hf409;
             14'h337f 	:	val_out <= 16'hf40a;
             14'h3380 	:	val_out <= 16'hf40c;
             14'h3381 	:	val_out <= 16'hf40e;
             14'h3382 	:	val_out <= 16'hf410;
             14'h3383 	:	val_out <= 16'hf412;
             14'h3384 	:	val_out <= 16'hf414;
             14'h3385 	:	val_out <= 16'hf416;
             14'h3386 	:	val_out <= 16'hf418;
             14'h3387 	:	val_out <= 16'hf41a;
             14'h3388 	:	val_out <= 16'hf41b;
             14'h3389 	:	val_out <= 16'hf41d;
             14'h338a 	:	val_out <= 16'hf41f;
             14'h338b 	:	val_out <= 16'hf421;
             14'h338c 	:	val_out <= 16'hf423;
             14'h338d 	:	val_out <= 16'hf425;
             14'h338e 	:	val_out <= 16'hf427;
             14'h338f 	:	val_out <= 16'hf429;
             14'h3390 	:	val_out <= 16'hf42b;
             14'h3391 	:	val_out <= 16'hf42c;
             14'h3392 	:	val_out <= 16'hf42e;
             14'h3393 	:	val_out <= 16'hf430;
             14'h3394 	:	val_out <= 16'hf432;
             14'h3395 	:	val_out <= 16'hf434;
             14'h3396 	:	val_out <= 16'hf436;
             14'h3397 	:	val_out <= 16'hf438;
             14'h3398 	:	val_out <= 16'hf43a;
             14'h3399 	:	val_out <= 16'hf43c;
             14'h339a 	:	val_out <= 16'hf43d;
             14'h339b 	:	val_out <= 16'hf43f;
             14'h339c 	:	val_out <= 16'hf441;
             14'h339d 	:	val_out <= 16'hf443;
             14'h339e 	:	val_out <= 16'hf445;
             14'h339f 	:	val_out <= 16'hf447;
             14'h33a0 	:	val_out <= 16'hf449;
             14'h33a1 	:	val_out <= 16'hf44b;
             14'h33a2 	:	val_out <= 16'hf44c;
             14'h33a3 	:	val_out <= 16'hf44e;
             14'h33a4 	:	val_out <= 16'hf450;
             14'h33a5 	:	val_out <= 16'hf452;
             14'h33a6 	:	val_out <= 16'hf454;
             14'h33a7 	:	val_out <= 16'hf456;
             14'h33a8 	:	val_out <= 16'hf458;
             14'h33a9 	:	val_out <= 16'hf45a;
             14'h33aa 	:	val_out <= 16'hf45b;
             14'h33ab 	:	val_out <= 16'hf45d;
             14'h33ac 	:	val_out <= 16'hf45f;
             14'h33ad 	:	val_out <= 16'hf461;
             14'h33ae 	:	val_out <= 16'hf463;
             14'h33af 	:	val_out <= 16'hf465;
             14'h33b0 	:	val_out <= 16'hf467;
             14'h33b1 	:	val_out <= 16'hf469;
             14'h33b2 	:	val_out <= 16'hf46a;
             14'h33b3 	:	val_out <= 16'hf46c;
             14'h33b4 	:	val_out <= 16'hf46e;
             14'h33b5 	:	val_out <= 16'hf470;
             14'h33b6 	:	val_out <= 16'hf472;
             14'h33b7 	:	val_out <= 16'hf474;
             14'h33b8 	:	val_out <= 16'hf476;
             14'h33b9 	:	val_out <= 16'hf478;
             14'h33ba 	:	val_out <= 16'hf479;
             14'h33bb 	:	val_out <= 16'hf47b;
             14'h33bc 	:	val_out <= 16'hf47d;
             14'h33bd 	:	val_out <= 16'hf47f;
             14'h33be 	:	val_out <= 16'hf481;
             14'h33bf 	:	val_out <= 16'hf483;
             14'h33c0 	:	val_out <= 16'hf485;
             14'h33c1 	:	val_out <= 16'hf486;
             14'h33c2 	:	val_out <= 16'hf488;
             14'h33c3 	:	val_out <= 16'hf48a;
             14'h33c4 	:	val_out <= 16'hf48c;
             14'h33c5 	:	val_out <= 16'hf48e;
             14'h33c6 	:	val_out <= 16'hf490;
             14'h33c7 	:	val_out <= 16'hf492;
             14'h33c8 	:	val_out <= 16'hf493;
             14'h33c9 	:	val_out <= 16'hf495;
             14'h33ca 	:	val_out <= 16'hf497;
             14'h33cb 	:	val_out <= 16'hf499;
             14'h33cc 	:	val_out <= 16'hf49b;
             14'h33cd 	:	val_out <= 16'hf49d;
             14'h33ce 	:	val_out <= 16'hf49f;
             14'h33cf 	:	val_out <= 16'hf4a0;
             14'h33d0 	:	val_out <= 16'hf4a2;
             14'h33d1 	:	val_out <= 16'hf4a4;
             14'h33d2 	:	val_out <= 16'hf4a6;
             14'h33d3 	:	val_out <= 16'hf4a8;
             14'h33d4 	:	val_out <= 16'hf4aa;
             14'h33d5 	:	val_out <= 16'hf4ac;
             14'h33d6 	:	val_out <= 16'hf4ad;
             14'h33d7 	:	val_out <= 16'hf4af;
             14'h33d8 	:	val_out <= 16'hf4b1;
             14'h33d9 	:	val_out <= 16'hf4b3;
             14'h33da 	:	val_out <= 16'hf4b5;
             14'h33db 	:	val_out <= 16'hf4b7;
             14'h33dc 	:	val_out <= 16'hf4b8;
             14'h33dd 	:	val_out <= 16'hf4ba;
             14'h33de 	:	val_out <= 16'hf4bc;
             14'h33df 	:	val_out <= 16'hf4be;
             14'h33e0 	:	val_out <= 16'hf4c0;
             14'h33e1 	:	val_out <= 16'hf4c2;
             14'h33e2 	:	val_out <= 16'hf4c3;
             14'h33e3 	:	val_out <= 16'hf4c5;
             14'h33e4 	:	val_out <= 16'hf4c7;
             14'h33e5 	:	val_out <= 16'hf4c9;
             14'h33e6 	:	val_out <= 16'hf4cb;
             14'h33e7 	:	val_out <= 16'hf4cd;
             14'h33e8 	:	val_out <= 16'hf4cf;
             14'h33e9 	:	val_out <= 16'hf4d0;
             14'h33ea 	:	val_out <= 16'hf4d2;
             14'h33eb 	:	val_out <= 16'hf4d4;
             14'h33ec 	:	val_out <= 16'hf4d6;
             14'h33ed 	:	val_out <= 16'hf4d8;
             14'h33ee 	:	val_out <= 16'hf4da;
             14'h33ef 	:	val_out <= 16'hf4db;
             14'h33f0 	:	val_out <= 16'hf4dd;
             14'h33f1 	:	val_out <= 16'hf4df;
             14'h33f2 	:	val_out <= 16'hf4e1;
             14'h33f3 	:	val_out <= 16'hf4e3;
             14'h33f4 	:	val_out <= 16'hf4e5;
             14'h33f5 	:	val_out <= 16'hf4e6;
             14'h33f6 	:	val_out <= 16'hf4e8;
             14'h33f7 	:	val_out <= 16'hf4ea;
             14'h33f8 	:	val_out <= 16'hf4ec;
             14'h33f9 	:	val_out <= 16'hf4ee;
             14'h33fa 	:	val_out <= 16'hf4f0;
             14'h33fb 	:	val_out <= 16'hf4f1;
             14'h33fc 	:	val_out <= 16'hf4f3;
             14'h33fd 	:	val_out <= 16'hf4f5;
             14'h33fe 	:	val_out <= 16'hf4f7;
             14'h33ff 	:	val_out <= 16'hf4f9;
             14'h3400 	:	val_out <= 16'hf4fa;
             14'h3401 	:	val_out <= 16'hf4fc;
             14'h3402 	:	val_out <= 16'hf4fe;
             14'h3403 	:	val_out <= 16'hf500;
             14'h3404 	:	val_out <= 16'hf502;
             14'h3405 	:	val_out <= 16'hf504;
             14'h3406 	:	val_out <= 16'hf505;
             14'h3407 	:	val_out <= 16'hf507;
             14'h3408 	:	val_out <= 16'hf509;
             14'h3409 	:	val_out <= 16'hf50b;
             14'h340a 	:	val_out <= 16'hf50d;
             14'h340b 	:	val_out <= 16'hf50e;
             14'h340c 	:	val_out <= 16'hf510;
             14'h340d 	:	val_out <= 16'hf512;
             14'h340e 	:	val_out <= 16'hf514;
             14'h340f 	:	val_out <= 16'hf516;
             14'h3410 	:	val_out <= 16'hf518;
             14'h3411 	:	val_out <= 16'hf519;
             14'h3412 	:	val_out <= 16'hf51b;
             14'h3413 	:	val_out <= 16'hf51d;
             14'h3414 	:	val_out <= 16'hf51f;
             14'h3415 	:	val_out <= 16'hf521;
             14'h3416 	:	val_out <= 16'hf522;
             14'h3417 	:	val_out <= 16'hf524;
             14'h3418 	:	val_out <= 16'hf526;
             14'h3419 	:	val_out <= 16'hf528;
             14'h341a 	:	val_out <= 16'hf52a;
             14'h341b 	:	val_out <= 16'hf52b;
             14'h341c 	:	val_out <= 16'hf52d;
             14'h341d 	:	val_out <= 16'hf52f;
             14'h341e 	:	val_out <= 16'hf531;
             14'h341f 	:	val_out <= 16'hf533;
             14'h3420 	:	val_out <= 16'hf535;
             14'h3421 	:	val_out <= 16'hf536;
             14'h3422 	:	val_out <= 16'hf538;
             14'h3423 	:	val_out <= 16'hf53a;
             14'h3424 	:	val_out <= 16'hf53c;
             14'h3425 	:	val_out <= 16'hf53e;
             14'h3426 	:	val_out <= 16'hf53f;
             14'h3427 	:	val_out <= 16'hf541;
             14'h3428 	:	val_out <= 16'hf543;
             14'h3429 	:	val_out <= 16'hf545;
             14'h342a 	:	val_out <= 16'hf547;
             14'h342b 	:	val_out <= 16'hf548;
             14'h342c 	:	val_out <= 16'hf54a;
             14'h342d 	:	val_out <= 16'hf54c;
             14'h342e 	:	val_out <= 16'hf54e;
             14'h342f 	:	val_out <= 16'hf550;
             14'h3430 	:	val_out <= 16'hf551;
             14'h3431 	:	val_out <= 16'hf553;
             14'h3432 	:	val_out <= 16'hf555;
             14'h3433 	:	val_out <= 16'hf557;
             14'h3434 	:	val_out <= 16'hf559;
             14'h3435 	:	val_out <= 16'hf55a;
             14'h3436 	:	val_out <= 16'hf55c;
             14'h3437 	:	val_out <= 16'hf55e;
             14'h3438 	:	val_out <= 16'hf560;
             14'h3439 	:	val_out <= 16'hf561;
             14'h343a 	:	val_out <= 16'hf563;
             14'h343b 	:	val_out <= 16'hf565;
             14'h343c 	:	val_out <= 16'hf567;
             14'h343d 	:	val_out <= 16'hf569;
             14'h343e 	:	val_out <= 16'hf56a;
             14'h343f 	:	val_out <= 16'hf56c;
             14'h3440 	:	val_out <= 16'hf56e;
             14'h3441 	:	val_out <= 16'hf570;
             14'h3442 	:	val_out <= 16'hf572;
             14'h3443 	:	val_out <= 16'hf573;
             14'h3444 	:	val_out <= 16'hf575;
             14'h3445 	:	val_out <= 16'hf577;
             14'h3446 	:	val_out <= 16'hf579;
             14'h3447 	:	val_out <= 16'hf57a;
             14'h3448 	:	val_out <= 16'hf57c;
             14'h3449 	:	val_out <= 16'hf57e;
             14'h344a 	:	val_out <= 16'hf580;
             14'h344b 	:	val_out <= 16'hf582;
             14'h344c 	:	val_out <= 16'hf583;
             14'h344d 	:	val_out <= 16'hf585;
             14'h344e 	:	val_out <= 16'hf587;
             14'h344f 	:	val_out <= 16'hf589;
             14'h3450 	:	val_out <= 16'hf58a;
             14'h3451 	:	val_out <= 16'hf58c;
             14'h3452 	:	val_out <= 16'hf58e;
             14'h3453 	:	val_out <= 16'hf590;
             14'h3454 	:	val_out <= 16'hf592;
             14'h3455 	:	val_out <= 16'hf593;
             14'h3456 	:	val_out <= 16'hf595;
             14'h3457 	:	val_out <= 16'hf597;
             14'h3458 	:	val_out <= 16'hf599;
             14'h3459 	:	val_out <= 16'hf59a;
             14'h345a 	:	val_out <= 16'hf59c;
             14'h345b 	:	val_out <= 16'hf59e;
             14'h345c 	:	val_out <= 16'hf5a0;
             14'h345d 	:	val_out <= 16'hf5a2;
             14'h345e 	:	val_out <= 16'hf5a3;
             14'h345f 	:	val_out <= 16'hf5a5;
             14'h3460 	:	val_out <= 16'hf5a7;
             14'h3461 	:	val_out <= 16'hf5a9;
             14'h3462 	:	val_out <= 16'hf5aa;
             14'h3463 	:	val_out <= 16'hf5ac;
             14'h3464 	:	val_out <= 16'hf5ae;
             14'h3465 	:	val_out <= 16'hf5b0;
             14'h3466 	:	val_out <= 16'hf5b1;
             14'h3467 	:	val_out <= 16'hf5b3;
             14'h3468 	:	val_out <= 16'hf5b5;
             14'h3469 	:	val_out <= 16'hf5b7;
             14'h346a 	:	val_out <= 16'hf5b9;
             14'h346b 	:	val_out <= 16'hf5ba;
             14'h346c 	:	val_out <= 16'hf5bc;
             14'h346d 	:	val_out <= 16'hf5be;
             14'h346e 	:	val_out <= 16'hf5c0;
             14'h346f 	:	val_out <= 16'hf5c1;
             14'h3470 	:	val_out <= 16'hf5c3;
             14'h3471 	:	val_out <= 16'hf5c5;
             14'h3472 	:	val_out <= 16'hf5c7;
             14'h3473 	:	val_out <= 16'hf5c8;
             14'h3474 	:	val_out <= 16'hf5ca;
             14'h3475 	:	val_out <= 16'hf5cc;
             14'h3476 	:	val_out <= 16'hf5ce;
             14'h3477 	:	val_out <= 16'hf5cf;
             14'h3478 	:	val_out <= 16'hf5d1;
             14'h3479 	:	val_out <= 16'hf5d3;
             14'h347a 	:	val_out <= 16'hf5d5;
             14'h347b 	:	val_out <= 16'hf5d6;
             14'h347c 	:	val_out <= 16'hf5d8;
             14'h347d 	:	val_out <= 16'hf5da;
             14'h347e 	:	val_out <= 16'hf5dc;
             14'h347f 	:	val_out <= 16'hf5dd;
             14'h3480 	:	val_out <= 16'hf5df;
             14'h3481 	:	val_out <= 16'hf5e1;
             14'h3482 	:	val_out <= 16'hf5e3;
             14'h3483 	:	val_out <= 16'hf5e4;
             14'h3484 	:	val_out <= 16'hf5e6;
             14'h3485 	:	val_out <= 16'hf5e8;
             14'h3486 	:	val_out <= 16'hf5ea;
             14'h3487 	:	val_out <= 16'hf5eb;
             14'h3488 	:	val_out <= 16'hf5ed;
             14'h3489 	:	val_out <= 16'hf5ef;
             14'h348a 	:	val_out <= 16'hf5f1;
             14'h348b 	:	val_out <= 16'hf5f2;
             14'h348c 	:	val_out <= 16'hf5f4;
             14'h348d 	:	val_out <= 16'hf5f6;
             14'h348e 	:	val_out <= 16'hf5f8;
             14'h348f 	:	val_out <= 16'hf5f9;
             14'h3490 	:	val_out <= 16'hf5fb;
             14'h3491 	:	val_out <= 16'hf5fd;
             14'h3492 	:	val_out <= 16'hf5ff;
             14'h3493 	:	val_out <= 16'hf600;
             14'h3494 	:	val_out <= 16'hf602;
             14'h3495 	:	val_out <= 16'hf604;
             14'h3496 	:	val_out <= 16'hf606;
             14'h3497 	:	val_out <= 16'hf607;
             14'h3498 	:	val_out <= 16'hf609;
             14'h3499 	:	val_out <= 16'hf60b;
             14'h349a 	:	val_out <= 16'hf60c;
             14'h349b 	:	val_out <= 16'hf60e;
             14'h349c 	:	val_out <= 16'hf610;
             14'h349d 	:	val_out <= 16'hf612;
             14'h349e 	:	val_out <= 16'hf613;
             14'h349f 	:	val_out <= 16'hf615;
             14'h34a0 	:	val_out <= 16'hf617;
             14'h34a1 	:	val_out <= 16'hf619;
             14'h34a2 	:	val_out <= 16'hf61a;
             14'h34a3 	:	val_out <= 16'hf61c;
             14'h34a4 	:	val_out <= 16'hf61e;
             14'h34a5 	:	val_out <= 16'hf61f;
             14'h34a6 	:	val_out <= 16'hf621;
             14'h34a7 	:	val_out <= 16'hf623;
             14'h34a8 	:	val_out <= 16'hf625;
             14'h34a9 	:	val_out <= 16'hf626;
             14'h34aa 	:	val_out <= 16'hf628;
             14'h34ab 	:	val_out <= 16'hf62a;
             14'h34ac 	:	val_out <= 16'hf62c;
             14'h34ad 	:	val_out <= 16'hf62d;
             14'h34ae 	:	val_out <= 16'hf62f;
             14'h34af 	:	val_out <= 16'hf631;
             14'h34b0 	:	val_out <= 16'hf632;
             14'h34b1 	:	val_out <= 16'hf634;
             14'h34b2 	:	val_out <= 16'hf636;
             14'h34b3 	:	val_out <= 16'hf638;
             14'h34b4 	:	val_out <= 16'hf639;
             14'h34b5 	:	val_out <= 16'hf63b;
             14'h34b6 	:	val_out <= 16'hf63d;
             14'h34b7 	:	val_out <= 16'hf63f;
             14'h34b8 	:	val_out <= 16'hf640;
             14'h34b9 	:	val_out <= 16'hf642;
             14'h34ba 	:	val_out <= 16'hf644;
             14'h34bb 	:	val_out <= 16'hf645;
             14'h34bc 	:	val_out <= 16'hf647;
             14'h34bd 	:	val_out <= 16'hf649;
             14'h34be 	:	val_out <= 16'hf64b;
             14'h34bf 	:	val_out <= 16'hf64c;
             14'h34c0 	:	val_out <= 16'hf64e;
             14'h34c1 	:	val_out <= 16'hf650;
             14'h34c2 	:	val_out <= 16'hf651;
             14'h34c3 	:	val_out <= 16'hf653;
             14'h34c4 	:	val_out <= 16'hf655;
             14'h34c5 	:	val_out <= 16'hf657;
             14'h34c6 	:	val_out <= 16'hf658;
             14'h34c7 	:	val_out <= 16'hf65a;
             14'h34c8 	:	val_out <= 16'hf65c;
             14'h34c9 	:	val_out <= 16'hf65d;
             14'h34ca 	:	val_out <= 16'hf65f;
             14'h34cb 	:	val_out <= 16'hf661;
             14'h34cc 	:	val_out <= 16'hf662;
             14'h34cd 	:	val_out <= 16'hf664;
             14'h34ce 	:	val_out <= 16'hf666;
             14'h34cf 	:	val_out <= 16'hf668;
             14'h34d0 	:	val_out <= 16'hf669;
             14'h34d1 	:	val_out <= 16'hf66b;
             14'h34d2 	:	val_out <= 16'hf66d;
             14'h34d3 	:	val_out <= 16'hf66e;
             14'h34d4 	:	val_out <= 16'hf670;
             14'h34d5 	:	val_out <= 16'hf672;
             14'h34d6 	:	val_out <= 16'hf673;
             14'h34d7 	:	val_out <= 16'hf675;
             14'h34d8 	:	val_out <= 16'hf677;
             14'h34d9 	:	val_out <= 16'hf679;
             14'h34da 	:	val_out <= 16'hf67a;
             14'h34db 	:	val_out <= 16'hf67c;
             14'h34dc 	:	val_out <= 16'hf67e;
             14'h34dd 	:	val_out <= 16'hf67f;
             14'h34de 	:	val_out <= 16'hf681;
             14'h34df 	:	val_out <= 16'hf683;
             14'h34e0 	:	val_out <= 16'hf684;
             14'h34e1 	:	val_out <= 16'hf686;
             14'h34e2 	:	val_out <= 16'hf688;
             14'h34e3 	:	val_out <= 16'hf68a;
             14'h34e4 	:	val_out <= 16'hf68b;
             14'h34e5 	:	val_out <= 16'hf68d;
             14'h34e6 	:	val_out <= 16'hf68f;
             14'h34e7 	:	val_out <= 16'hf690;
             14'h34e8 	:	val_out <= 16'hf692;
             14'h34e9 	:	val_out <= 16'hf694;
             14'h34ea 	:	val_out <= 16'hf695;
             14'h34eb 	:	val_out <= 16'hf697;
             14'h34ec 	:	val_out <= 16'hf699;
             14'h34ed 	:	val_out <= 16'hf69a;
             14'h34ee 	:	val_out <= 16'hf69c;
             14'h34ef 	:	val_out <= 16'hf69e;
             14'h34f0 	:	val_out <= 16'hf69f;
             14'h34f1 	:	val_out <= 16'hf6a1;
             14'h34f2 	:	val_out <= 16'hf6a3;
             14'h34f3 	:	val_out <= 16'hf6a5;
             14'h34f4 	:	val_out <= 16'hf6a6;
             14'h34f5 	:	val_out <= 16'hf6a8;
             14'h34f6 	:	val_out <= 16'hf6aa;
             14'h34f7 	:	val_out <= 16'hf6ab;
             14'h34f8 	:	val_out <= 16'hf6ad;
             14'h34f9 	:	val_out <= 16'hf6af;
             14'h34fa 	:	val_out <= 16'hf6b0;
             14'h34fb 	:	val_out <= 16'hf6b2;
             14'h34fc 	:	val_out <= 16'hf6b4;
             14'h34fd 	:	val_out <= 16'hf6b5;
             14'h34fe 	:	val_out <= 16'hf6b7;
             14'h34ff 	:	val_out <= 16'hf6b9;
             14'h3500 	:	val_out <= 16'hf6ba;
             14'h3501 	:	val_out <= 16'hf6bc;
             14'h3502 	:	val_out <= 16'hf6be;
             14'h3503 	:	val_out <= 16'hf6bf;
             14'h3504 	:	val_out <= 16'hf6c1;
             14'h3505 	:	val_out <= 16'hf6c3;
             14'h3506 	:	val_out <= 16'hf6c4;
             14'h3507 	:	val_out <= 16'hf6c6;
             14'h3508 	:	val_out <= 16'hf6c8;
             14'h3509 	:	val_out <= 16'hf6c9;
             14'h350a 	:	val_out <= 16'hf6cb;
             14'h350b 	:	val_out <= 16'hf6cd;
             14'h350c 	:	val_out <= 16'hf6ce;
             14'h350d 	:	val_out <= 16'hf6d0;
             14'h350e 	:	val_out <= 16'hf6d2;
             14'h350f 	:	val_out <= 16'hf6d3;
             14'h3510 	:	val_out <= 16'hf6d5;
             14'h3511 	:	val_out <= 16'hf6d7;
             14'h3512 	:	val_out <= 16'hf6d8;
             14'h3513 	:	val_out <= 16'hf6da;
             14'h3514 	:	val_out <= 16'hf6dc;
             14'h3515 	:	val_out <= 16'hf6dd;
             14'h3516 	:	val_out <= 16'hf6df;
             14'h3517 	:	val_out <= 16'hf6e1;
             14'h3518 	:	val_out <= 16'hf6e2;
             14'h3519 	:	val_out <= 16'hf6e4;
             14'h351a 	:	val_out <= 16'hf6e6;
             14'h351b 	:	val_out <= 16'hf6e7;
             14'h351c 	:	val_out <= 16'hf6e9;
             14'h351d 	:	val_out <= 16'hf6eb;
             14'h351e 	:	val_out <= 16'hf6ec;
             14'h351f 	:	val_out <= 16'hf6ee;
             14'h3520 	:	val_out <= 16'hf6f0;
             14'h3521 	:	val_out <= 16'hf6f1;
             14'h3522 	:	val_out <= 16'hf6f3;
             14'h3523 	:	val_out <= 16'hf6f5;
             14'h3524 	:	val_out <= 16'hf6f6;
             14'h3525 	:	val_out <= 16'hf6f8;
             14'h3526 	:	val_out <= 16'hf6fa;
             14'h3527 	:	val_out <= 16'hf6fb;
             14'h3528 	:	val_out <= 16'hf6fd;
             14'h3529 	:	val_out <= 16'hf6ff;
             14'h352a 	:	val_out <= 16'hf700;
             14'h352b 	:	val_out <= 16'hf702;
             14'h352c 	:	val_out <= 16'hf704;
             14'h352d 	:	val_out <= 16'hf705;
             14'h352e 	:	val_out <= 16'hf707;
             14'h352f 	:	val_out <= 16'hf708;
             14'h3530 	:	val_out <= 16'hf70a;
             14'h3531 	:	val_out <= 16'hf70c;
             14'h3532 	:	val_out <= 16'hf70d;
             14'h3533 	:	val_out <= 16'hf70f;
             14'h3534 	:	val_out <= 16'hf711;
             14'h3535 	:	val_out <= 16'hf712;
             14'h3536 	:	val_out <= 16'hf714;
             14'h3537 	:	val_out <= 16'hf716;
             14'h3538 	:	val_out <= 16'hf717;
             14'h3539 	:	val_out <= 16'hf719;
             14'h353a 	:	val_out <= 16'hf71b;
             14'h353b 	:	val_out <= 16'hf71c;
             14'h353c 	:	val_out <= 16'hf71e;
             14'h353d 	:	val_out <= 16'hf71f;
             14'h353e 	:	val_out <= 16'hf721;
             14'h353f 	:	val_out <= 16'hf723;
             14'h3540 	:	val_out <= 16'hf724;
             14'h3541 	:	val_out <= 16'hf726;
             14'h3542 	:	val_out <= 16'hf728;
             14'h3543 	:	val_out <= 16'hf729;
             14'h3544 	:	val_out <= 16'hf72b;
             14'h3545 	:	val_out <= 16'hf72d;
             14'h3546 	:	val_out <= 16'hf72e;
             14'h3547 	:	val_out <= 16'hf730;
             14'h3548 	:	val_out <= 16'hf731;
             14'h3549 	:	val_out <= 16'hf733;
             14'h354a 	:	val_out <= 16'hf735;
             14'h354b 	:	val_out <= 16'hf736;
             14'h354c 	:	val_out <= 16'hf738;
             14'h354d 	:	val_out <= 16'hf73a;
             14'h354e 	:	val_out <= 16'hf73b;
             14'h354f 	:	val_out <= 16'hf73d;
             14'h3550 	:	val_out <= 16'hf73f;
             14'h3551 	:	val_out <= 16'hf740;
             14'h3552 	:	val_out <= 16'hf742;
             14'h3553 	:	val_out <= 16'hf743;
             14'h3554 	:	val_out <= 16'hf745;
             14'h3555 	:	val_out <= 16'hf747;
             14'h3556 	:	val_out <= 16'hf748;
             14'h3557 	:	val_out <= 16'hf74a;
             14'h3558 	:	val_out <= 16'hf74c;
             14'h3559 	:	val_out <= 16'hf74d;
             14'h355a 	:	val_out <= 16'hf74f;
             14'h355b 	:	val_out <= 16'hf750;
             14'h355c 	:	val_out <= 16'hf752;
             14'h355d 	:	val_out <= 16'hf754;
             14'h355e 	:	val_out <= 16'hf755;
             14'h355f 	:	val_out <= 16'hf757;
             14'h3560 	:	val_out <= 16'hf759;
             14'h3561 	:	val_out <= 16'hf75a;
             14'h3562 	:	val_out <= 16'hf75c;
             14'h3563 	:	val_out <= 16'hf75d;
             14'h3564 	:	val_out <= 16'hf75f;
             14'h3565 	:	val_out <= 16'hf761;
             14'h3566 	:	val_out <= 16'hf762;
             14'h3567 	:	val_out <= 16'hf764;
             14'h3568 	:	val_out <= 16'hf765;
             14'h3569 	:	val_out <= 16'hf767;
             14'h356a 	:	val_out <= 16'hf769;
             14'h356b 	:	val_out <= 16'hf76a;
             14'h356c 	:	val_out <= 16'hf76c;
             14'h356d 	:	val_out <= 16'hf76e;
             14'h356e 	:	val_out <= 16'hf76f;
             14'h356f 	:	val_out <= 16'hf771;
             14'h3570 	:	val_out <= 16'hf772;
             14'h3571 	:	val_out <= 16'hf774;
             14'h3572 	:	val_out <= 16'hf776;
             14'h3573 	:	val_out <= 16'hf777;
             14'h3574 	:	val_out <= 16'hf779;
             14'h3575 	:	val_out <= 16'hf77a;
             14'h3576 	:	val_out <= 16'hf77c;
             14'h3577 	:	val_out <= 16'hf77e;
             14'h3578 	:	val_out <= 16'hf77f;
             14'h3579 	:	val_out <= 16'hf781;
             14'h357a 	:	val_out <= 16'hf782;
             14'h357b 	:	val_out <= 16'hf784;
             14'h357c 	:	val_out <= 16'hf786;
             14'h357d 	:	val_out <= 16'hf787;
             14'h357e 	:	val_out <= 16'hf789;
             14'h357f 	:	val_out <= 16'hf78a;
             14'h3580 	:	val_out <= 16'hf78c;
             14'h3581 	:	val_out <= 16'hf78e;
             14'h3582 	:	val_out <= 16'hf78f;
             14'h3583 	:	val_out <= 16'hf791;
             14'h3584 	:	val_out <= 16'hf792;
             14'h3585 	:	val_out <= 16'hf794;
             14'h3586 	:	val_out <= 16'hf796;
             14'h3587 	:	val_out <= 16'hf797;
             14'h3588 	:	val_out <= 16'hf799;
             14'h3589 	:	val_out <= 16'hf79a;
             14'h358a 	:	val_out <= 16'hf79c;
             14'h358b 	:	val_out <= 16'hf79e;
             14'h358c 	:	val_out <= 16'hf79f;
             14'h358d 	:	val_out <= 16'hf7a1;
             14'h358e 	:	val_out <= 16'hf7a2;
             14'h358f 	:	val_out <= 16'hf7a4;
             14'h3590 	:	val_out <= 16'hf7a6;
             14'h3591 	:	val_out <= 16'hf7a7;
             14'h3592 	:	val_out <= 16'hf7a9;
             14'h3593 	:	val_out <= 16'hf7aa;
             14'h3594 	:	val_out <= 16'hf7ac;
             14'h3595 	:	val_out <= 16'hf7ae;
             14'h3596 	:	val_out <= 16'hf7af;
             14'h3597 	:	val_out <= 16'hf7b1;
             14'h3598 	:	val_out <= 16'hf7b2;
             14'h3599 	:	val_out <= 16'hf7b4;
             14'h359a 	:	val_out <= 16'hf7b6;
             14'h359b 	:	val_out <= 16'hf7b7;
             14'h359c 	:	val_out <= 16'hf7b9;
             14'h359d 	:	val_out <= 16'hf7ba;
             14'h359e 	:	val_out <= 16'hf7bc;
             14'h359f 	:	val_out <= 16'hf7bd;
             14'h35a0 	:	val_out <= 16'hf7bf;
             14'h35a1 	:	val_out <= 16'hf7c1;
             14'h35a2 	:	val_out <= 16'hf7c2;
             14'h35a3 	:	val_out <= 16'hf7c4;
             14'h35a4 	:	val_out <= 16'hf7c5;
             14'h35a5 	:	val_out <= 16'hf7c7;
             14'h35a6 	:	val_out <= 16'hf7c8;
             14'h35a7 	:	val_out <= 16'hf7ca;
             14'h35a8 	:	val_out <= 16'hf7cc;
             14'h35a9 	:	val_out <= 16'hf7cd;
             14'h35aa 	:	val_out <= 16'hf7cf;
             14'h35ab 	:	val_out <= 16'hf7d0;
             14'h35ac 	:	val_out <= 16'hf7d2;
             14'h35ad 	:	val_out <= 16'hf7d4;
             14'h35ae 	:	val_out <= 16'hf7d5;
             14'h35af 	:	val_out <= 16'hf7d7;
             14'h35b0 	:	val_out <= 16'hf7d8;
             14'h35b1 	:	val_out <= 16'hf7da;
             14'h35b2 	:	val_out <= 16'hf7db;
             14'h35b3 	:	val_out <= 16'hf7dd;
             14'h35b4 	:	val_out <= 16'hf7df;
             14'h35b5 	:	val_out <= 16'hf7e0;
             14'h35b6 	:	val_out <= 16'hf7e2;
             14'h35b7 	:	val_out <= 16'hf7e3;
             14'h35b8 	:	val_out <= 16'hf7e5;
             14'h35b9 	:	val_out <= 16'hf7e6;
             14'h35ba 	:	val_out <= 16'hf7e8;
             14'h35bb 	:	val_out <= 16'hf7ea;
             14'h35bc 	:	val_out <= 16'hf7eb;
             14'h35bd 	:	val_out <= 16'hf7ed;
             14'h35be 	:	val_out <= 16'hf7ee;
             14'h35bf 	:	val_out <= 16'hf7f0;
             14'h35c0 	:	val_out <= 16'hf7f1;
             14'h35c1 	:	val_out <= 16'hf7f3;
             14'h35c2 	:	val_out <= 16'hf7f4;
             14'h35c3 	:	val_out <= 16'hf7f6;
             14'h35c4 	:	val_out <= 16'hf7f8;
             14'h35c5 	:	val_out <= 16'hf7f9;
             14'h35c6 	:	val_out <= 16'hf7fb;
             14'h35c7 	:	val_out <= 16'hf7fc;
             14'h35c8 	:	val_out <= 16'hf7fe;
             14'h35c9 	:	val_out <= 16'hf7ff;
             14'h35ca 	:	val_out <= 16'hf801;
             14'h35cb 	:	val_out <= 16'hf803;
             14'h35cc 	:	val_out <= 16'hf804;
             14'h35cd 	:	val_out <= 16'hf806;
             14'h35ce 	:	val_out <= 16'hf807;
             14'h35cf 	:	val_out <= 16'hf809;
             14'h35d0 	:	val_out <= 16'hf80a;
             14'h35d1 	:	val_out <= 16'hf80c;
             14'h35d2 	:	val_out <= 16'hf80d;
             14'h35d3 	:	val_out <= 16'hf80f;
             14'h35d4 	:	val_out <= 16'hf811;
             14'h35d5 	:	val_out <= 16'hf812;
             14'h35d6 	:	val_out <= 16'hf814;
             14'h35d7 	:	val_out <= 16'hf815;
             14'h35d8 	:	val_out <= 16'hf817;
             14'h35d9 	:	val_out <= 16'hf818;
             14'h35da 	:	val_out <= 16'hf81a;
             14'h35db 	:	val_out <= 16'hf81b;
             14'h35dc 	:	val_out <= 16'hf81d;
             14'h35dd 	:	val_out <= 16'hf81e;
             14'h35de 	:	val_out <= 16'hf820;
             14'h35df 	:	val_out <= 16'hf822;
             14'h35e0 	:	val_out <= 16'hf823;
             14'h35e1 	:	val_out <= 16'hf825;
             14'h35e2 	:	val_out <= 16'hf826;
             14'h35e3 	:	val_out <= 16'hf828;
             14'h35e4 	:	val_out <= 16'hf829;
             14'h35e5 	:	val_out <= 16'hf82b;
             14'h35e6 	:	val_out <= 16'hf82c;
             14'h35e7 	:	val_out <= 16'hf82e;
             14'h35e8 	:	val_out <= 16'hf82f;
             14'h35e9 	:	val_out <= 16'hf831;
             14'h35ea 	:	val_out <= 16'hf833;
             14'h35eb 	:	val_out <= 16'hf834;
             14'h35ec 	:	val_out <= 16'hf836;
             14'h35ed 	:	val_out <= 16'hf837;
             14'h35ee 	:	val_out <= 16'hf839;
             14'h35ef 	:	val_out <= 16'hf83a;
             14'h35f0 	:	val_out <= 16'hf83c;
             14'h35f1 	:	val_out <= 16'hf83d;
             14'h35f2 	:	val_out <= 16'hf83f;
             14'h35f3 	:	val_out <= 16'hf840;
             14'h35f4 	:	val_out <= 16'hf842;
             14'h35f5 	:	val_out <= 16'hf843;
             14'h35f6 	:	val_out <= 16'hf845;
             14'h35f7 	:	val_out <= 16'hf846;
             14'h35f8 	:	val_out <= 16'hf848;
             14'h35f9 	:	val_out <= 16'hf84a;
             14'h35fa 	:	val_out <= 16'hf84b;
             14'h35fb 	:	val_out <= 16'hf84d;
             14'h35fc 	:	val_out <= 16'hf84e;
             14'h35fd 	:	val_out <= 16'hf850;
             14'h35fe 	:	val_out <= 16'hf851;
             14'h35ff 	:	val_out <= 16'hf853;
             14'h3600 	:	val_out <= 16'hf854;
             14'h3601 	:	val_out <= 16'hf856;
             14'h3602 	:	val_out <= 16'hf857;
             14'h3603 	:	val_out <= 16'hf859;
             14'h3604 	:	val_out <= 16'hf85a;
             14'h3605 	:	val_out <= 16'hf85c;
             14'h3606 	:	val_out <= 16'hf85d;
             14'h3607 	:	val_out <= 16'hf85f;
             14'h3608 	:	val_out <= 16'hf860;
             14'h3609 	:	val_out <= 16'hf862;
             14'h360a 	:	val_out <= 16'hf863;
             14'h360b 	:	val_out <= 16'hf865;
             14'h360c 	:	val_out <= 16'hf867;
             14'h360d 	:	val_out <= 16'hf868;
             14'h360e 	:	val_out <= 16'hf86a;
             14'h360f 	:	val_out <= 16'hf86b;
             14'h3610 	:	val_out <= 16'hf86d;
             14'h3611 	:	val_out <= 16'hf86e;
             14'h3612 	:	val_out <= 16'hf870;
             14'h3613 	:	val_out <= 16'hf871;
             14'h3614 	:	val_out <= 16'hf873;
             14'h3615 	:	val_out <= 16'hf874;
             14'h3616 	:	val_out <= 16'hf876;
             14'h3617 	:	val_out <= 16'hf877;
             14'h3618 	:	val_out <= 16'hf879;
             14'h3619 	:	val_out <= 16'hf87a;
             14'h361a 	:	val_out <= 16'hf87c;
             14'h361b 	:	val_out <= 16'hf87d;
             14'h361c 	:	val_out <= 16'hf87f;
             14'h361d 	:	val_out <= 16'hf880;
             14'h361e 	:	val_out <= 16'hf882;
             14'h361f 	:	val_out <= 16'hf883;
             14'h3620 	:	val_out <= 16'hf885;
             14'h3621 	:	val_out <= 16'hf886;
             14'h3622 	:	val_out <= 16'hf888;
             14'h3623 	:	val_out <= 16'hf889;
             14'h3624 	:	val_out <= 16'hf88b;
             14'h3625 	:	val_out <= 16'hf88c;
             14'h3626 	:	val_out <= 16'hf88e;
             14'h3627 	:	val_out <= 16'hf88f;
             14'h3628 	:	val_out <= 16'hf891;
             14'h3629 	:	val_out <= 16'hf892;
             14'h362a 	:	val_out <= 16'hf894;
             14'h362b 	:	val_out <= 16'hf895;
             14'h362c 	:	val_out <= 16'hf897;
             14'h362d 	:	val_out <= 16'hf898;
             14'h362e 	:	val_out <= 16'hf89a;
             14'h362f 	:	val_out <= 16'hf89b;
             14'h3630 	:	val_out <= 16'hf89d;
             14'h3631 	:	val_out <= 16'hf89e;
             14'h3632 	:	val_out <= 16'hf8a0;
             14'h3633 	:	val_out <= 16'hf8a1;
             14'h3634 	:	val_out <= 16'hf8a3;
             14'h3635 	:	val_out <= 16'hf8a4;
             14'h3636 	:	val_out <= 16'hf8a6;
             14'h3637 	:	val_out <= 16'hf8a7;
             14'h3638 	:	val_out <= 16'hf8a9;
             14'h3639 	:	val_out <= 16'hf8aa;
             14'h363a 	:	val_out <= 16'hf8ac;
             14'h363b 	:	val_out <= 16'hf8ad;
             14'h363c 	:	val_out <= 16'hf8af;
             14'h363d 	:	val_out <= 16'hf8b0;
             14'h363e 	:	val_out <= 16'hf8b2;
             14'h363f 	:	val_out <= 16'hf8b3;
             14'h3640 	:	val_out <= 16'hf8b5;
             14'h3641 	:	val_out <= 16'hf8b6;
             14'h3642 	:	val_out <= 16'hf8b8;
             14'h3643 	:	val_out <= 16'hf8b9;
             14'h3644 	:	val_out <= 16'hf8bb;
             14'h3645 	:	val_out <= 16'hf8bc;
             14'h3646 	:	val_out <= 16'hf8be;
             14'h3647 	:	val_out <= 16'hf8bf;
             14'h3648 	:	val_out <= 16'hf8c1;
             14'h3649 	:	val_out <= 16'hf8c2;
             14'h364a 	:	val_out <= 16'hf8c4;
             14'h364b 	:	val_out <= 16'hf8c5;
             14'h364c 	:	val_out <= 16'hf8c7;
             14'h364d 	:	val_out <= 16'hf8c8;
             14'h364e 	:	val_out <= 16'hf8ca;
             14'h364f 	:	val_out <= 16'hf8cb;
             14'h3650 	:	val_out <= 16'hf8cc;
             14'h3651 	:	val_out <= 16'hf8ce;
             14'h3652 	:	val_out <= 16'hf8cf;
             14'h3653 	:	val_out <= 16'hf8d1;
             14'h3654 	:	val_out <= 16'hf8d2;
             14'h3655 	:	val_out <= 16'hf8d4;
             14'h3656 	:	val_out <= 16'hf8d5;
             14'h3657 	:	val_out <= 16'hf8d7;
             14'h3658 	:	val_out <= 16'hf8d8;
             14'h3659 	:	val_out <= 16'hf8da;
             14'h365a 	:	val_out <= 16'hf8db;
             14'h365b 	:	val_out <= 16'hf8dd;
             14'h365c 	:	val_out <= 16'hf8de;
             14'h365d 	:	val_out <= 16'hf8e0;
             14'h365e 	:	val_out <= 16'hf8e1;
             14'h365f 	:	val_out <= 16'hf8e3;
             14'h3660 	:	val_out <= 16'hf8e4;
             14'h3661 	:	val_out <= 16'hf8e6;
             14'h3662 	:	val_out <= 16'hf8e7;
             14'h3663 	:	val_out <= 16'hf8e8;
             14'h3664 	:	val_out <= 16'hf8ea;
             14'h3665 	:	val_out <= 16'hf8eb;
             14'h3666 	:	val_out <= 16'hf8ed;
             14'h3667 	:	val_out <= 16'hf8ee;
             14'h3668 	:	val_out <= 16'hf8f0;
             14'h3669 	:	val_out <= 16'hf8f1;
             14'h366a 	:	val_out <= 16'hf8f3;
             14'h366b 	:	val_out <= 16'hf8f4;
             14'h366c 	:	val_out <= 16'hf8f6;
             14'h366d 	:	val_out <= 16'hf8f7;
             14'h366e 	:	val_out <= 16'hf8f9;
             14'h366f 	:	val_out <= 16'hf8fa;
             14'h3670 	:	val_out <= 16'hf8fc;
             14'h3671 	:	val_out <= 16'hf8fd;
             14'h3672 	:	val_out <= 16'hf8fe;
             14'h3673 	:	val_out <= 16'hf900;
             14'h3674 	:	val_out <= 16'hf901;
             14'h3675 	:	val_out <= 16'hf903;
             14'h3676 	:	val_out <= 16'hf904;
             14'h3677 	:	val_out <= 16'hf906;
             14'h3678 	:	val_out <= 16'hf907;
             14'h3679 	:	val_out <= 16'hf909;
             14'h367a 	:	val_out <= 16'hf90a;
             14'h367b 	:	val_out <= 16'hf90c;
             14'h367c 	:	val_out <= 16'hf90d;
             14'h367d 	:	val_out <= 16'hf90e;
             14'h367e 	:	val_out <= 16'hf910;
             14'h367f 	:	val_out <= 16'hf911;
             14'h3680 	:	val_out <= 16'hf913;
             14'h3681 	:	val_out <= 16'hf914;
             14'h3682 	:	val_out <= 16'hf916;
             14'h3683 	:	val_out <= 16'hf917;
             14'h3684 	:	val_out <= 16'hf919;
             14'h3685 	:	val_out <= 16'hf91a;
             14'h3686 	:	val_out <= 16'hf91c;
             14'h3687 	:	val_out <= 16'hf91d;
             14'h3688 	:	val_out <= 16'hf91e;
             14'h3689 	:	val_out <= 16'hf920;
             14'h368a 	:	val_out <= 16'hf921;
             14'h368b 	:	val_out <= 16'hf923;
             14'h368c 	:	val_out <= 16'hf924;
             14'h368d 	:	val_out <= 16'hf926;
             14'h368e 	:	val_out <= 16'hf927;
             14'h368f 	:	val_out <= 16'hf929;
             14'h3690 	:	val_out <= 16'hf92a;
             14'h3691 	:	val_out <= 16'hf92b;
             14'h3692 	:	val_out <= 16'hf92d;
             14'h3693 	:	val_out <= 16'hf92e;
             14'h3694 	:	val_out <= 16'hf930;
             14'h3695 	:	val_out <= 16'hf931;
             14'h3696 	:	val_out <= 16'hf933;
             14'h3697 	:	val_out <= 16'hf934;
             14'h3698 	:	val_out <= 16'hf935;
             14'h3699 	:	val_out <= 16'hf937;
             14'h369a 	:	val_out <= 16'hf938;
             14'h369b 	:	val_out <= 16'hf93a;
             14'h369c 	:	val_out <= 16'hf93b;
             14'h369d 	:	val_out <= 16'hf93d;
             14'h369e 	:	val_out <= 16'hf93e;
             14'h369f 	:	val_out <= 16'hf940;
             14'h36a0 	:	val_out <= 16'hf941;
             14'h36a1 	:	val_out <= 16'hf942;
             14'h36a2 	:	val_out <= 16'hf944;
             14'h36a3 	:	val_out <= 16'hf945;
             14'h36a4 	:	val_out <= 16'hf947;
             14'h36a5 	:	val_out <= 16'hf948;
             14'h36a6 	:	val_out <= 16'hf94a;
             14'h36a7 	:	val_out <= 16'hf94b;
             14'h36a8 	:	val_out <= 16'hf94c;
             14'h36a9 	:	val_out <= 16'hf94e;
             14'h36aa 	:	val_out <= 16'hf94f;
             14'h36ab 	:	val_out <= 16'hf951;
             14'h36ac 	:	val_out <= 16'hf952;
             14'h36ad 	:	val_out <= 16'hf954;
             14'h36ae 	:	val_out <= 16'hf955;
             14'h36af 	:	val_out <= 16'hf956;
             14'h36b0 	:	val_out <= 16'hf958;
             14'h36b1 	:	val_out <= 16'hf959;
             14'h36b2 	:	val_out <= 16'hf95b;
             14'h36b3 	:	val_out <= 16'hf95c;
             14'h36b4 	:	val_out <= 16'hf95e;
             14'h36b5 	:	val_out <= 16'hf95f;
             14'h36b6 	:	val_out <= 16'hf960;
             14'h36b7 	:	val_out <= 16'hf962;
             14'h36b8 	:	val_out <= 16'hf963;
             14'h36b9 	:	val_out <= 16'hf965;
             14'h36ba 	:	val_out <= 16'hf966;
             14'h36bb 	:	val_out <= 16'hf967;
             14'h36bc 	:	val_out <= 16'hf969;
             14'h36bd 	:	val_out <= 16'hf96a;
             14'h36be 	:	val_out <= 16'hf96c;
             14'h36bf 	:	val_out <= 16'hf96d;
             14'h36c0 	:	val_out <= 16'hf96f;
             14'h36c1 	:	val_out <= 16'hf970;
             14'h36c2 	:	val_out <= 16'hf971;
             14'h36c3 	:	val_out <= 16'hf973;
             14'h36c4 	:	val_out <= 16'hf974;
             14'h36c5 	:	val_out <= 16'hf976;
             14'h36c6 	:	val_out <= 16'hf977;
             14'h36c7 	:	val_out <= 16'hf978;
             14'h36c8 	:	val_out <= 16'hf97a;
             14'h36c9 	:	val_out <= 16'hf97b;
             14'h36ca 	:	val_out <= 16'hf97d;
             14'h36cb 	:	val_out <= 16'hf97e;
             14'h36cc 	:	val_out <= 16'hf97f;
             14'h36cd 	:	val_out <= 16'hf981;
             14'h36ce 	:	val_out <= 16'hf982;
             14'h36cf 	:	val_out <= 16'hf984;
             14'h36d0 	:	val_out <= 16'hf985;
             14'h36d1 	:	val_out <= 16'hf986;
             14'h36d2 	:	val_out <= 16'hf988;
             14'h36d3 	:	val_out <= 16'hf989;
             14'h36d4 	:	val_out <= 16'hf98b;
             14'h36d5 	:	val_out <= 16'hf98c;
             14'h36d6 	:	val_out <= 16'hf98d;
             14'h36d7 	:	val_out <= 16'hf98f;
             14'h36d8 	:	val_out <= 16'hf990;
             14'h36d9 	:	val_out <= 16'hf992;
             14'h36da 	:	val_out <= 16'hf993;
             14'h36db 	:	val_out <= 16'hf994;
             14'h36dc 	:	val_out <= 16'hf996;
             14'h36dd 	:	val_out <= 16'hf997;
             14'h36de 	:	val_out <= 16'hf999;
             14'h36df 	:	val_out <= 16'hf99a;
             14'h36e0 	:	val_out <= 16'hf99b;
             14'h36e1 	:	val_out <= 16'hf99d;
             14'h36e2 	:	val_out <= 16'hf99e;
             14'h36e3 	:	val_out <= 16'hf9a0;
             14'h36e4 	:	val_out <= 16'hf9a1;
             14'h36e5 	:	val_out <= 16'hf9a2;
             14'h36e6 	:	val_out <= 16'hf9a4;
             14'h36e7 	:	val_out <= 16'hf9a5;
             14'h36e8 	:	val_out <= 16'hf9a7;
             14'h36e9 	:	val_out <= 16'hf9a8;
             14'h36ea 	:	val_out <= 16'hf9a9;
             14'h36eb 	:	val_out <= 16'hf9ab;
             14'h36ec 	:	val_out <= 16'hf9ac;
             14'h36ed 	:	val_out <= 16'hf9ae;
             14'h36ee 	:	val_out <= 16'hf9af;
             14'h36ef 	:	val_out <= 16'hf9b0;
             14'h36f0 	:	val_out <= 16'hf9b2;
             14'h36f1 	:	val_out <= 16'hf9b3;
             14'h36f2 	:	val_out <= 16'hf9b4;
             14'h36f3 	:	val_out <= 16'hf9b6;
             14'h36f4 	:	val_out <= 16'hf9b7;
             14'h36f5 	:	val_out <= 16'hf9b9;
             14'h36f6 	:	val_out <= 16'hf9ba;
             14'h36f7 	:	val_out <= 16'hf9bb;
             14'h36f8 	:	val_out <= 16'hf9bd;
             14'h36f9 	:	val_out <= 16'hf9be;
             14'h36fa 	:	val_out <= 16'hf9c0;
             14'h36fb 	:	val_out <= 16'hf9c1;
             14'h36fc 	:	val_out <= 16'hf9c2;
             14'h36fd 	:	val_out <= 16'hf9c4;
             14'h36fe 	:	val_out <= 16'hf9c5;
             14'h36ff 	:	val_out <= 16'hf9c6;
             14'h3700 	:	val_out <= 16'hf9c8;
             14'h3701 	:	val_out <= 16'hf9c9;
             14'h3702 	:	val_out <= 16'hf9cb;
             14'h3703 	:	val_out <= 16'hf9cc;
             14'h3704 	:	val_out <= 16'hf9cd;
             14'h3705 	:	val_out <= 16'hf9cf;
             14'h3706 	:	val_out <= 16'hf9d0;
             14'h3707 	:	val_out <= 16'hf9d1;
             14'h3708 	:	val_out <= 16'hf9d3;
             14'h3709 	:	val_out <= 16'hf9d4;
             14'h370a 	:	val_out <= 16'hf9d6;
             14'h370b 	:	val_out <= 16'hf9d7;
             14'h370c 	:	val_out <= 16'hf9d8;
             14'h370d 	:	val_out <= 16'hf9da;
             14'h370e 	:	val_out <= 16'hf9db;
             14'h370f 	:	val_out <= 16'hf9dc;
             14'h3710 	:	val_out <= 16'hf9de;
             14'h3711 	:	val_out <= 16'hf9df;
             14'h3712 	:	val_out <= 16'hf9e0;
             14'h3713 	:	val_out <= 16'hf9e2;
             14'h3714 	:	val_out <= 16'hf9e3;
             14'h3715 	:	val_out <= 16'hf9e5;
             14'h3716 	:	val_out <= 16'hf9e6;
             14'h3717 	:	val_out <= 16'hf9e7;
             14'h3718 	:	val_out <= 16'hf9e9;
             14'h3719 	:	val_out <= 16'hf9ea;
             14'h371a 	:	val_out <= 16'hf9eb;
             14'h371b 	:	val_out <= 16'hf9ed;
             14'h371c 	:	val_out <= 16'hf9ee;
             14'h371d 	:	val_out <= 16'hf9ef;
             14'h371e 	:	val_out <= 16'hf9f1;
             14'h371f 	:	val_out <= 16'hf9f2;
             14'h3720 	:	val_out <= 16'hf9f4;
             14'h3721 	:	val_out <= 16'hf9f5;
             14'h3722 	:	val_out <= 16'hf9f6;
             14'h3723 	:	val_out <= 16'hf9f8;
             14'h3724 	:	val_out <= 16'hf9f9;
             14'h3725 	:	val_out <= 16'hf9fa;
             14'h3726 	:	val_out <= 16'hf9fc;
             14'h3727 	:	val_out <= 16'hf9fd;
             14'h3728 	:	val_out <= 16'hf9fe;
             14'h3729 	:	val_out <= 16'hfa00;
             14'h372a 	:	val_out <= 16'hfa01;
             14'h372b 	:	val_out <= 16'hfa02;
             14'h372c 	:	val_out <= 16'hfa04;
             14'h372d 	:	val_out <= 16'hfa05;
             14'h372e 	:	val_out <= 16'hfa06;
             14'h372f 	:	val_out <= 16'hfa08;
             14'h3730 	:	val_out <= 16'hfa09;
             14'h3731 	:	val_out <= 16'hfa0b;
             14'h3732 	:	val_out <= 16'hfa0c;
             14'h3733 	:	val_out <= 16'hfa0d;
             14'h3734 	:	val_out <= 16'hfa0f;
             14'h3735 	:	val_out <= 16'hfa10;
             14'h3736 	:	val_out <= 16'hfa11;
             14'h3737 	:	val_out <= 16'hfa13;
             14'h3738 	:	val_out <= 16'hfa14;
             14'h3739 	:	val_out <= 16'hfa15;
             14'h373a 	:	val_out <= 16'hfa17;
             14'h373b 	:	val_out <= 16'hfa18;
             14'h373c 	:	val_out <= 16'hfa19;
             14'h373d 	:	val_out <= 16'hfa1b;
             14'h373e 	:	val_out <= 16'hfa1c;
             14'h373f 	:	val_out <= 16'hfa1d;
             14'h3740 	:	val_out <= 16'hfa1f;
             14'h3741 	:	val_out <= 16'hfa20;
             14'h3742 	:	val_out <= 16'hfa21;
             14'h3743 	:	val_out <= 16'hfa23;
             14'h3744 	:	val_out <= 16'hfa24;
             14'h3745 	:	val_out <= 16'hfa25;
             14'h3746 	:	val_out <= 16'hfa27;
             14'h3747 	:	val_out <= 16'hfa28;
             14'h3748 	:	val_out <= 16'hfa29;
             14'h3749 	:	val_out <= 16'hfa2b;
             14'h374a 	:	val_out <= 16'hfa2c;
             14'h374b 	:	val_out <= 16'hfa2d;
             14'h374c 	:	val_out <= 16'hfa2f;
             14'h374d 	:	val_out <= 16'hfa30;
             14'h374e 	:	val_out <= 16'hfa31;
             14'h374f 	:	val_out <= 16'hfa33;
             14'h3750 	:	val_out <= 16'hfa34;
             14'h3751 	:	val_out <= 16'hfa35;
             14'h3752 	:	val_out <= 16'hfa37;
             14'h3753 	:	val_out <= 16'hfa38;
             14'h3754 	:	val_out <= 16'hfa39;
             14'h3755 	:	val_out <= 16'hfa3b;
             14'h3756 	:	val_out <= 16'hfa3c;
             14'h3757 	:	val_out <= 16'hfa3d;
             14'h3758 	:	val_out <= 16'hfa3f;
             14'h3759 	:	val_out <= 16'hfa40;
             14'h375a 	:	val_out <= 16'hfa41;
             14'h375b 	:	val_out <= 16'hfa43;
             14'h375c 	:	val_out <= 16'hfa44;
             14'h375d 	:	val_out <= 16'hfa45;
             14'h375e 	:	val_out <= 16'hfa47;
             14'h375f 	:	val_out <= 16'hfa48;
             14'h3760 	:	val_out <= 16'hfa49;
             14'h3761 	:	val_out <= 16'hfa4b;
             14'h3762 	:	val_out <= 16'hfa4c;
             14'h3763 	:	val_out <= 16'hfa4d;
             14'h3764 	:	val_out <= 16'hfa4e;
             14'h3765 	:	val_out <= 16'hfa50;
             14'h3766 	:	val_out <= 16'hfa51;
             14'h3767 	:	val_out <= 16'hfa52;
             14'h3768 	:	val_out <= 16'hfa54;
             14'h3769 	:	val_out <= 16'hfa55;
             14'h376a 	:	val_out <= 16'hfa56;
             14'h376b 	:	val_out <= 16'hfa58;
             14'h376c 	:	val_out <= 16'hfa59;
             14'h376d 	:	val_out <= 16'hfa5a;
             14'h376e 	:	val_out <= 16'hfa5c;
             14'h376f 	:	val_out <= 16'hfa5d;
             14'h3770 	:	val_out <= 16'hfa5e;
             14'h3771 	:	val_out <= 16'hfa60;
             14'h3772 	:	val_out <= 16'hfa61;
             14'h3773 	:	val_out <= 16'hfa62;
             14'h3774 	:	val_out <= 16'hfa64;
             14'h3775 	:	val_out <= 16'hfa65;
             14'h3776 	:	val_out <= 16'hfa66;
             14'h3777 	:	val_out <= 16'hfa67;
             14'h3778 	:	val_out <= 16'hfa69;
             14'h3779 	:	val_out <= 16'hfa6a;
             14'h377a 	:	val_out <= 16'hfa6b;
             14'h377b 	:	val_out <= 16'hfa6d;
             14'h377c 	:	val_out <= 16'hfa6e;
             14'h377d 	:	val_out <= 16'hfa6f;
             14'h377e 	:	val_out <= 16'hfa71;
             14'h377f 	:	val_out <= 16'hfa72;
             14'h3780 	:	val_out <= 16'hfa73;
             14'h3781 	:	val_out <= 16'hfa74;
             14'h3782 	:	val_out <= 16'hfa76;
             14'h3783 	:	val_out <= 16'hfa77;
             14'h3784 	:	val_out <= 16'hfa78;
             14'h3785 	:	val_out <= 16'hfa7a;
             14'h3786 	:	val_out <= 16'hfa7b;
             14'h3787 	:	val_out <= 16'hfa7c;
             14'h3788 	:	val_out <= 16'hfa7e;
             14'h3789 	:	val_out <= 16'hfa7f;
             14'h378a 	:	val_out <= 16'hfa80;
             14'h378b 	:	val_out <= 16'hfa81;
             14'h378c 	:	val_out <= 16'hfa83;
             14'h378d 	:	val_out <= 16'hfa84;
             14'h378e 	:	val_out <= 16'hfa85;
             14'h378f 	:	val_out <= 16'hfa87;
             14'h3790 	:	val_out <= 16'hfa88;
             14'h3791 	:	val_out <= 16'hfa89;
             14'h3792 	:	val_out <= 16'hfa8a;
             14'h3793 	:	val_out <= 16'hfa8c;
             14'h3794 	:	val_out <= 16'hfa8d;
             14'h3795 	:	val_out <= 16'hfa8e;
             14'h3796 	:	val_out <= 16'hfa90;
             14'h3797 	:	val_out <= 16'hfa91;
             14'h3798 	:	val_out <= 16'hfa92;
             14'h3799 	:	val_out <= 16'hfa93;
             14'h379a 	:	val_out <= 16'hfa95;
             14'h379b 	:	val_out <= 16'hfa96;
             14'h379c 	:	val_out <= 16'hfa97;
             14'h379d 	:	val_out <= 16'hfa99;
             14'h379e 	:	val_out <= 16'hfa9a;
             14'h379f 	:	val_out <= 16'hfa9b;
             14'h37a0 	:	val_out <= 16'hfa9c;
             14'h37a1 	:	val_out <= 16'hfa9e;
             14'h37a2 	:	val_out <= 16'hfa9f;
             14'h37a3 	:	val_out <= 16'hfaa0;
             14'h37a4 	:	val_out <= 16'hfaa2;
             14'h37a5 	:	val_out <= 16'hfaa3;
             14'h37a6 	:	val_out <= 16'hfaa4;
             14'h37a7 	:	val_out <= 16'hfaa5;
             14'h37a8 	:	val_out <= 16'hfaa7;
             14'h37a9 	:	val_out <= 16'hfaa8;
             14'h37aa 	:	val_out <= 16'hfaa9;
             14'h37ab 	:	val_out <= 16'hfaab;
             14'h37ac 	:	val_out <= 16'hfaac;
             14'h37ad 	:	val_out <= 16'hfaad;
             14'h37ae 	:	val_out <= 16'hfaae;
             14'h37af 	:	val_out <= 16'hfab0;
             14'h37b0 	:	val_out <= 16'hfab1;
             14'h37b1 	:	val_out <= 16'hfab2;
             14'h37b2 	:	val_out <= 16'hfab3;
             14'h37b3 	:	val_out <= 16'hfab5;
             14'h37b4 	:	val_out <= 16'hfab6;
             14'h37b5 	:	val_out <= 16'hfab7;
             14'h37b6 	:	val_out <= 16'hfab9;
             14'h37b7 	:	val_out <= 16'hfaba;
             14'h37b8 	:	val_out <= 16'hfabb;
             14'h37b9 	:	val_out <= 16'hfabc;
             14'h37ba 	:	val_out <= 16'hfabe;
             14'h37bb 	:	val_out <= 16'hfabf;
             14'h37bc 	:	val_out <= 16'hfac0;
             14'h37bd 	:	val_out <= 16'hfac1;
             14'h37be 	:	val_out <= 16'hfac3;
             14'h37bf 	:	val_out <= 16'hfac4;
             14'h37c0 	:	val_out <= 16'hfac5;
             14'h37c1 	:	val_out <= 16'hfac6;
             14'h37c2 	:	val_out <= 16'hfac8;
             14'h37c3 	:	val_out <= 16'hfac9;
             14'h37c4 	:	val_out <= 16'hfaca;
             14'h37c5 	:	val_out <= 16'hfacc;
             14'h37c6 	:	val_out <= 16'hfacd;
             14'h37c7 	:	val_out <= 16'hface;
             14'h37c8 	:	val_out <= 16'hfacf;
             14'h37c9 	:	val_out <= 16'hfad1;
             14'h37ca 	:	val_out <= 16'hfad2;
             14'h37cb 	:	val_out <= 16'hfad3;
             14'h37cc 	:	val_out <= 16'hfad4;
             14'h37cd 	:	val_out <= 16'hfad6;
             14'h37ce 	:	val_out <= 16'hfad7;
             14'h37cf 	:	val_out <= 16'hfad8;
             14'h37d0 	:	val_out <= 16'hfad9;
             14'h37d1 	:	val_out <= 16'hfadb;
             14'h37d2 	:	val_out <= 16'hfadc;
             14'h37d3 	:	val_out <= 16'hfadd;
             14'h37d4 	:	val_out <= 16'hfade;
             14'h37d5 	:	val_out <= 16'hfae0;
             14'h37d6 	:	val_out <= 16'hfae1;
             14'h37d7 	:	val_out <= 16'hfae2;
             14'h37d8 	:	val_out <= 16'hfae3;
             14'h37d9 	:	val_out <= 16'hfae5;
             14'h37da 	:	val_out <= 16'hfae6;
             14'h37db 	:	val_out <= 16'hfae7;
             14'h37dc 	:	val_out <= 16'hfae8;
             14'h37dd 	:	val_out <= 16'hfaea;
             14'h37de 	:	val_out <= 16'hfaeb;
             14'h37df 	:	val_out <= 16'hfaec;
             14'h37e0 	:	val_out <= 16'hfaed;
             14'h37e1 	:	val_out <= 16'hfaef;
             14'h37e2 	:	val_out <= 16'hfaf0;
             14'h37e3 	:	val_out <= 16'hfaf1;
             14'h37e4 	:	val_out <= 16'hfaf2;
             14'h37e5 	:	val_out <= 16'hfaf4;
             14'h37e6 	:	val_out <= 16'hfaf5;
             14'h37e7 	:	val_out <= 16'hfaf6;
             14'h37e8 	:	val_out <= 16'hfaf7;
             14'h37e9 	:	val_out <= 16'hfaf9;
             14'h37ea 	:	val_out <= 16'hfafa;
             14'h37eb 	:	val_out <= 16'hfafb;
             14'h37ec 	:	val_out <= 16'hfafc;
             14'h37ed 	:	val_out <= 16'hfafd;
             14'h37ee 	:	val_out <= 16'hfaff;
             14'h37ef 	:	val_out <= 16'hfb00;
             14'h37f0 	:	val_out <= 16'hfb01;
             14'h37f1 	:	val_out <= 16'hfb02;
             14'h37f2 	:	val_out <= 16'hfb04;
             14'h37f3 	:	val_out <= 16'hfb05;
             14'h37f4 	:	val_out <= 16'hfb06;
             14'h37f5 	:	val_out <= 16'hfb07;
             14'h37f6 	:	val_out <= 16'hfb09;
             14'h37f7 	:	val_out <= 16'hfb0a;
             14'h37f8 	:	val_out <= 16'hfb0b;
             14'h37f9 	:	val_out <= 16'hfb0c;
             14'h37fa 	:	val_out <= 16'hfb0d;
             14'h37fb 	:	val_out <= 16'hfb0f;
             14'h37fc 	:	val_out <= 16'hfb10;
             14'h37fd 	:	val_out <= 16'hfb11;
             14'h37fe 	:	val_out <= 16'hfb12;
             14'h37ff 	:	val_out <= 16'hfb14;
             14'h3800 	:	val_out <= 16'hfb15;
             14'h3801 	:	val_out <= 16'hfb16;
             14'h3802 	:	val_out <= 16'hfb17;
             14'h3803 	:	val_out <= 16'hfb19;
             14'h3804 	:	val_out <= 16'hfb1a;
             14'h3805 	:	val_out <= 16'hfb1b;
             14'h3806 	:	val_out <= 16'hfb1c;
             14'h3807 	:	val_out <= 16'hfb1d;
             14'h3808 	:	val_out <= 16'hfb1f;
             14'h3809 	:	val_out <= 16'hfb20;
             14'h380a 	:	val_out <= 16'hfb21;
             14'h380b 	:	val_out <= 16'hfb22;
             14'h380c 	:	val_out <= 16'hfb24;
             14'h380d 	:	val_out <= 16'hfb25;
             14'h380e 	:	val_out <= 16'hfb26;
             14'h380f 	:	val_out <= 16'hfb27;
             14'h3810 	:	val_out <= 16'hfb28;
             14'h3811 	:	val_out <= 16'hfb2a;
             14'h3812 	:	val_out <= 16'hfb2b;
             14'h3813 	:	val_out <= 16'hfb2c;
             14'h3814 	:	val_out <= 16'hfb2d;
             14'h3815 	:	val_out <= 16'hfb2e;
             14'h3816 	:	val_out <= 16'hfb30;
             14'h3817 	:	val_out <= 16'hfb31;
             14'h3818 	:	val_out <= 16'hfb32;
             14'h3819 	:	val_out <= 16'hfb33;
             14'h381a 	:	val_out <= 16'hfb35;
             14'h381b 	:	val_out <= 16'hfb36;
             14'h381c 	:	val_out <= 16'hfb37;
             14'h381d 	:	val_out <= 16'hfb38;
             14'h381e 	:	val_out <= 16'hfb39;
             14'h381f 	:	val_out <= 16'hfb3b;
             14'h3820 	:	val_out <= 16'hfb3c;
             14'h3821 	:	val_out <= 16'hfb3d;
             14'h3822 	:	val_out <= 16'hfb3e;
             14'h3823 	:	val_out <= 16'hfb3f;
             14'h3824 	:	val_out <= 16'hfb41;
             14'h3825 	:	val_out <= 16'hfb42;
             14'h3826 	:	val_out <= 16'hfb43;
             14'h3827 	:	val_out <= 16'hfb44;
             14'h3828 	:	val_out <= 16'hfb45;
             14'h3829 	:	val_out <= 16'hfb47;
             14'h382a 	:	val_out <= 16'hfb48;
             14'h382b 	:	val_out <= 16'hfb49;
             14'h382c 	:	val_out <= 16'hfb4a;
             14'h382d 	:	val_out <= 16'hfb4b;
             14'h382e 	:	val_out <= 16'hfb4d;
             14'h382f 	:	val_out <= 16'hfb4e;
             14'h3830 	:	val_out <= 16'hfb4f;
             14'h3831 	:	val_out <= 16'hfb50;
             14'h3832 	:	val_out <= 16'hfb51;
             14'h3833 	:	val_out <= 16'hfb53;
             14'h3834 	:	val_out <= 16'hfb54;
             14'h3835 	:	val_out <= 16'hfb55;
             14'h3836 	:	val_out <= 16'hfb56;
             14'h3837 	:	val_out <= 16'hfb57;
             14'h3838 	:	val_out <= 16'hfb59;
             14'h3839 	:	val_out <= 16'hfb5a;
             14'h383a 	:	val_out <= 16'hfb5b;
             14'h383b 	:	val_out <= 16'hfb5c;
             14'h383c 	:	val_out <= 16'hfb5d;
             14'h383d 	:	val_out <= 16'hfb5f;
             14'h383e 	:	val_out <= 16'hfb60;
             14'h383f 	:	val_out <= 16'hfb61;
             14'h3840 	:	val_out <= 16'hfb62;
             14'h3841 	:	val_out <= 16'hfb63;
             14'h3842 	:	val_out <= 16'hfb64;
             14'h3843 	:	val_out <= 16'hfb66;
             14'h3844 	:	val_out <= 16'hfb67;
             14'h3845 	:	val_out <= 16'hfb68;
             14'h3846 	:	val_out <= 16'hfb69;
             14'h3847 	:	val_out <= 16'hfb6a;
             14'h3848 	:	val_out <= 16'hfb6c;
             14'h3849 	:	val_out <= 16'hfb6d;
             14'h384a 	:	val_out <= 16'hfb6e;
             14'h384b 	:	val_out <= 16'hfb6f;
             14'h384c 	:	val_out <= 16'hfb70;
             14'h384d 	:	val_out <= 16'hfb71;
             14'h384e 	:	val_out <= 16'hfb73;
             14'h384f 	:	val_out <= 16'hfb74;
             14'h3850 	:	val_out <= 16'hfb75;
             14'h3851 	:	val_out <= 16'hfb76;
             14'h3852 	:	val_out <= 16'hfb77;
             14'h3853 	:	val_out <= 16'hfb79;
             14'h3854 	:	val_out <= 16'hfb7a;
             14'h3855 	:	val_out <= 16'hfb7b;
             14'h3856 	:	val_out <= 16'hfb7c;
             14'h3857 	:	val_out <= 16'hfb7d;
             14'h3858 	:	val_out <= 16'hfb7e;
             14'h3859 	:	val_out <= 16'hfb80;
             14'h385a 	:	val_out <= 16'hfb81;
             14'h385b 	:	val_out <= 16'hfb82;
             14'h385c 	:	val_out <= 16'hfb83;
             14'h385d 	:	val_out <= 16'hfb84;
             14'h385e 	:	val_out <= 16'hfb85;
             14'h385f 	:	val_out <= 16'hfb87;
             14'h3860 	:	val_out <= 16'hfb88;
             14'h3861 	:	val_out <= 16'hfb89;
             14'h3862 	:	val_out <= 16'hfb8a;
             14'h3863 	:	val_out <= 16'hfb8b;
             14'h3864 	:	val_out <= 16'hfb8c;
             14'h3865 	:	val_out <= 16'hfb8e;
             14'h3866 	:	val_out <= 16'hfb8f;
             14'h3867 	:	val_out <= 16'hfb90;
             14'h3868 	:	val_out <= 16'hfb91;
             14'h3869 	:	val_out <= 16'hfb92;
             14'h386a 	:	val_out <= 16'hfb93;
             14'h386b 	:	val_out <= 16'hfb95;
             14'h386c 	:	val_out <= 16'hfb96;
             14'h386d 	:	val_out <= 16'hfb97;
             14'h386e 	:	val_out <= 16'hfb98;
             14'h386f 	:	val_out <= 16'hfb99;
             14'h3870 	:	val_out <= 16'hfb9a;
             14'h3871 	:	val_out <= 16'hfb9c;
             14'h3872 	:	val_out <= 16'hfb9d;
             14'h3873 	:	val_out <= 16'hfb9e;
             14'h3874 	:	val_out <= 16'hfb9f;
             14'h3875 	:	val_out <= 16'hfba0;
             14'h3876 	:	val_out <= 16'hfba1;
             14'h3877 	:	val_out <= 16'hfba3;
             14'h3878 	:	val_out <= 16'hfba4;
             14'h3879 	:	val_out <= 16'hfba5;
             14'h387a 	:	val_out <= 16'hfba6;
             14'h387b 	:	val_out <= 16'hfba7;
             14'h387c 	:	val_out <= 16'hfba8;
             14'h387d 	:	val_out <= 16'hfba9;
             14'h387e 	:	val_out <= 16'hfbab;
             14'h387f 	:	val_out <= 16'hfbac;
             14'h3880 	:	val_out <= 16'hfbad;
             14'h3881 	:	val_out <= 16'hfbae;
             14'h3882 	:	val_out <= 16'hfbaf;
             14'h3883 	:	val_out <= 16'hfbb0;
             14'h3884 	:	val_out <= 16'hfbb1;
             14'h3885 	:	val_out <= 16'hfbb3;
             14'h3886 	:	val_out <= 16'hfbb4;
             14'h3887 	:	val_out <= 16'hfbb5;
             14'h3888 	:	val_out <= 16'hfbb6;
             14'h3889 	:	val_out <= 16'hfbb7;
             14'h388a 	:	val_out <= 16'hfbb8;
             14'h388b 	:	val_out <= 16'hfbb9;
             14'h388c 	:	val_out <= 16'hfbbb;
             14'h388d 	:	val_out <= 16'hfbbc;
             14'h388e 	:	val_out <= 16'hfbbd;
             14'h388f 	:	val_out <= 16'hfbbe;
             14'h3890 	:	val_out <= 16'hfbbf;
             14'h3891 	:	val_out <= 16'hfbc0;
             14'h3892 	:	val_out <= 16'hfbc1;
             14'h3893 	:	val_out <= 16'hfbc3;
             14'h3894 	:	val_out <= 16'hfbc4;
             14'h3895 	:	val_out <= 16'hfbc5;
             14'h3896 	:	val_out <= 16'hfbc6;
             14'h3897 	:	val_out <= 16'hfbc7;
             14'h3898 	:	val_out <= 16'hfbc8;
             14'h3899 	:	val_out <= 16'hfbc9;
             14'h389a 	:	val_out <= 16'hfbcb;
             14'h389b 	:	val_out <= 16'hfbcc;
             14'h389c 	:	val_out <= 16'hfbcd;
             14'h389d 	:	val_out <= 16'hfbce;
             14'h389e 	:	val_out <= 16'hfbcf;
             14'h389f 	:	val_out <= 16'hfbd0;
             14'h38a0 	:	val_out <= 16'hfbd1;
             14'h38a1 	:	val_out <= 16'hfbd2;
             14'h38a2 	:	val_out <= 16'hfbd4;
             14'h38a3 	:	val_out <= 16'hfbd5;
             14'h38a4 	:	val_out <= 16'hfbd6;
             14'h38a5 	:	val_out <= 16'hfbd7;
             14'h38a6 	:	val_out <= 16'hfbd8;
             14'h38a7 	:	val_out <= 16'hfbd9;
             14'h38a8 	:	val_out <= 16'hfbda;
             14'h38a9 	:	val_out <= 16'hfbdc;
             14'h38aa 	:	val_out <= 16'hfbdd;
             14'h38ab 	:	val_out <= 16'hfbde;
             14'h38ac 	:	val_out <= 16'hfbdf;
             14'h38ad 	:	val_out <= 16'hfbe0;
             14'h38ae 	:	val_out <= 16'hfbe1;
             14'h38af 	:	val_out <= 16'hfbe2;
             14'h38b0 	:	val_out <= 16'hfbe3;
             14'h38b1 	:	val_out <= 16'hfbe5;
             14'h38b2 	:	val_out <= 16'hfbe6;
             14'h38b3 	:	val_out <= 16'hfbe7;
             14'h38b4 	:	val_out <= 16'hfbe8;
             14'h38b5 	:	val_out <= 16'hfbe9;
             14'h38b6 	:	val_out <= 16'hfbea;
             14'h38b7 	:	val_out <= 16'hfbeb;
             14'h38b8 	:	val_out <= 16'hfbec;
             14'h38b9 	:	val_out <= 16'hfbed;
             14'h38ba 	:	val_out <= 16'hfbef;
             14'h38bb 	:	val_out <= 16'hfbf0;
             14'h38bc 	:	val_out <= 16'hfbf1;
             14'h38bd 	:	val_out <= 16'hfbf2;
             14'h38be 	:	val_out <= 16'hfbf3;
             14'h38bf 	:	val_out <= 16'hfbf4;
             14'h38c0 	:	val_out <= 16'hfbf5;
             14'h38c1 	:	val_out <= 16'hfbf6;
             14'h38c2 	:	val_out <= 16'hfbf7;
             14'h38c3 	:	val_out <= 16'hfbf9;
             14'h38c4 	:	val_out <= 16'hfbfa;
             14'h38c5 	:	val_out <= 16'hfbfb;
             14'h38c6 	:	val_out <= 16'hfbfc;
             14'h38c7 	:	val_out <= 16'hfbfd;
             14'h38c8 	:	val_out <= 16'hfbfe;
             14'h38c9 	:	val_out <= 16'hfbff;
             14'h38ca 	:	val_out <= 16'hfc00;
             14'h38cb 	:	val_out <= 16'hfc01;
             14'h38cc 	:	val_out <= 16'hfc03;
             14'h38cd 	:	val_out <= 16'hfc04;
             14'h38ce 	:	val_out <= 16'hfc05;
             14'h38cf 	:	val_out <= 16'hfc06;
             14'h38d0 	:	val_out <= 16'hfc07;
             14'h38d1 	:	val_out <= 16'hfc08;
             14'h38d2 	:	val_out <= 16'hfc09;
             14'h38d3 	:	val_out <= 16'hfc0a;
             14'h38d4 	:	val_out <= 16'hfc0b;
             14'h38d5 	:	val_out <= 16'hfc0c;
             14'h38d6 	:	val_out <= 16'hfc0e;
             14'h38d7 	:	val_out <= 16'hfc0f;
             14'h38d8 	:	val_out <= 16'hfc10;
             14'h38d9 	:	val_out <= 16'hfc11;
             14'h38da 	:	val_out <= 16'hfc12;
             14'h38db 	:	val_out <= 16'hfc13;
             14'h38dc 	:	val_out <= 16'hfc14;
             14'h38dd 	:	val_out <= 16'hfc15;
             14'h38de 	:	val_out <= 16'hfc16;
             14'h38df 	:	val_out <= 16'hfc17;
             14'h38e0 	:	val_out <= 16'hfc19;
             14'h38e1 	:	val_out <= 16'hfc1a;
             14'h38e2 	:	val_out <= 16'hfc1b;
             14'h38e3 	:	val_out <= 16'hfc1c;
             14'h38e4 	:	val_out <= 16'hfc1d;
             14'h38e5 	:	val_out <= 16'hfc1e;
             14'h38e6 	:	val_out <= 16'hfc1f;
             14'h38e7 	:	val_out <= 16'hfc20;
             14'h38e8 	:	val_out <= 16'hfc21;
             14'h38e9 	:	val_out <= 16'hfc22;
             14'h38ea 	:	val_out <= 16'hfc23;
             14'h38eb 	:	val_out <= 16'hfc25;
             14'h38ec 	:	val_out <= 16'hfc26;
             14'h38ed 	:	val_out <= 16'hfc27;
             14'h38ee 	:	val_out <= 16'hfc28;
             14'h38ef 	:	val_out <= 16'hfc29;
             14'h38f0 	:	val_out <= 16'hfc2a;
             14'h38f1 	:	val_out <= 16'hfc2b;
             14'h38f2 	:	val_out <= 16'hfc2c;
             14'h38f3 	:	val_out <= 16'hfc2d;
             14'h38f4 	:	val_out <= 16'hfc2e;
             14'h38f5 	:	val_out <= 16'hfc2f;
             14'h38f6 	:	val_out <= 16'hfc30;
             14'h38f7 	:	val_out <= 16'hfc32;
             14'h38f8 	:	val_out <= 16'hfc33;
             14'h38f9 	:	val_out <= 16'hfc34;
             14'h38fa 	:	val_out <= 16'hfc35;
             14'h38fb 	:	val_out <= 16'hfc36;
             14'h38fc 	:	val_out <= 16'hfc37;
             14'h38fd 	:	val_out <= 16'hfc38;
             14'h38fe 	:	val_out <= 16'hfc39;
             14'h38ff 	:	val_out <= 16'hfc3a;
             14'h3900 	:	val_out <= 16'hfc3b;
             14'h3901 	:	val_out <= 16'hfc3c;
             14'h3902 	:	val_out <= 16'hfc3d;
             14'h3903 	:	val_out <= 16'hfc3e;
             14'h3904 	:	val_out <= 16'hfc3f;
             14'h3905 	:	val_out <= 16'hfc41;
             14'h3906 	:	val_out <= 16'hfc42;
             14'h3907 	:	val_out <= 16'hfc43;
             14'h3908 	:	val_out <= 16'hfc44;
             14'h3909 	:	val_out <= 16'hfc45;
             14'h390a 	:	val_out <= 16'hfc46;
             14'h390b 	:	val_out <= 16'hfc47;
             14'h390c 	:	val_out <= 16'hfc48;
             14'h390d 	:	val_out <= 16'hfc49;
             14'h390e 	:	val_out <= 16'hfc4a;
             14'h390f 	:	val_out <= 16'hfc4b;
             14'h3910 	:	val_out <= 16'hfc4c;
             14'h3911 	:	val_out <= 16'hfc4d;
             14'h3912 	:	val_out <= 16'hfc4e;
             14'h3913 	:	val_out <= 16'hfc4f;
             14'h3914 	:	val_out <= 16'hfc51;
             14'h3915 	:	val_out <= 16'hfc52;
             14'h3916 	:	val_out <= 16'hfc53;
             14'h3917 	:	val_out <= 16'hfc54;
             14'h3918 	:	val_out <= 16'hfc55;
             14'h3919 	:	val_out <= 16'hfc56;
             14'h391a 	:	val_out <= 16'hfc57;
             14'h391b 	:	val_out <= 16'hfc58;
             14'h391c 	:	val_out <= 16'hfc59;
             14'h391d 	:	val_out <= 16'hfc5a;
             14'h391e 	:	val_out <= 16'hfc5b;
             14'h391f 	:	val_out <= 16'hfc5c;
             14'h3920 	:	val_out <= 16'hfc5d;
             14'h3921 	:	val_out <= 16'hfc5e;
             14'h3922 	:	val_out <= 16'hfc5f;
             14'h3923 	:	val_out <= 16'hfc60;
             14'h3924 	:	val_out <= 16'hfc61;
             14'h3925 	:	val_out <= 16'hfc63;
             14'h3926 	:	val_out <= 16'hfc64;
             14'h3927 	:	val_out <= 16'hfc65;
             14'h3928 	:	val_out <= 16'hfc66;
             14'h3929 	:	val_out <= 16'hfc67;
             14'h392a 	:	val_out <= 16'hfc68;
             14'h392b 	:	val_out <= 16'hfc69;
             14'h392c 	:	val_out <= 16'hfc6a;
             14'h392d 	:	val_out <= 16'hfc6b;
             14'h392e 	:	val_out <= 16'hfc6c;
             14'h392f 	:	val_out <= 16'hfc6d;
             14'h3930 	:	val_out <= 16'hfc6e;
             14'h3931 	:	val_out <= 16'hfc6f;
             14'h3932 	:	val_out <= 16'hfc70;
             14'h3933 	:	val_out <= 16'hfc71;
             14'h3934 	:	val_out <= 16'hfc72;
             14'h3935 	:	val_out <= 16'hfc73;
             14'h3936 	:	val_out <= 16'hfc74;
             14'h3937 	:	val_out <= 16'hfc75;
             14'h3938 	:	val_out <= 16'hfc76;
             14'h3939 	:	val_out <= 16'hfc77;
             14'h393a 	:	val_out <= 16'hfc78;
             14'h393b 	:	val_out <= 16'hfc7a;
             14'h393c 	:	val_out <= 16'hfc7b;
             14'h393d 	:	val_out <= 16'hfc7c;
             14'h393e 	:	val_out <= 16'hfc7d;
             14'h393f 	:	val_out <= 16'hfc7e;
             14'h3940 	:	val_out <= 16'hfc7f;
             14'h3941 	:	val_out <= 16'hfc80;
             14'h3942 	:	val_out <= 16'hfc81;
             14'h3943 	:	val_out <= 16'hfc82;
             14'h3944 	:	val_out <= 16'hfc83;
             14'h3945 	:	val_out <= 16'hfc84;
             14'h3946 	:	val_out <= 16'hfc85;
             14'h3947 	:	val_out <= 16'hfc86;
             14'h3948 	:	val_out <= 16'hfc87;
             14'h3949 	:	val_out <= 16'hfc88;
             14'h394a 	:	val_out <= 16'hfc89;
             14'h394b 	:	val_out <= 16'hfc8a;
             14'h394c 	:	val_out <= 16'hfc8b;
             14'h394d 	:	val_out <= 16'hfc8c;
             14'h394e 	:	val_out <= 16'hfc8d;
             14'h394f 	:	val_out <= 16'hfc8e;
             14'h3950 	:	val_out <= 16'hfc8f;
             14'h3951 	:	val_out <= 16'hfc90;
             14'h3952 	:	val_out <= 16'hfc91;
             14'h3953 	:	val_out <= 16'hfc92;
             14'h3954 	:	val_out <= 16'hfc93;
             14'h3955 	:	val_out <= 16'hfc94;
             14'h3956 	:	val_out <= 16'hfc95;
             14'h3957 	:	val_out <= 16'hfc96;
             14'h3958 	:	val_out <= 16'hfc97;
             14'h3959 	:	val_out <= 16'hfc98;
             14'h395a 	:	val_out <= 16'hfc99;
             14'h395b 	:	val_out <= 16'hfc9a;
             14'h395c 	:	val_out <= 16'hfc9b;
             14'h395d 	:	val_out <= 16'hfc9c;
             14'h395e 	:	val_out <= 16'hfc9e;
             14'h395f 	:	val_out <= 16'hfc9f;
             14'h3960 	:	val_out <= 16'hfca0;
             14'h3961 	:	val_out <= 16'hfca1;
             14'h3962 	:	val_out <= 16'hfca2;
             14'h3963 	:	val_out <= 16'hfca3;
             14'h3964 	:	val_out <= 16'hfca4;
             14'h3965 	:	val_out <= 16'hfca5;
             14'h3966 	:	val_out <= 16'hfca6;
             14'h3967 	:	val_out <= 16'hfca7;
             14'h3968 	:	val_out <= 16'hfca8;
             14'h3969 	:	val_out <= 16'hfca9;
             14'h396a 	:	val_out <= 16'hfcaa;
             14'h396b 	:	val_out <= 16'hfcab;
             14'h396c 	:	val_out <= 16'hfcac;
             14'h396d 	:	val_out <= 16'hfcad;
             14'h396e 	:	val_out <= 16'hfcae;
             14'h396f 	:	val_out <= 16'hfcaf;
             14'h3970 	:	val_out <= 16'hfcb0;
             14'h3971 	:	val_out <= 16'hfcb1;
             14'h3972 	:	val_out <= 16'hfcb2;
             14'h3973 	:	val_out <= 16'hfcb3;
             14'h3974 	:	val_out <= 16'hfcb4;
             14'h3975 	:	val_out <= 16'hfcb5;
             14'h3976 	:	val_out <= 16'hfcb6;
             14'h3977 	:	val_out <= 16'hfcb7;
             14'h3978 	:	val_out <= 16'hfcb8;
             14'h3979 	:	val_out <= 16'hfcb9;
             14'h397a 	:	val_out <= 16'hfcba;
             14'h397b 	:	val_out <= 16'hfcbb;
             14'h397c 	:	val_out <= 16'hfcbc;
             14'h397d 	:	val_out <= 16'hfcbd;
             14'h397e 	:	val_out <= 16'hfcbe;
             14'h397f 	:	val_out <= 16'hfcbf;
             14'h3980 	:	val_out <= 16'hfcc0;
             14'h3981 	:	val_out <= 16'hfcc1;
             14'h3982 	:	val_out <= 16'hfcc2;
             14'h3983 	:	val_out <= 16'hfcc3;
             14'h3984 	:	val_out <= 16'hfcc4;
             14'h3985 	:	val_out <= 16'hfcc5;
             14'h3986 	:	val_out <= 16'hfcc6;
             14'h3987 	:	val_out <= 16'hfcc7;
             14'h3988 	:	val_out <= 16'hfcc8;
             14'h3989 	:	val_out <= 16'hfcc9;
             14'h398a 	:	val_out <= 16'hfcca;
             14'h398b 	:	val_out <= 16'hfccb;
             14'h398c 	:	val_out <= 16'hfccc;
             14'h398d 	:	val_out <= 16'hfccd;
             14'h398e 	:	val_out <= 16'hfcce;
             14'h398f 	:	val_out <= 16'hfccf;
             14'h3990 	:	val_out <= 16'hfcd0;
             14'h3991 	:	val_out <= 16'hfcd1;
             14'h3992 	:	val_out <= 16'hfcd2;
             14'h3993 	:	val_out <= 16'hfcd3;
             14'h3994 	:	val_out <= 16'hfcd4;
             14'h3995 	:	val_out <= 16'hfcd5;
             14'h3996 	:	val_out <= 16'hfcd6;
             14'h3997 	:	val_out <= 16'hfcd7;
             14'h3998 	:	val_out <= 16'hfcd8;
             14'h3999 	:	val_out <= 16'hfcd9;
             14'h399a 	:	val_out <= 16'hfcda;
             14'h399b 	:	val_out <= 16'hfcdb;
             14'h399c 	:	val_out <= 16'hfcdb;
             14'h399d 	:	val_out <= 16'hfcdc;
             14'h399e 	:	val_out <= 16'hfcdd;
             14'h399f 	:	val_out <= 16'hfcde;
             14'h39a0 	:	val_out <= 16'hfcdf;
             14'h39a1 	:	val_out <= 16'hfce0;
             14'h39a2 	:	val_out <= 16'hfce1;
             14'h39a3 	:	val_out <= 16'hfce2;
             14'h39a4 	:	val_out <= 16'hfce3;
             14'h39a5 	:	val_out <= 16'hfce4;
             14'h39a6 	:	val_out <= 16'hfce5;
             14'h39a7 	:	val_out <= 16'hfce6;
             14'h39a8 	:	val_out <= 16'hfce7;
             14'h39a9 	:	val_out <= 16'hfce8;
             14'h39aa 	:	val_out <= 16'hfce9;
             14'h39ab 	:	val_out <= 16'hfcea;
             14'h39ac 	:	val_out <= 16'hfceb;
             14'h39ad 	:	val_out <= 16'hfcec;
             14'h39ae 	:	val_out <= 16'hfced;
             14'h39af 	:	val_out <= 16'hfcee;
             14'h39b0 	:	val_out <= 16'hfcef;
             14'h39b1 	:	val_out <= 16'hfcf0;
             14'h39b2 	:	val_out <= 16'hfcf1;
             14'h39b3 	:	val_out <= 16'hfcf2;
             14'h39b4 	:	val_out <= 16'hfcf3;
             14'h39b5 	:	val_out <= 16'hfcf4;
             14'h39b6 	:	val_out <= 16'hfcf5;
             14'h39b7 	:	val_out <= 16'hfcf6;
             14'h39b8 	:	val_out <= 16'hfcf7;
             14'h39b9 	:	val_out <= 16'hfcf8;
             14'h39ba 	:	val_out <= 16'hfcf9;
             14'h39bb 	:	val_out <= 16'hfcfa;
             14'h39bc 	:	val_out <= 16'hfcfb;
             14'h39bd 	:	val_out <= 16'hfcfc;
             14'h39be 	:	val_out <= 16'hfcfd;
             14'h39bf 	:	val_out <= 16'hfcfd;
             14'h39c0 	:	val_out <= 16'hfcfe;
             14'h39c1 	:	val_out <= 16'hfcff;
             14'h39c2 	:	val_out <= 16'hfd00;
             14'h39c3 	:	val_out <= 16'hfd01;
             14'h39c4 	:	val_out <= 16'hfd02;
             14'h39c5 	:	val_out <= 16'hfd03;
             14'h39c6 	:	val_out <= 16'hfd04;
             14'h39c7 	:	val_out <= 16'hfd05;
             14'h39c8 	:	val_out <= 16'hfd06;
             14'h39c9 	:	val_out <= 16'hfd07;
             14'h39ca 	:	val_out <= 16'hfd08;
             14'h39cb 	:	val_out <= 16'hfd09;
             14'h39cc 	:	val_out <= 16'hfd0a;
             14'h39cd 	:	val_out <= 16'hfd0b;
             14'h39ce 	:	val_out <= 16'hfd0c;
             14'h39cf 	:	val_out <= 16'hfd0d;
             14'h39d0 	:	val_out <= 16'hfd0e;
             14'h39d1 	:	val_out <= 16'hfd0f;
             14'h39d2 	:	val_out <= 16'hfd10;
             14'h39d3 	:	val_out <= 16'hfd11;
             14'h39d4 	:	val_out <= 16'hfd12;
             14'h39d5 	:	val_out <= 16'hfd12;
             14'h39d6 	:	val_out <= 16'hfd13;
             14'h39d7 	:	val_out <= 16'hfd14;
             14'h39d8 	:	val_out <= 16'hfd15;
             14'h39d9 	:	val_out <= 16'hfd16;
             14'h39da 	:	val_out <= 16'hfd17;
             14'h39db 	:	val_out <= 16'hfd18;
             14'h39dc 	:	val_out <= 16'hfd19;
             14'h39dd 	:	val_out <= 16'hfd1a;
             14'h39de 	:	val_out <= 16'hfd1b;
             14'h39df 	:	val_out <= 16'hfd1c;
             14'h39e0 	:	val_out <= 16'hfd1d;
             14'h39e1 	:	val_out <= 16'hfd1e;
             14'h39e2 	:	val_out <= 16'hfd1f;
             14'h39e3 	:	val_out <= 16'hfd20;
             14'h39e4 	:	val_out <= 16'hfd21;
             14'h39e5 	:	val_out <= 16'hfd22;
             14'h39e6 	:	val_out <= 16'hfd22;
             14'h39e7 	:	val_out <= 16'hfd23;
             14'h39e8 	:	val_out <= 16'hfd24;
             14'h39e9 	:	val_out <= 16'hfd25;
             14'h39ea 	:	val_out <= 16'hfd26;
             14'h39eb 	:	val_out <= 16'hfd27;
             14'h39ec 	:	val_out <= 16'hfd28;
             14'h39ed 	:	val_out <= 16'hfd29;
             14'h39ee 	:	val_out <= 16'hfd2a;
             14'h39ef 	:	val_out <= 16'hfd2b;
             14'h39f0 	:	val_out <= 16'hfd2c;
             14'h39f1 	:	val_out <= 16'hfd2d;
             14'h39f2 	:	val_out <= 16'hfd2e;
             14'h39f3 	:	val_out <= 16'hfd2f;
             14'h39f4 	:	val_out <= 16'hfd30;
             14'h39f5 	:	val_out <= 16'hfd30;
             14'h39f6 	:	val_out <= 16'hfd31;
             14'h39f7 	:	val_out <= 16'hfd32;
             14'h39f8 	:	val_out <= 16'hfd33;
             14'h39f9 	:	val_out <= 16'hfd34;
             14'h39fa 	:	val_out <= 16'hfd35;
             14'h39fb 	:	val_out <= 16'hfd36;
             14'h39fc 	:	val_out <= 16'hfd37;
             14'h39fd 	:	val_out <= 16'hfd38;
             14'h39fe 	:	val_out <= 16'hfd39;
             14'h39ff 	:	val_out <= 16'hfd3a;
             14'h3a00 	:	val_out <= 16'hfd3b;
             14'h3a01 	:	val_out <= 16'hfd3c;
             14'h3a02 	:	val_out <= 16'hfd3c;
             14'h3a03 	:	val_out <= 16'hfd3d;
             14'h3a04 	:	val_out <= 16'hfd3e;
             14'h3a05 	:	val_out <= 16'hfd3f;
             14'h3a06 	:	val_out <= 16'hfd40;
             14'h3a07 	:	val_out <= 16'hfd41;
             14'h3a08 	:	val_out <= 16'hfd42;
             14'h3a09 	:	val_out <= 16'hfd43;
             14'h3a0a 	:	val_out <= 16'hfd44;
             14'h3a0b 	:	val_out <= 16'hfd45;
             14'h3a0c 	:	val_out <= 16'hfd46;
             14'h3a0d 	:	val_out <= 16'hfd47;
             14'h3a0e 	:	val_out <= 16'hfd47;
             14'h3a0f 	:	val_out <= 16'hfd48;
             14'h3a10 	:	val_out <= 16'hfd49;
             14'h3a11 	:	val_out <= 16'hfd4a;
             14'h3a12 	:	val_out <= 16'hfd4b;
             14'h3a13 	:	val_out <= 16'hfd4c;
             14'h3a14 	:	val_out <= 16'hfd4d;
             14'h3a15 	:	val_out <= 16'hfd4e;
             14'h3a16 	:	val_out <= 16'hfd4f;
             14'h3a17 	:	val_out <= 16'hfd50;
             14'h3a18 	:	val_out <= 16'hfd51;
             14'h3a19 	:	val_out <= 16'hfd51;
             14'h3a1a 	:	val_out <= 16'hfd52;
             14'h3a1b 	:	val_out <= 16'hfd53;
             14'h3a1c 	:	val_out <= 16'hfd54;
             14'h3a1d 	:	val_out <= 16'hfd55;
             14'h3a1e 	:	val_out <= 16'hfd56;
             14'h3a1f 	:	val_out <= 16'hfd57;
             14'h3a20 	:	val_out <= 16'hfd58;
             14'h3a21 	:	val_out <= 16'hfd59;
             14'h3a22 	:	val_out <= 16'hfd5a;
             14'h3a23 	:	val_out <= 16'hfd5b;
             14'h3a24 	:	val_out <= 16'hfd5b;
             14'h3a25 	:	val_out <= 16'hfd5c;
             14'h3a26 	:	val_out <= 16'hfd5d;
             14'h3a27 	:	val_out <= 16'hfd5e;
             14'h3a28 	:	val_out <= 16'hfd5f;
             14'h3a29 	:	val_out <= 16'hfd60;
             14'h3a2a 	:	val_out <= 16'hfd61;
             14'h3a2b 	:	val_out <= 16'hfd62;
             14'h3a2c 	:	val_out <= 16'hfd63;
             14'h3a2d 	:	val_out <= 16'hfd64;
             14'h3a2e 	:	val_out <= 16'hfd64;
             14'h3a2f 	:	val_out <= 16'hfd65;
             14'h3a30 	:	val_out <= 16'hfd66;
             14'h3a31 	:	val_out <= 16'hfd67;
             14'h3a32 	:	val_out <= 16'hfd68;
             14'h3a33 	:	val_out <= 16'hfd69;
             14'h3a34 	:	val_out <= 16'hfd6a;
             14'h3a35 	:	val_out <= 16'hfd6b;
             14'h3a36 	:	val_out <= 16'hfd6c;
             14'h3a37 	:	val_out <= 16'hfd6c;
             14'h3a38 	:	val_out <= 16'hfd6d;
             14'h3a39 	:	val_out <= 16'hfd6e;
             14'h3a3a 	:	val_out <= 16'hfd6f;
             14'h3a3b 	:	val_out <= 16'hfd70;
             14'h3a3c 	:	val_out <= 16'hfd71;
             14'h3a3d 	:	val_out <= 16'hfd72;
             14'h3a3e 	:	val_out <= 16'hfd73;
             14'h3a3f 	:	val_out <= 16'hfd74;
             14'h3a40 	:	val_out <= 16'hfd74;
             14'h3a41 	:	val_out <= 16'hfd75;
             14'h3a42 	:	val_out <= 16'hfd76;
             14'h3a43 	:	val_out <= 16'hfd77;
             14'h3a44 	:	val_out <= 16'hfd78;
             14'h3a45 	:	val_out <= 16'hfd79;
             14'h3a46 	:	val_out <= 16'hfd7a;
             14'h3a47 	:	val_out <= 16'hfd7b;
             14'h3a48 	:	val_out <= 16'hfd7b;
             14'h3a49 	:	val_out <= 16'hfd7c;
             14'h3a4a 	:	val_out <= 16'hfd7d;
             14'h3a4b 	:	val_out <= 16'hfd7e;
             14'h3a4c 	:	val_out <= 16'hfd7f;
             14'h3a4d 	:	val_out <= 16'hfd80;
             14'h3a4e 	:	val_out <= 16'hfd81;
             14'h3a4f 	:	val_out <= 16'hfd82;
             14'h3a50 	:	val_out <= 16'hfd82;
             14'h3a51 	:	val_out <= 16'hfd83;
             14'h3a52 	:	val_out <= 16'hfd84;
             14'h3a53 	:	val_out <= 16'hfd85;
             14'h3a54 	:	val_out <= 16'hfd86;
             14'h3a55 	:	val_out <= 16'hfd87;
             14'h3a56 	:	val_out <= 16'hfd88;
             14'h3a57 	:	val_out <= 16'hfd89;
             14'h3a58 	:	val_out <= 16'hfd89;
             14'h3a59 	:	val_out <= 16'hfd8a;
             14'h3a5a 	:	val_out <= 16'hfd8b;
             14'h3a5b 	:	val_out <= 16'hfd8c;
             14'h3a5c 	:	val_out <= 16'hfd8d;
             14'h3a5d 	:	val_out <= 16'hfd8e;
             14'h3a5e 	:	val_out <= 16'hfd8f;
             14'h3a5f 	:	val_out <= 16'hfd8f;
             14'h3a60 	:	val_out <= 16'hfd90;
             14'h3a61 	:	val_out <= 16'hfd91;
             14'h3a62 	:	val_out <= 16'hfd92;
             14'h3a63 	:	val_out <= 16'hfd93;
             14'h3a64 	:	val_out <= 16'hfd94;
             14'h3a65 	:	val_out <= 16'hfd95;
             14'h3a66 	:	val_out <= 16'hfd96;
             14'h3a67 	:	val_out <= 16'hfd96;
             14'h3a68 	:	val_out <= 16'hfd97;
             14'h3a69 	:	val_out <= 16'hfd98;
             14'h3a6a 	:	val_out <= 16'hfd99;
             14'h3a6b 	:	val_out <= 16'hfd9a;
             14'h3a6c 	:	val_out <= 16'hfd9b;
             14'h3a6d 	:	val_out <= 16'hfd9c;
             14'h3a6e 	:	val_out <= 16'hfd9c;
             14'h3a6f 	:	val_out <= 16'hfd9d;
             14'h3a70 	:	val_out <= 16'hfd9e;
             14'h3a71 	:	val_out <= 16'hfd9f;
             14'h3a72 	:	val_out <= 16'hfda0;
             14'h3a73 	:	val_out <= 16'hfda1;
             14'h3a74 	:	val_out <= 16'hfda2;
             14'h3a75 	:	val_out <= 16'hfda2;
             14'h3a76 	:	val_out <= 16'hfda3;
             14'h3a77 	:	val_out <= 16'hfda4;
             14'h3a78 	:	val_out <= 16'hfda5;
             14'h3a79 	:	val_out <= 16'hfda6;
             14'h3a7a 	:	val_out <= 16'hfda7;
             14'h3a7b 	:	val_out <= 16'hfda7;
             14'h3a7c 	:	val_out <= 16'hfda8;
             14'h3a7d 	:	val_out <= 16'hfda9;
             14'h3a7e 	:	val_out <= 16'hfdaa;
             14'h3a7f 	:	val_out <= 16'hfdab;
             14'h3a80 	:	val_out <= 16'hfdac;
             14'h3a81 	:	val_out <= 16'hfdad;
             14'h3a82 	:	val_out <= 16'hfdad;
             14'h3a83 	:	val_out <= 16'hfdae;
             14'h3a84 	:	val_out <= 16'hfdaf;
             14'h3a85 	:	val_out <= 16'hfdb0;
             14'h3a86 	:	val_out <= 16'hfdb1;
             14'h3a87 	:	val_out <= 16'hfdb2;
             14'h3a88 	:	val_out <= 16'hfdb2;
             14'h3a89 	:	val_out <= 16'hfdb3;
             14'h3a8a 	:	val_out <= 16'hfdb4;
             14'h3a8b 	:	val_out <= 16'hfdb5;
             14'h3a8c 	:	val_out <= 16'hfdb6;
             14'h3a8d 	:	val_out <= 16'hfdb7;
             14'h3a8e 	:	val_out <= 16'hfdb7;
             14'h3a8f 	:	val_out <= 16'hfdb8;
             14'h3a90 	:	val_out <= 16'hfdb9;
             14'h3a91 	:	val_out <= 16'hfdba;
             14'h3a92 	:	val_out <= 16'hfdbb;
             14'h3a93 	:	val_out <= 16'hfdbc;
             14'h3a94 	:	val_out <= 16'hfdbd;
             14'h3a95 	:	val_out <= 16'hfdbd;
             14'h3a96 	:	val_out <= 16'hfdbe;
             14'h3a97 	:	val_out <= 16'hfdbf;
             14'h3a98 	:	val_out <= 16'hfdc0;
             14'h3a99 	:	val_out <= 16'hfdc1;
             14'h3a9a 	:	val_out <= 16'hfdc1;
             14'h3a9b 	:	val_out <= 16'hfdc2;
             14'h3a9c 	:	val_out <= 16'hfdc3;
             14'h3a9d 	:	val_out <= 16'hfdc4;
             14'h3a9e 	:	val_out <= 16'hfdc5;
             14'h3a9f 	:	val_out <= 16'hfdc6;
             14'h3aa0 	:	val_out <= 16'hfdc6;
             14'h3aa1 	:	val_out <= 16'hfdc7;
             14'h3aa2 	:	val_out <= 16'hfdc8;
             14'h3aa3 	:	val_out <= 16'hfdc9;
             14'h3aa4 	:	val_out <= 16'hfdca;
             14'h3aa5 	:	val_out <= 16'hfdcb;
             14'h3aa6 	:	val_out <= 16'hfdcb;
             14'h3aa7 	:	val_out <= 16'hfdcc;
             14'h3aa8 	:	val_out <= 16'hfdcd;
             14'h3aa9 	:	val_out <= 16'hfdce;
             14'h3aaa 	:	val_out <= 16'hfdcf;
             14'h3aab 	:	val_out <= 16'hfdd0;
             14'h3aac 	:	val_out <= 16'hfdd0;
             14'h3aad 	:	val_out <= 16'hfdd1;
             14'h3aae 	:	val_out <= 16'hfdd2;
             14'h3aaf 	:	val_out <= 16'hfdd3;
             14'h3ab0 	:	val_out <= 16'hfdd4;
             14'h3ab1 	:	val_out <= 16'hfdd4;
             14'h3ab2 	:	val_out <= 16'hfdd5;
             14'h3ab3 	:	val_out <= 16'hfdd6;
             14'h3ab4 	:	val_out <= 16'hfdd7;
             14'h3ab5 	:	val_out <= 16'hfdd8;
             14'h3ab6 	:	val_out <= 16'hfdd8;
             14'h3ab7 	:	val_out <= 16'hfdd9;
             14'h3ab8 	:	val_out <= 16'hfdda;
             14'h3ab9 	:	val_out <= 16'hfddb;
             14'h3aba 	:	val_out <= 16'hfddc;
             14'h3abb 	:	val_out <= 16'hfddd;
             14'h3abc 	:	val_out <= 16'hfddd;
             14'h3abd 	:	val_out <= 16'hfdde;
             14'h3abe 	:	val_out <= 16'hfddf;
             14'h3abf 	:	val_out <= 16'hfde0;
             14'h3ac0 	:	val_out <= 16'hfde1;
             14'h3ac1 	:	val_out <= 16'hfde1;
             14'h3ac2 	:	val_out <= 16'hfde2;
             14'h3ac3 	:	val_out <= 16'hfde3;
             14'h3ac4 	:	val_out <= 16'hfde4;
             14'h3ac5 	:	val_out <= 16'hfde5;
             14'h3ac6 	:	val_out <= 16'hfde5;
             14'h3ac7 	:	val_out <= 16'hfde6;
             14'h3ac8 	:	val_out <= 16'hfde7;
             14'h3ac9 	:	val_out <= 16'hfde8;
             14'h3aca 	:	val_out <= 16'hfde9;
             14'h3acb 	:	val_out <= 16'hfde9;
             14'h3acc 	:	val_out <= 16'hfdea;
             14'h3acd 	:	val_out <= 16'hfdeb;
             14'h3ace 	:	val_out <= 16'hfdec;
             14'h3acf 	:	val_out <= 16'hfded;
             14'h3ad0 	:	val_out <= 16'hfded;
             14'h3ad1 	:	val_out <= 16'hfdee;
             14'h3ad2 	:	val_out <= 16'hfdef;
             14'h3ad3 	:	val_out <= 16'hfdf0;
             14'h3ad4 	:	val_out <= 16'hfdf1;
             14'h3ad5 	:	val_out <= 16'hfdf1;
             14'h3ad6 	:	val_out <= 16'hfdf2;
             14'h3ad7 	:	val_out <= 16'hfdf3;
             14'h3ad8 	:	val_out <= 16'hfdf4;
             14'h3ad9 	:	val_out <= 16'hfdf5;
             14'h3ada 	:	val_out <= 16'hfdf5;
             14'h3adb 	:	val_out <= 16'hfdf6;
             14'h3adc 	:	val_out <= 16'hfdf7;
             14'h3add 	:	val_out <= 16'hfdf8;
             14'h3ade 	:	val_out <= 16'hfdf9;
             14'h3adf 	:	val_out <= 16'hfdf9;
             14'h3ae0 	:	val_out <= 16'hfdfa;
             14'h3ae1 	:	val_out <= 16'hfdfb;
             14'h3ae2 	:	val_out <= 16'hfdfc;
             14'h3ae3 	:	val_out <= 16'hfdfc;
             14'h3ae4 	:	val_out <= 16'hfdfd;
             14'h3ae5 	:	val_out <= 16'hfdfe;
             14'h3ae6 	:	val_out <= 16'hfdff;
             14'h3ae7 	:	val_out <= 16'hfe00;
             14'h3ae8 	:	val_out <= 16'hfe00;
             14'h3ae9 	:	val_out <= 16'hfe01;
             14'h3aea 	:	val_out <= 16'hfe02;
             14'h3aeb 	:	val_out <= 16'hfe03;
             14'h3aec 	:	val_out <= 16'hfe04;
             14'h3aed 	:	val_out <= 16'hfe04;
             14'h3aee 	:	val_out <= 16'hfe05;
             14'h3aef 	:	val_out <= 16'hfe06;
             14'h3af0 	:	val_out <= 16'hfe07;
             14'h3af1 	:	val_out <= 16'hfe07;
             14'h3af2 	:	val_out <= 16'hfe08;
             14'h3af3 	:	val_out <= 16'hfe09;
             14'h3af4 	:	val_out <= 16'hfe0a;
             14'h3af5 	:	val_out <= 16'hfe0b;
             14'h3af6 	:	val_out <= 16'hfe0b;
             14'h3af7 	:	val_out <= 16'hfe0c;
             14'h3af8 	:	val_out <= 16'hfe0d;
             14'h3af9 	:	val_out <= 16'hfe0e;
             14'h3afa 	:	val_out <= 16'hfe0e;
             14'h3afb 	:	val_out <= 16'hfe0f;
             14'h3afc 	:	val_out <= 16'hfe10;
             14'h3afd 	:	val_out <= 16'hfe11;
             14'h3afe 	:	val_out <= 16'hfe11;
             14'h3aff 	:	val_out <= 16'hfe12;
             14'h3b00 	:	val_out <= 16'hfe13;
             14'h3b01 	:	val_out <= 16'hfe14;
             14'h3b02 	:	val_out <= 16'hfe15;
             14'h3b03 	:	val_out <= 16'hfe15;
             14'h3b04 	:	val_out <= 16'hfe16;
             14'h3b05 	:	val_out <= 16'hfe17;
             14'h3b06 	:	val_out <= 16'hfe18;
             14'h3b07 	:	val_out <= 16'hfe18;
             14'h3b08 	:	val_out <= 16'hfe19;
             14'h3b09 	:	val_out <= 16'hfe1a;
             14'h3b0a 	:	val_out <= 16'hfe1b;
             14'h3b0b 	:	val_out <= 16'hfe1b;
             14'h3b0c 	:	val_out <= 16'hfe1c;
             14'h3b0d 	:	val_out <= 16'hfe1d;
             14'h3b0e 	:	val_out <= 16'hfe1e;
             14'h3b0f 	:	val_out <= 16'hfe1e;
             14'h3b10 	:	val_out <= 16'hfe1f;
             14'h3b11 	:	val_out <= 16'hfe20;
             14'h3b12 	:	val_out <= 16'hfe21;
             14'h3b13 	:	val_out <= 16'hfe22;
             14'h3b14 	:	val_out <= 16'hfe22;
             14'h3b15 	:	val_out <= 16'hfe23;
             14'h3b16 	:	val_out <= 16'hfe24;
             14'h3b17 	:	val_out <= 16'hfe25;
             14'h3b18 	:	val_out <= 16'hfe25;
             14'h3b19 	:	val_out <= 16'hfe26;
             14'h3b1a 	:	val_out <= 16'hfe27;
             14'h3b1b 	:	val_out <= 16'hfe28;
             14'h3b1c 	:	val_out <= 16'hfe28;
             14'h3b1d 	:	val_out <= 16'hfe29;
             14'h3b1e 	:	val_out <= 16'hfe2a;
             14'h3b1f 	:	val_out <= 16'hfe2b;
             14'h3b20 	:	val_out <= 16'hfe2b;
             14'h3b21 	:	val_out <= 16'hfe2c;
             14'h3b22 	:	val_out <= 16'hfe2d;
             14'h3b23 	:	val_out <= 16'hfe2e;
             14'h3b24 	:	val_out <= 16'hfe2e;
             14'h3b25 	:	val_out <= 16'hfe2f;
             14'h3b26 	:	val_out <= 16'hfe30;
             14'h3b27 	:	val_out <= 16'hfe31;
             14'h3b28 	:	val_out <= 16'hfe31;
             14'h3b29 	:	val_out <= 16'hfe32;
             14'h3b2a 	:	val_out <= 16'hfe33;
             14'h3b2b 	:	val_out <= 16'hfe34;
             14'h3b2c 	:	val_out <= 16'hfe34;
             14'h3b2d 	:	val_out <= 16'hfe35;
             14'h3b2e 	:	val_out <= 16'hfe36;
             14'h3b2f 	:	val_out <= 16'hfe36;
             14'h3b30 	:	val_out <= 16'hfe37;
             14'h3b31 	:	val_out <= 16'hfe38;
             14'h3b32 	:	val_out <= 16'hfe39;
             14'h3b33 	:	val_out <= 16'hfe39;
             14'h3b34 	:	val_out <= 16'hfe3a;
             14'h3b35 	:	val_out <= 16'hfe3b;
             14'h3b36 	:	val_out <= 16'hfe3c;
             14'h3b37 	:	val_out <= 16'hfe3c;
             14'h3b38 	:	val_out <= 16'hfe3d;
             14'h3b39 	:	val_out <= 16'hfe3e;
             14'h3b3a 	:	val_out <= 16'hfe3f;
             14'h3b3b 	:	val_out <= 16'hfe3f;
             14'h3b3c 	:	val_out <= 16'hfe40;
             14'h3b3d 	:	val_out <= 16'hfe41;
             14'h3b3e 	:	val_out <= 16'hfe42;
             14'h3b3f 	:	val_out <= 16'hfe42;
             14'h3b40 	:	val_out <= 16'hfe43;
             14'h3b41 	:	val_out <= 16'hfe44;
             14'h3b42 	:	val_out <= 16'hfe44;
             14'h3b43 	:	val_out <= 16'hfe45;
             14'h3b44 	:	val_out <= 16'hfe46;
             14'h3b45 	:	val_out <= 16'hfe47;
             14'h3b46 	:	val_out <= 16'hfe47;
             14'h3b47 	:	val_out <= 16'hfe48;
             14'h3b48 	:	val_out <= 16'hfe49;
             14'h3b49 	:	val_out <= 16'hfe4a;
             14'h3b4a 	:	val_out <= 16'hfe4a;
             14'h3b4b 	:	val_out <= 16'hfe4b;
             14'h3b4c 	:	val_out <= 16'hfe4c;
             14'h3b4d 	:	val_out <= 16'hfe4c;
             14'h3b4e 	:	val_out <= 16'hfe4d;
             14'h3b4f 	:	val_out <= 16'hfe4e;
             14'h3b50 	:	val_out <= 16'hfe4f;
             14'h3b51 	:	val_out <= 16'hfe4f;
             14'h3b52 	:	val_out <= 16'hfe50;
             14'h3b53 	:	val_out <= 16'hfe51;
             14'h3b54 	:	val_out <= 16'hfe51;
             14'h3b55 	:	val_out <= 16'hfe52;
             14'h3b56 	:	val_out <= 16'hfe53;
             14'h3b57 	:	val_out <= 16'hfe54;
             14'h3b58 	:	val_out <= 16'hfe54;
             14'h3b59 	:	val_out <= 16'hfe55;
             14'h3b5a 	:	val_out <= 16'hfe56;
             14'h3b5b 	:	val_out <= 16'hfe57;
             14'h3b5c 	:	val_out <= 16'hfe57;
             14'h3b5d 	:	val_out <= 16'hfe58;
             14'h3b5e 	:	val_out <= 16'hfe59;
             14'h3b5f 	:	val_out <= 16'hfe59;
             14'h3b60 	:	val_out <= 16'hfe5a;
             14'h3b61 	:	val_out <= 16'hfe5b;
             14'h3b62 	:	val_out <= 16'hfe5b;
             14'h3b63 	:	val_out <= 16'hfe5c;
             14'h3b64 	:	val_out <= 16'hfe5d;
             14'h3b65 	:	val_out <= 16'hfe5e;
             14'h3b66 	:	val_out <= 16'hfe5e;
             14'h3b67 	:	val_out <= 16'hfe5f;
             14'h3b68 	:	val_out <= 16'hfe60;
             14'h3b69 	:	val_out <= 16'hfe60;
             14'h3b6a 	:	val_out <= 16'hfe61;
             14'h3b6b 	:	val_out <= 16'hfe62;
             14'h3b6c 	:	val_out <= 16'hfe63;
             14'h3b6d 	:	val_out <= 16'hfe63;
             14'h3b6e 	:	val_out <= 16'hfe64;
             14'h3b6f 	:	val_out <= 16'hfe65;
             14'h3b70 	:	val_out <= 16'hfe65;
             14'h3b71 	:	val_out <= 16'hfe66;
             14'h3b72 	:	val_out <= 16'hfe67;
             14'h3b73 	:	val_out <= 16'hfe67;
             14'h3b74 	:	val_out <= 16'hfe68;
             14'h3b75 	:	val_out <= 16'hfe69;
             14'h3b76 	:	val_out <= 16'hfe6a;
             14'h3b77 	:	val_out <= 16'hfe6a;
             14'h3b78 	:	val_out <= 16'hfe6b;
             14'h3b79 	:	val_out <= 16'hfe6c;
             14'h3b7a 	:	val_out <= 16'hfe6c;
             14'h3b7b 	:	val_out <= 16'hfe6d;
             14'h3b7c 	:	val_out <= 16'hfe6e;
             14'h3b7d 	:	val_out <= 16'hfe6e;
             14'h3b7e 	:	val_out <= 16'hfe6f;
             14'h3b7f 	:	val_out <= 16'hfe70;
             14'h3b80 	:	val_out <= 16'hfe71;
             14'h3b81 	:	val_out <= 16'hfe71;
             14'h3b82 	:	val_out <= 16'hfe72;
             14'h3b83 	:	val_out <= 16'hfe73;
             14'h3b84 	:	val_out <= 16'hfe73;
             14'h3b85 	:	val_out <= 16'hfe74;
             14'h3b86 	:	val_out <= 16'hfe75;
             14'h3b87 	:	val_out <= 16'hfe75;
             14'h3b88 	:	val_out <= 16'hfe76;
             14'h3b89 	:	val_out <= 16'hfe77;
             14'h3b8a 	:	val_out <= 16'hfe77;
             14'h3b8b 	:	val_out <= 16'hfe78;
             14'h3b8c 	:	val_out <= 16'hfe79;
             14'h3b8d 	:	val_out <= 16'hfe79;
             14'h3b8e 	:	val_out <= 16'hfe7a;
             14'h3b8f 	:	val_out <= 16'hfe7b;
             14'h3b90 	:	val_out <= 16'hfe7c;
             14'h3b91 	:	val_out <= 16'hfe7c;
             14'h3b92 	:	val_out <= 16'hfe7d;
             14'h3b93 	:	val_out <= 16'hfe7e;
             14'h3b94 	:	val_out <= 16'hfe7e;
             14'h3b95 	:	val_out <= 16'hfe7f;
             14'h3b96 	:	val_out <= 16'hfe80;
             14'h3b97 	:	val_out <= 16'hfe80;
             14'h3b98 	:	val_out <= 16'hfe81;
             14'h3b99 	:	val_out <= 16'hfe82;
             14'h3b9a 	:	val_out <= 16'hfe82;
             14'h3b9b 	:	val_out <= 16'hfe83;
             14'h3b9c 	:	val_out <= 16'hfe84;
             14'h3b9d 	:	val_out <= 16'hfe84;
             14'h3b9e 	:	val_out <= 16'hfe85;
             14'h3b9f 	:	val_out <= 16'hfe86;
             14'h3ba0 	:	val_out <= 16'hfe86;
             14'h3ba1 	:	val_out <= 16'hfe87;
             14'h3ba2 	:	val_out <= 16'hfe88;
             14'h3ba3 	:	val_out <= 16'hfe88;
             14'h3ba4 	:	val_out <= 16'hfe89;
             14'h3ba5 	:	val_out <= 16'hfe8a;
             14'h3ba6 	:	val_out <= 16'hfe8a;
             14'h3ba7 	:	val_out <= 16'hfe8b;
             14'h3ba8 	:	val_out <= 16'hfe8c;
             14'h3ba9 	:	val_out <= 16'hfe8c;
             14'h3baa 	:	val_out <= 16'hfe8d;
             14'h3bab 	:	val_out <= 16'hfe8e;
             14'h3bac 	:	val_out <= 16'hfe8e;
             14'h3bad 	:	val_out <= 16'hfe8f;
             14'h3bae 	:	val_out <= 16'hfe90;
             14'h3baf 	:	val_out <= 16'hfe90;
             14'h3bb0 	:	val_out <= 16'hfe91;
             14'h3bb1 	:	val_out <= 16'hfe92;
             14'h3bb2 	:	val_out <= 16'hfe92;
             14'h3bb3 	:	val_out <= 16'hfe93;
             14'h3bb4 	:	val_out <= 16'hfe94;
             14'h3bb5 	:	val_out <= 16'hfe94;
             14'h3bb6 	:	val_out <= 16'hfe95;
             14'h3bb7 	:	val_out <= 16'hfe96;
             14'h3bb8 	:	val_out <= 16'hfe96;
             14'h3bb9 	:	val_out <= 16'hfe97;
             14'h3bba 	:	val_out <= 16'hfe98;
             14'h3bbb 	:	val_out <= 16'hfe98;
             14'h3bbc 	:	val_out <= 16'hfe99;
             14'h3bbd 	:	val_out <= 16'hfe9a;
             14'h3bbe 	:	val_out <= 16'hfe9a;
             14'h3bbf 	:	val_out <= 16'hfe9b;
             14'h3bc0 	:	val_out <= 16'hfe9c;
             14'h3bc1 	:	val_out <= 16'hfe9c;
             14'h3bc2 	:	val_out <= 16'hfe9d;
             14'h3bc3 	:	val_out <= 16'hfe9e;
             14'h3bc4 	:	val_out <= 16'hfe9e;
             14'h3bc5 	:	val_out <= 16'hfe9f;
             14'h3bc6 	:	val_out <= 16'hfea0;
             14'h3bc7 	:	val_out <= 16'hfea0;
             14'h3bc8 	:	val_out <= 16'hfea1;
             14'h3bc9 	:	val_out <= 16'hfea1;
             14'h3bca 	:	val_out <= 16'hfea2;
             14'h3bcb 	:	val_out <= 16'hfea3;
             14'h3bcc 	:	val_out <= 16'hfea3;
             14'h3bcd 	:	val_out <= 16'hfea4;
             14'h3bce 	:	val_out <= 16'hfea5;
             14'h3bcf 	:	val_out <= 16'hfea5;
             14'h3bd0 	:	val_out <= 16'hfea6;
             14'h3bd1 	:	val_out <= 16'hfea7;
             14'h3bd2 	:	val_out <= 16'hfea7;
             14'h3bd3 	:	val_out <= 16'hfea8;
             14'h3bd4 	:	val_out <= 16'hfea9;
             14'h3bd5 	:	val_out <= 16'hfea9;
             14'h3bd6 	:	val_out <= 16'hfeaa;
             14'h3bd7 	:	val_out <= 16'hfeaa;
             14'h3bd8 	:	val_out <= 16'hfeab;
             14'h3bd9 	:	val_out <= 16'hfeac;
             14'h3bda 	:	val_out <= 16'hfeac;
             14'h3bdb 	:	val_out <= 16'hfead;
             14'h3bdc 	:	val_out <= 16'hfeae;
             14'h3bdd 	:	val_out <= 16'hfeae;
             14'h3bde 	:	val_out <= 16'hfeaf;
             14'h3bdf 	:	val_out <= 16'hfeb0;
             14'h3be0 	:	val_out <= 16'hfeb0;
             14'h3be1 	:	val_out <= 16'hfeb1;
             14'h3be2 	:	val_out <= 16'hfeb1;
             14'h3be3 	:	val_out <= 16'hfeb2;
             14'h3be4 	:	val_out <= 16'hfeb3;
             14'h3be5 	:	val_out <= 16'hfeb3;
             14'h3be6 	:	val_out <= 16'hfeb4;
             14'h3be7 	:	val_out <= 16'hfeb5;
             14'h3be8 	:	val_out <= 16'hfeb5;
             14'h3be9 	:	val_out <= 16'hfeb6;
             14'h3bea 	:	val_out <= 16'hfeb7;
             14'h3beb 	:	val_out <= 16'hfeb7;
             14'h3bec 	:	val_out <= 16'hfeb8;
             14'h3bed 	:	val_out <= 16'hfeb8;
             14'h3bee 	:	val_out <= 16'hfeb9;
             14'h3bef 	:	val_out <= 16'hfeba;
             14'h3bf0 	:	val_out <= 16'hfeba;
             14'h3bf1 	:	val_out <= 16'hfebb;
             14'h3bf2 	:	val_out <= 16'hfebc;
             14'h3bf3 	:	val_out <= 16'hfebc;
             14'h3bf4 	:	val_out <= 16'hfebd;
             14'h3bf5 	:	val_out <= 16'hfebd;
             14'h3bf6 	:	val_out <= 16'hfebe;
             14'h3bf7 	:	val_out <= 16'hfebf;
             14'h3bf8 	:	val_out <= 16'hfebf;
             14'h3bf9 	:	val_out <= 16'hfec0;
             14'h3bfa 	:	val_out <= 16'hfec1;
             14'h3bfb 	:	val_out <= 16'hfec1;
             14'h3bfc 	:	val_out <= 16'hfec2;
             14'h3bfd 	:	val_out <= 16'hfec2;
             14'h3bfe 	:	val_out <= 16'hfec3;
             14'h3bff 	:	val_out <= 16'hfec4;
             14'h3c00 	:	val_out <= 16'hfec4;
             14'h3c01 	:	val_out <= 16'hfec5;
             14'h3c02 	:	val_out <= 16'hfec5;
             14'h3c03 	:	val_out <= 16'hfec6;
             14'h3c04 	:	val_out <= 16'hfec7;
             14'h3c05 	:	val_out <= 16'hfec7;
             14'h3c06 	:	val_out <= 16'hfec8;
             14'h3c07 	:	val_out <= 16'hfec9;
             14'h3c08 	:	val_out <= 16'hfec9;
             14'h3c09 	:	val_out <= 16'hfeca;
             14'h3c0a 	:	val_out <= 16'hfeca;
             14'h3c0b 	:	val_out <= 16'hfecb;
             14'h3c0c 	:	val_out <= 16'hfecc;
             14'h3c0d 	:	val_out <= 16'hfecc;
             14'h3c0e 	:	val_out <= 16'hfecd;
             14'h3c0f 	:	val_out <= 16'hfecd;
             14'h3c10 	:	val_out <= 16'hfece;
             14'h3c11 	:	val_out <= 16'hfecf;
             14'h3c12 	:	val_out <= 16'hfecf;
             14'h3c13 	:	val_out <= 16'hfed0;
             14'h3c14 	:	val_out <= 16'hfed0;
             14'h3c15 	:	val_out <= 16'hfed1;
             14'h3c16 	:	val_out <= 16'hfed2;
             14'h3c17 	:	val_out <= 16'hfed2;
             14'h3c18 	:	val_out <= 16'hfed3;
             14'h3c19 	:	val_out <= 16'hfed3;
             14'h3c1a 	:	val_out <= 16'hfed4;
             14'h3c1b 	:	val_out <= 16'hfed5;
             14'h3c1c 	:	val_out <= 16'hfed5;
             14'h3c1d 	:	val_out <= 16'hfed6;
             14'h3c1e 	:	val_out <= 16'hfed6;
             14'h3c1f 	:	val_out <= 16'hfed7;
             14'h3c20 	:	val_out <= 16'hfed8;
             14'h3c21 	:	val_out <= 16'hfed8;
             14'h3c22 	:	val_out <= 16'hfed9;
             14'h3c23 	:	val_out <= 16'hfed9;
             14'h3c24 	:	val_out <= 16'hfeda;
             14'h3c25 	:	val_out <= 16'hfedb;
             14'h3c26 	:	val_out <= 16'hfedb;
             14'h3c27 	:	val_out <= 16'hfedc;
             14'h3c28 	:	val_out <= 16'hfedc;
             14'h3c29 	:	val_out <= 16'hfedd;
             14'h3c2a 	:	val_out <= 16'hfede;
             14'h3c2b 	:	val_out <= 16'hfede;
             14'h3c2c 	:	val_out <= 16'hfedf;
             14'h3c2d 	:	val_out <= 16'hfedf;
             14'h3c2e 	:	val_out <= 16'hfee0;
             14'h3c2f 	:	val_out <= 16'hfee1;
             14'h3c30 	:	val_out <= 16'hfee1;
             14'h3c31 	:	val_out <= 16'hfee2;
             14'h3c32 	:	val_out <= 16'hfee2;
             14'h3c33 	:	val_out <= 16'hfee3;
             14'h3c34 	:	val_out <= 16'hfee3;
             14'h3c35 	:	val_out <= 16'hfee4;
             14'h3c36 	:	val_out <= 16'hfee5;
             14'h3c37 	:	val_out <= 16'hfee5;
             14'h3c38 	:	val_out <= 16'hfee6;
             14'h3c39 	:	val_out <= 16'hfee6;
             14'h3c3a 	:	val_out <= 16'hfee7;
             14'h3c3b 	:	val_out <= 16'hfee8;
             14'h3c3c 	:	val_out <= 16'hfee8;
             14'h3c3d 	:	val_out <= 16'hfee9;
             14'h3c3e 	:	val_out <= 16'hfee9;
             14'h3c3f 	:	val_out <= 16'hfeea;
             14'h3c40 	:	val_out <= 16'hfeea;
             14'h3c41 	:	val_out <= 16'hfeeb;
             14'h3c42 	:	val_out <= 16'hfeec;
             14'h3c43 	:	val_out <= 16'hfeec;
             14'h3c44 	:	val_out <= 16'hfeed;
             14'h3c45 	:	val_out <= 16'hfeed;
             14'h3c46 	:	val_out <= 16'hfeee;
             14'h3c47 	:	val_out <= 16'hfeee;
             14'h3c48 	:	val_out <= 16'hfeef;
             14'h3c49 	:	val_out <= 16'hfef0;
             14'h3c4a 	:	val_out <= 16'hfef0;
             14'h3c4b 	:	val_out <= 16'hfef1;
             14'h3c4c 	:	val_out <= 16'hfef1;
             14'h3c4d 	:	val_out <= 16'hfef2;
             14'h3c4e 	:	val_out <= 16'hfef2;
             14'h3c4f 	:	val_out <= 16'hfef3;
             14'h3c50 	:	val_out <= 16'hfef4;
             14'h3c51 	:	val_out <= 16'hfef4;
             14'h3c52 	:	val_out <= 16'hfef5;
             14'h3c53 	:	val_out <= 16'hfef5;
             14'h3c54 	:	val_out <= 16'hfef6;
             14'h3c55 	:	val_out <= 16'hfef6;
             14'h3c56 	:	val_out <= 16'hfef7;
             14'h3c57 	:	val_out <= 16'hfef8;
             14'h3c58 	:	val_out <= 16'hfef8;
             14'h3c59 	:	val_out <= 16'hfef9;
             14'h3c5a 	:	val_out <= 16'hfef9;
             14'h3c5b 	:	val_out <= 16'hfefa;
             14'h3c5c 	:	val_out <= 16'hfefa;
             14'h3c5d 	:	val_out <= 16'hfefb;
             14'h3c5e 	:	val_out <= 16'hfefb;
             14'h3c5f 	:	val_out <= 16'hfefc;
             14'h3c60 	:	val_out <= 16'hfefd;
             14'h3c61 	:	val_out <= 16'hfefd;
             14'h3c62 	:	val_out <= 16'hfefe;
             14'h3c63 	:	val_out <= 16'hfefe;
             14'h3c64 	:	val_out <= 16'hfeff;
             14'h3c65 	:	val_out <= 16'hfeff;
             14'h3c66 	:	val_out <= 16'hff00;
             14'h3c67 	:	val_out <= 16'hff00;
             14'h3c68 	:	val_out <= 16'hff01;
             14'h3c69 	:	val_out <= 16'hff02;
             14'h3c6a 	:	val_out <= 16'hff02;
             14'h3c6b 	:	val_out <= 16'hff03;
             14'h3c6c 	:	val_out <= 16'hff03;
             14'h3c6d 	:	val_out <= 16'hff04;
             14'h3c6e 	:	val_out <= 16'hff04;
             14'h3c6f 	:	val_out <= 16'hff05;
             14'h3c70 	:	val_out <= 16'hff05;
             14'h3c71 	:	val_out <= 16'hff06;
             14'h3c72 	:	val_out <= 16'hff07;
             14'h3c73 	:	val_out <= 16'hff07;
             14'h3c74 	:	val_out <= 16'hff08;
             14'h3c75 	:	val_out <= 16'hff08;
             14'h3c76 	:	val_out <= 16'hff09;
             14'h3c77 	:	val_out <= 16'hff09;
             14'h3c78 	:	val_out <= 16'hff0a;
             14'h3c79 	:	val_out <= 16'hff0a;
             14'h3c7a 	:	val_out <= 16'hff0b;
             14'h3c7b 	:	val_out <= 16'hff0b;
             14'h3c7c 	:	val_out <= 16'hff0c;
             14'h3c7d 	:	val_out <= 16'hff0c;
             14'h3c7e 	:	val_out <= 16'hff0d;
             14'h3c7f 	:	val_out <= 16'hff0e;
             14'h3c80 	:	val_out <= 16'hff0e;
             14'h3c81 	:	val_out <= 16'hff0f;
             14'h3c82 	:	val_out <= 16'hff0f;
             14'h3c83 	:	val_out <= 16'hff10;
             14'h3c84 	:	val_out <= 16'hff10;
             14'h3c85 	:	val_out <= 16'hff11;
             14'h3c86 	:	val_out <= 16'hff11;
             14'h3c87 	:	val_out <= 16'hff12;
             14'h3c88 	:	val_out <= 16'hff12;
             14'h3c89 	:	val_out <= 16'hff13;
             14'h3c8a 	:	val_out <= 16'hff13;
             14'h3c8b 	:	val_out <= 16'hff14;
             14'h3c8c 	:	val_out <= 16'hff15;
             14'h3c8d 	:	val_out <= 16'hff15;
             14'h3c8e 	:	val_out <= 16'hff16;
             14'h3c8f 	:	val_out <= 16'hff16;
             14'h3c90 	:	val_out <= 16'hff17;
             14'h3c91 	:	val_out <= 16'hff17;
             14'h3c92 	:	val_out <= 16'hff18;
             14'h3c93 	:	val_out <= 16'hff18;
             14'h3c94 	:	val_out <= 16'hff19;
             14'h3c95 	:	val_out <= 16'hff19;
             14'h3c96 	:	val_out <= 16'hff1a;
             14'h3c97 	:	val_out <= 16'hff1a;
             14'h3c98 	:	val_out <= 16'hff1b;
             14'h3c99 	:	val_out <= 16'hff1b;
             14'h3c9a 	:	val_out <= 16'hff1c;
             14'h3c9b 	:	val_out <= 16'hff1c;
             14'h3c9c 	:	val_out <= 16'hff1d;
             14'h3c9d 	:	val_out <= 16'hff1d;
             14'h3c9e 	:	val_out <= 16'hff1e;
             14'h3c9f 	:	val_out <= 16'hff1f;
             14'h3ca0 	:	val_out <= 16'hff1f;
             14'h3ca1 	:	val_out <= 16'hff20;
             14'h3ca2 	:	val_out <= 16'hff20;
             14'h3ca3 	:	val_out <= 16'hff21;
             14'h3ca4 	:	val_out <= 16'hff21;
             14'h3ca5 	:	val_out <= 16'hff22;
             14'h3ca6 	:	val_out <= 16'hff22;
             14'h3ca7 	:	val_out <= 16'hff23;
             14'h3ca8 	:	val_out <= 16'hff23;
             14'h3ca9 	:	val_out <= 16'hff24;
             14'h3caa 	:	val_out <= 16'hff24;
             14'h3cab 	:	val_out <= 16'hff25;
             14'h3cac 	:	val_out <= 16'hff25;
             14'h3cad 	:	val_out <= 16'hff26;
             14'h3cae 	:	val_out <= 16'hff26;
             14'h3caf 	:	val_out <= 16'hff27;
             14'h3cb0 	:	val_out <= 16'hff27;
             14'h3cb1 	:	val_out <= 16'hff28;
             14'h3cb2 	:	val_out <= 16'hff28;
             14'h3cb3 	:	val_out <= 16'hff29;
             14'h3cb4 	:	val_out <= 16'hff29;
             14'h3cb5 	:	val_out <= 16'hff2a;
             14'h3cb6 	:	val_out <= 16'hff2a;
             14'h3cb7 	:	val_out <= 16'hff2b;
             14'h3cb8 	:	val_out <= 16'hff2b;
             14'h3cb9 	:	val_out <= 16'hff2c;
             14'h3cba 	:	val_out <= 16'hff2c;
             14'h3cbb 	:	val_out <= 16'hff2d;
             14'h3cbc 	:	val_out <= 16'hff2d;
             14'h3cbd 	:	val_out <= 16'hff2e;
             14'h3cbe 	:	val_out <= 16'hff2e;
             14'h3cbf 	:	val_out <= 16'hff2f;
             14'h3cc0 	:	val_out <= 16'hff2f;
             14'h3cc1 	:	val_out <= 16'hff30;
             14'h3cc2 	:	val_out <= 16'hff30;
             14'h3cc3 	:	val_out <= 16'hff31;
             14'h3cc4 	:	val_out <= 16'hff31;
             14'h3cc5 	:	val_out <= 16'hff32;
             14'h3cc6 	:	val_out <= 16'hff32;
             14'h3cc7 	:	val_out <= 16'hff33;
             14'h3cc8 	:	val_out <= 16'hff33;
             14'h3cc9 	:	val_out <= 16'hff34;
             14'h3cca 	:	val_out <= 16'hff34;
             14'h3ccb 	:	val_out <= 16'hff35;
             14'h3ccc 	:	val_out <= 16'hff35;
             14'h3ccd 	:	val_out <= 16'hff36;
             14'h3cce 	:	val_out <= 16'hff36;
             14'h3ccf 	:	val_out <= 16'hff37;
             14'h3cd0 	:	val_out <= 16'hff37;
             14'h3cd1 	:	val_out <= 16'hff38;
             14'h3cd2 	:	val_out <= 16'hff38;
             14'h3cd3 	:	val_out <= 16'hff39;
             14'h3cd4 	:	val_out <= 16'hff39;
             14'h3cd5 	:	val_out <= 16'hff3a;
             14'h3cd6 	:	val_out <= 16'hff3a;
             14'h3cd7 	:	val_out <= 16'hff3b;
             14'h3cd8 	:	val_out <= 16'hff3b;
             14'h3cd9 	:	val_out <= 16'hff3c;
             14'h3cda 	:	val_out <= 16'hff3c;
             14'h3cdb 	:	val_out <= 16'hff3d;
             14'h3cdc 	:	val_out <= 16'hff3d;
             14'h3cdd 	:	val_out <= 16'hff3e;
             14'h3cde 	:	val_out <= 16'hff3e;
             14'h3cdf 	:	val_out <= 16'hff3f;
             14'h3ce0 	:	val_out <= 16'hff3f;
             14'h3ce1 	:	val_out <= 16'hff40;
             14'h3ce2 	:	val_out <= 16'hff40;
             14'h3ce3 	:	val_out <= 16'hff41;
             14'h3ce4 	:	val_out <= 16'hff41;
             14'h3ce5 	:	val_out <= 16'hff41;
             14'h3ce6 	:	val_out <= 16'hff42;
             14'h3ce7 	:	val_out <= 16'hff42;
             14'h3ce8 	:	val_out <= 16'hff43;
             14'h3ce9 	:	val_out <= 16'hff43;
             14'h3cea 	:	val_out <= 16'hff44;
             14'h3ceb 	:	val_out <= 16'hff44;
             14'h3cec 	:	val_out <= 16'hff45;
             14'h3ced 	:	val_out <= 16'hff45;
             14'h3cee 	:	val_out <= 16'hff46;
             14'h3cef 	:	val_out <= 16'hff46;
             14'h3cf0 	:	val_out <= 16'hff47;
             14'h3cf1 	:	val_out <= 16'hff47;
             14'h3cf2 	:	val_out <= 16'hff48;
             14'h3cf3 	:	val_out <= 16'hff48;
             14'h3cf4 	:	val_out <= 16'hff49;
             14'h3cf5 	:	val_out <= 16'hff49;
             14'h3cf6 	:	val_out <= 16'hff4a;
             14'h3cf7 	:	val_out <= 16'hff4a;
             14'h3cf8 	:	val_out <= 16'hff4a;
             14'h3cf9 	:	val_out <= 16'hff4b;
             14'h3cfa 	:	val_out <= 16'hff4b;
             14'h3cfb 	:	val_out <= 16'hff4c;
             14'h3cfc 	:	val_out <= 16'hff4c;
             14'h3cfd 	:	val_out <= 16'hff4d;
             14'h3cfe 	:	val_out <= 16'hff4d;
             14'h3cff 	:	val_out <= 16'hff4e;
             14'h3d00 	:	val_out <= 16'hff4e;
             14'h3d01 	:	val_out <= 16'hff4f;
             14'h3d02 	:	val_out <= 16'hff4f;
             14'h3d03 	:	val_out <= 16'hff50;
             14'h3d04 	:	val_out <= 16'hff50;
             14'h3d05 	:	val_out <= 16'hff50;
             14'h3d06 	:	val_out <= 16'hff51;
             14'h3d07 	:	val_out <= 16'hff51;
             14'h3d08 	:	val_out <= 16'hff52;
             14'h3d09 	:	val_out <= 16'hff52;
             14'h3d0a 	:	val_out <= 16'hff53;
             14'h3d0b 	:	val_out <= 16'hff53;
             14'h3d0c 	:	val_out <= 16'hff54;
             14'h3d0d 	:	val_out <= 16'hff54;
             14'h3d0e 	:	val_out <= 16'hff55;
             14'h3d0f 	:	val_out <= 16'hff55;
             14'h3d10 	:	val_out <= 16'hff55;
             14'h3d11 	:	val_out <= 16'hff56;
             14'h3d12 	:	val_out <= 16'hff56;
             14'h3d13 	:	val_out <= 16'hff57;
             14'h3d14 	:	val_out <= 16'hff57;
             14'h3d15 	:	val_out <= 16'hff58;
             14'h3d16 	:	val_out <= 16'hff58;
             14'h3d17 	:	val_out <= 16'hff59;
             14'h3d18 	:	val_out <= 16'hff59;
             14'h3d19 	:	val_out <= 16'hff5a;
             14'h3d1a 	:	val_out <= 16'hff5a;
             14'h3d1b 	:	val_out <= 16'hff5a;
             14'h3d1c 	:	val_out <= 16'hff5b;
             14'h3d1d 	:	val_out <= 16'hff5b;
             14'h3d1e 	:	val_out <= 16'hff5c;
             14'h3d1f 	:	val_out <= 16'hff5c;
             14'h3d20 	:	val_out <= 16'hff5d;
             14'h3d21 	:	val_out <= 16'hff5d;
             14'h3d22 	:	val_out <= 16'hff5e;
             14'h3d23 	:	val_out <= 16'hff5e;
             14'h3d24 	:	val_out <= 16'hff5e;
             14'h3d25 	:	val_out <= 16'hff5f;
             14'h3d26 	:	val_out <= 16'hff5f;
             14'h3d27 	:	val_out <= 16'hff60;
             14'h3d28 	:	val_out <= 16'hff60;
             14'h3d29 	:	val_out <= 16'hff61;
             14'h3d2a 	:	val_out <= 16'hff61;
             14'h3d2b 	:	val_out <= 16'hff61;
             14'h3d2c 	:	val_out <= 16'hff62;
             14'h3d2d 	:	val_out <= 16'hff62;
             14'h3d2e 	:	val_out <= 16'hff63;
             14'h3d2f 	:	val_out <= 16'hff63;
             14'h3d30 	:	val_out <= 16'hff64;
             14'h3d31 	:	val_out <= 16'hff64;
             14'h3d32 	:	val_out <= 16'hff65;
             14'h3d33 	:	val_out <= 16'hff65;
             14'h3d34 	:	val_out <= 16'hff65;
             14'h3d35 	:	val_out <= 16'hff66;
             14'h3d36 	:	val_out <= 16'hff66;
             14'h3d37 	:	val_out <= 16'hff67;
             14'h3d38 	:	val_out <= 16'hff67;
             14'h3d39 	:	val_out <= 16'hff68;
             14'h3d3a 	:	val_out <= 16'hff68;
             14'h3d3b 	:	val_out <= 16'hff68;
             14'h3d3c 	:	val_out <= 16'hff69;
             14'h3d3d 	:	val_out <= 16'hff69;
             14'h3d3e 	:	val_out <= 16'hff6a;
             14'h3d3f 	:	val_out <= 16'hff6a;
             14'h3d40 	:	val_out <= 16'hff6a;
             14'h3d41 	:	val_out <= 16'hff6b;
             14'h3d42 	:	val_out <= 16'hff6b;
             14'h3d43 	:	val_out <= 16'hff6c;
             14'h3d44 	:	val_out <= 16'hff6c;
             14'h3d45 	:	val_out <= 16'hff6d;
             14'h3d46 	:	val_out <= 16'hff6d;
             14'h3d47 	:	val_out <= 16'hff6d;
             14'h3d48 	:	val_out <= 16'hff6e;
             14'h3d49 	:	val_out <= 16'hff6e;
             14'h3d4a 	:	val_out <= 16'hff6f;
             14'h3d4b 	:	val_out <= 16'hff6f;
             14'h3d4c 	:	val_out <= 16'hff70;
             14'h3d4d 	:	val_out <= 16'hff70;
             14'h3d4e 	:	val_out <= 16'hff70;
             14'h3d4f 	:	val_out <= 16'hff71;
             14'h3d50 	:	val_out <= 16'hff71;
             14'h3d51 	:	val_out <= 16'hff72;
             14'h3d52 	:	val_out <= 16'hff72;
             14'h3d53 	:	val_out <= 16'hff72;
             14'h3d54 	:	val_out <= 16'hff73;
             14'h3d55 	:	val_out <= 16'hff73;
             14'h3d56 	:	val_out <= 16'hff74;
             14'h3d57 	:	val_out <= 16'hff74;
             14'h3d58 	:	val_out <= 16'hff74;
             14'h3d59 	:	val_out <= 16'hff75;
             14'h3d5a 	:	val_out <= 16'hff75;
             14'h3d5b 	:	val_out <= 16'hff76;
             14'h3d5c 	:	val_out <= 16'hff76;
             14'h3d5d 	:	val_out <= 16'hff77;
             14'h3d5e 	:	val_out <= 16'hff77;
             14'h3d5f 	:	val_out <= 16'hff77;
             14'h3d60 	:	val_out <= 16'hff78;
             14'h3d61 	:	val_out <= 16'hff78;
             14'h3d62 	:	val_out <= 16'hff79;
             14'h3d63 	:	val_out <= 16'hff79;
             14'h3d64 	:	val_out <= 16'hff79;
             14'h3d65 	:	val_out <= 16'hff7a;
             14'h3d66 	:	val_out <= 16'hff7a;
             14'h3d67 	:	val_out <= 16'hff7b;
             14'h3d68 	:	val_out <= 16'hff7b;
             14'h3d69 	:	val_out <= 16'hff7b;
             14'h3d6a 	:	val_out <= 16'hff7c;
             14'h3d6b 	:	val_out <= 16'hff7c;
             14'h3d6c 	:	val_out <= 16'hff7d;
             14'h3d6d 	:	val_out <= 16'hff7d;
             14'h3d6e 	:	val_out <= 16'hff7d;
             14'h3d6f 	:	val_out <= 16'hff7e;
             14'h3d70 	:	val_out <= 16'hff7e;
             14'h3d71 	:	val_out <= 16'hff7f;
             14'h3d72 	:	val_out <= 16'hff7f;
             14'h3d73 	:	val_out <= 16'hff7f;
             14'h3d74 	:	val_out <= 16'hff80;
             14'h3d75 	:	val_out <= 16'hff80;
             14'h3d76 	:	val_out <= 16'hff80;
             14'h3d77 	:	val_out <= 16'hff81;
             14'h3d78 	:	val_out <= 16'hff81;
             14'h3d79 	:	val_out <= 16'hff82;
             14'h3d7a 	:	val_out <= 16'hff82;
             14'h3d7b 	:	val_out <= 16'hff82;
             14'h3d7c 	:	val_out <= 16'hff83;
             14'h3d7d 	:	val_out <= 16'hff83;
             14'h3d7e 	:	val_out <= 16'hff84;
             14'h3d7f 	:	val_out <= 16'hff84;
             14'h3d80 	:	val_out <= 16'hff84;
             14'h3d81 	:	val_out <= 16'hff85;
             14'h3d82 	:	val_out <= 16'hff85;
             14'h3d83 	:	val_out <= 16'hff86;
             14'h3d84 	:	val_out <= 16'hff86;
             14'h3d85 	:	val_out <= 16'hff86;
             14'h3d86 	:	val_out <= 16'hff87;
             14'h3d87 	:	val_out <= 16'hff87;
             14'h3d88 	:	val_out <= 16'hff87;
             14'h3d89 	:	val_out <= 16'hff88;
             14'h3d8a 	:	val_out <= 16'hff88;
             14'h3d8b 	:	val_out <= 16'hff89;
             14'h3d8c 	:	val_out <= 16'hff89;
             14'h3d8d 	:	val_out <= 16'hff89;
             14'h3d8e 	:	val_out <= 16'hff8a;
             14'h3d8f 	:	val_out <= 16'hff8a;
             14'h3d90 	:	val_out <= 16'hff8a;
             14'h3d91 	:	val_out <= 16'hff8b;
             14'h3d92 	:	val_out <= 16'hff8b;
             14'h3d93 	:	val_out <= 16'hff8c;
             14'h3d94 	:	val_out <= 16'hff8c;
             14'h3d95 	:	val_out <= 16'hff8c;
             14'h3d96 	:	val_out <= 16'hff8d;
             14'h3d97 	:	val_out <= 16'hff8d;
             14'h3d98 	:	val_out <= 16'hff8d;
             14'h3d99 	:	val_out <= 16'hff8e;
             14'h3d9a 	:	val_out <= 16'hff8e;
             14'h3d9b 	:	val_out <= 16'hff8f;
             14'h3d9c 	:	val_out <= 16'hff8f;
             14'h3d9d 	:	val_out <= 16'hff8f;
             14'h3d9e 	:	val_out <= 16'hff90;
             14'h3d9f 	:	val_out <= 16'hff90;
             14'h3da0 	:	val_out <= 16'hff90;
             14'h3da1 	:	val_out <= 16'hff91;
             14'h3da2 	:	val_out <= 16'hff91;
             14'h3da3 	:	val_out <= 16'hff91;
             14'h3da4 	:	val_out <= 16'hff92;
             14'h3da5 	:	val_out <= 16'hff92;
             14'h3da6 	:	val_out <= 16'hff93;
             14'h3da7 	:	val_out <= 16'hff93;
             14'h3da8 	:	val_out <= 16'hff93;
             14'h3da9 	:	val_out <= 16'hff94;
             14'h3daa 	:	val_out <= 16'hff94;
             14'h3dab 	:	val_out <= 16'hff94;
             14'h3dac 	:	val_out <= 16'hff95;
             14'h3dad 	:	val_out <= 16'hff95;
             14'h3dae 	:	val_out <= 16'hff95;
             14'h3daf 	:	val_out <= 16'hff96;
             14'h3db0 	:	val_out <= 16'hff96;
             14'h3db1 	:	val_out <= 16'hff97;
             14'h3db2 	:	val_out <= 16'hff97;
             14'h3db3 	:	val_out <= 16'hff97;
             14'h3db4 	:	val_out <= 16'hff98;
             14'h3db5 	:	val_out <= 16'hff98;
             14'h3db6 	:	val_out <= 16'hff98;
             14'h3db7 	:	val_out <= 16'hff99;
             14'h3db8 	:	val_out <= 16'hff99;
             14'h3db9 	:	val_out <= 16'hff99;
             14'h3dba 	:	val_out <= 16'hff9a;
             14'h3dbb 	:	val_out <= 16'hff9a;
             14'h3dbc 	:	val_out <= 16'hff9a;
             14'h3dbd 	:	val_out <= 16'hff9b;
             14'h3dbe 	:	val_out <= 16'hff9b;
             14'h3dbf 	:	val_out <= 16'hff9b;
             14'h3dc0 	:	val_out <= 16'hff9c;
             14'h3dc1 	:	val_out <= 16'hff9c;
             14'h3dc2 	:	val_out <= 16'hff9c;
             14'h3dc3 	:	val_out <= 16'hff9d;
             14'h3dc4 	:	val_out <= 16'hff9d;
             14'h3dc5 	:	val_out <= 16'hff9d;
             14'h3dc6 	:	val_out <= 16'hff9e;
             14'h3dc7 	:	val_out <= 16'hff9e;
             14'h3dc8 	:	val_out <= 16'hff9f;
             14'h3dc9 	:	val_out <= 16'hff9f;
             14'h3dca 	:	val_out <= 16'hff9f;
             14'h3dcb 	:	val_out <= 16'hffa0;
             14'h3dcc 	:	val_out <= 16'hffa0;
             14'h3dcd 	:	val_out <= 16'hffa0;
             14'h3dce 	:	val_out <= 16'hffa1;
             14'h3dcf 	:	val_out <= 16'hffa1;
             14'h3dd0 	:	val_out <= 16'hffa1;
             14'h3dd1 	:	val_out <= 16'hffa2;
             14'h3dd2 	:	val_out <= 16'hffa2;
             14'h3dd3 	:	val_out <= 16'hffa2;
             14'h3dd4 	:	val_out <= 16'hffa3;
             14'h3dd5 	:	val_out <= 16'hffa3;
             14'h3dd6 	:	val_out <= 16'hffa3;
             14'h3dd7 	:	val_out <= 16'hffa4;
             14'h3dd8 	:	val_out <= 16'hffa4;
             14'h3dd9 	:	val_out <= 16'hffa4;
             14'h3dda 	:	val_out <= 16'hffa5;
             14'h3ddb 	:	val_out <= 16'hffa5;
             14'h3ddc 	:	val_out <= 16'hffa5;
             14'h3ddd 	:	val_out <= 16'hffa6;
             14'h3dde 	:	val_out <= 16'hffa6;
             14'h3ddf 	:	val_out <= 16'hffa6;
             14'h3de0 	:	val_out <= 16'hffa7;
             14'h3de1 	:	val_out <= 16'hffa7;
             14'h3de2 	:	val_out <= 16'hffa7;
             14'h3de3 	:	val_out <= 16'hffa8;
             14'h3de4 	:	val_out <= 16'hffa8;
             14'h3de5 	:	val_out <= 16'hffa8;
             14'h3de6 	:	val_out <= 16'hffa9;
             14'h3de7 	:	val_out <= 16'hffa9;
             14'h3de8 	:	val_out <= 16'hffa9;
             14'h3de9 	:	val_out <= 16'hffa9;
             14'h3dea 	:	val_out <= 16'hffaa;
             14'h3deb 	:	val_out <= 16'hffaa;
             14'h3dec 	:	val_out <= 16'hffaa;
             14'h3ded 	:	val_out <= 16'hffab;
             14'h3dee 	:	val_out <= 16'hffab;
             14'h3def 	:	val_out <= 16'hffab;
             14'h3df0 	:	val_out <= 16'hffac;
             14'h3df1 	:	val_out <= 16'hffac;
             14'h3df2 	:	val_out <= 16'hffac;
             14'h3df3 	:	val_out <= 16'hffad;
             14'h3df4 	:	val_out <= 16'hffad;
             14'h3df5 	:	val_out <= 16'hffad;
             14'h3df6 	:	val_out <= 16'hffae;
             14'h3df7 	:	val_out <= 16'hffae;
             14'h3df8 	:	val_out <= 16'hffae;
             14'h3df9 	:	val_out <= 16'hffaf;
             14'h3dfa 	:	val_out <= 16'hffaf;
             14'h3dfb 	:	val_out <= 16'hffaf;
             14'h3dfc 	:	val_out <= 16'hffaf;
             14'h3dfd 	:	val_out <= 16'hffb0;
             14'h3dfe 	:	val_out <= 16'hffb0;
             14'h3dff 	:	val_out <= 16'hffb0;
             14'h3e00 	:	val_out <= 16'hffb1;
             14'h3e01 	:	val_out <= 16'hffb1;
             14'h3e02 	:	val_out <= 16'hffb1;
             14'h3e03 	:	val_out <= 16'hffb2;
             14'h3e04 	:	val_out <= 16'hffb2;
             14'h3e05 	:	val_out <= 16'hffb2;
             14'h3e06 	:	val_out <= 16'hffb3;
             14'h3e07 	:	val_out <= 16'hffb3;
             14'h3e08 	:	val_out <= 16'hffb3;
             14'h3e09 	:	val_out <= 16'hffb3;
             14'h3e0a 	:	val_out <= 16'hffb4;
             14'h3e0b 	:	val_out <= 16'hffb4;
             14'h3e0c 	:	val_out <= 16'hffb4;
             14'h3e0d 	:	val_out <= 16'hffb5;
             14'h3e0e 	:	val_out <= 16'hffb5;
             14'h3e0f 	:	val_out <= 16'hffb5;
             14'h3e10 	:	val_out <= 16'hffb6;
             14'h3e11 	:	val_out <= 16'hffb6;
             14'h3e12 	:	val_out <= 16'hffb6;
             14'h3e13 	:	val_out <= 16'hffb6;
             14'h3e14 	:	val_out <= 16'hffb7;
             14'h3e15 	:	val_out <= 16'hffb7;
             14'h3e16 	:	val_out <= 16'hffb7;
             14'h3e17 	:	val_out <= 16'hffb8;
             14'h3e18 	:	val_out <= 16'hffb8;
             14'h3e19 	:	val_out <= 16'hffb8;
             14'h3e1a 	:	val_out <= 16'hffb9;
             14'h3e1b 	:	val_out <= 16'hffb9;
             14'h3e1c 	:	val_out <= 16'hffb9;
             14'h3e1d 	:	val_out <= 16'hffb9;
             14'h3e1e 	:	val_out <= 16'hffba;
             14'h3e1f 	:	val_out <= 16'hffba;
             14'h3e20 	:	val_out <= 16'hffba;
             14'h3e21 	:	val_out <= 16'hffbb;
             14'h3e22 	:	val_out <= 16'hffbb;
             14'h3e23 	:	val_out <= 16'hffbb;
             14'h3e24 	:	val_out <= 16'hffbb;
             14'h3e25 	:	val_out <= 16'hffbc;
             14'h3e26 	:	val_out <= 16'hffbc;
             14'h3e27 	:	val_out <= 16'hffbc;
             14'h3e28 	:	val_out <= 16'hffbd;
             14'h3e29 	:	val_out <= 16'hffbd;
             14'h3e2a 	:	val_out <= 16'hffbd;
             14'h3e2b 	:	val_out <= 16'hffbd;
             14'h3e2c 	:	val_out <= 16'hffbe;
             14'h3e2d 	:	val_out <= 16'hffbe;
             14'h3e2e 	:	val_out <= 16'hffbe;
             14'h3e2f 	:	val_out <= 16'hffbf;
             14'h3e30 	:	val_out <= 16'hffbf;
             14'h3e31 	:	val_out <= 16'hffbf;
             14'h3e32 	:	val_out <= 16'hffbf;
             14'h3e33 	:	val_out <= 16'hffc0;
             14'h3e34 	:	val_out <= 16'hffc0;
             14'h3e35 	:	val_out <= 16'hffc0;
             14'h3e36 	:	val_out <= 16'hffc0;
             14'h3e37 	:	val_out <= 16'hffc1;
             14'h3e38 	:	val_out <= 16'hffc1;
             14'h3e39 	:	val_out <= 16'hffc1;
             14'h3e3a 	:	val_out <= 16'hffc2;
             14'h3e3b 	:	val_out <= 16'hffc2;
             14'h3e3c 	:	val_out <= 16'hffc2;
             14'h3e3d 	:	val_out <= 16'hffc2;
             14'h3e3e 	:	val_out <= 16'hffc3;
             14'h3e3f 	:	val_out <= 16'hffc3;
             14'h3e40 	:	val_out <= 16'hffc3;
             14'h3e41 	:	val_out <= 16'hffc3;
             14'h3e42 	:	val_out <= 16'hffc4;
             14'h3e43 	:	val_out <= 16'hffc4;
             14'h3e44 	:	val_out <= 16'hffc4;
             14'h3e45 	:	val_out <= 16'hffc5;
             14'h3e46 	:	val_out <= 16'hffc5;
             14'h3e47 	:	val_out <= 16'hffc5;
             14'h3e48 	:	val_out <= 16'hffc5;
             14'h3e49 	:	val_out <= 16'hffc6;
             14'h3e4a 	:	val_out <= 16'hffc6;
             14'h3e4b 	:	val_out <= 16'hffc6;
             14'h3e4c 	:	val_out <= 16'hffc6;
             14'h3e4d 	:	val_out <= 16'hffc7;
             14'h3e4e 	:	val_out <= 16'hffc7;
             14'h3e4f 	:	val_out <= 16'hffc7;
             14'h3e50 	:	val_out <= 16'hffc7;
             14'h3e51 	:	val_out <= 16'hffc8;
             14'h3e52 	:	val_out <= 16'hffc8;
             14'h3e53 	:	val_out <= 16'hffc8;
             14'h3e54 	:	val_out <= 16'hffc8;
             14'h3e55 	:	val_out <= 16'hffc9;
             14'h3e56 	:	val_out <= 16'hffc9;
             14'h3e57 	:	val_out <= 16'hffc9;
             14'h3e58 	:	val_out <= 16'hffc9;
             14'h3e59 	:	val_out <= 16'hffca;
             14'h3e5a 	:	val_out <= 16'hffca;
             14'h3e5b 	:	val_out <= 16'hffca;
             14'h3e5c 	:	val_out <= 16'hffcb;
             14'h3e5d 	:	val_out <= 16'hffcb;
             14'h3e5e 	:	val_out <= 16'hffcb;
             14'h3e5f 	:	val_out <= 16'hffcb;
             14'h3e60 	:	val_out <= 16'hffcc;
             14'h3e61 	:	val_out <= 16'hffcc;
             14'h3e62 	:	val_out <= 16'hffcc;
             14'h3e63 	:	val_out <= 16'hffcc;
             14'h3e64 	:	val_out <= 16'hffcd;
             14'h3e65 	:	val_out <= 16'hffcd;
             14'h3e66 	:	val_out <= 16'hffcd;
             14'h3e67 	:	val_out <= 16'hffcd;
             14'h3e68 	:	val_out <= 16'hffcd;
             14'h3e69 	:	val_out <= 16'hffce;
             14'h3e6a 	:	val_out <= 16'hffce;
             14'h3e6b 	:	val_out <= 16'hffce;
             14'h3e6c 	:	val_out <= 16'hffce;
             14'h3e6d 	:	val_out <= 16'hffcf;
             14'h3e6e 	:	val_out <= 16'hffcf;
             14'h3e6f 	:	val_out <= 16'hffcf;
             14'h3e70 	:	val_out <= 16'hffcf;
             14'h3e71 	:	val_out <= 16'hffd0;
             14'h3e72 	:	val_out <= 16'hffd0;
             14'h3e73 	:	val_out <= 16'hffd0;
             14'h3e74 	:	val_out <= 16'hffd0;
             14'h3e75 	:	val_out <= 16'hffd1;
             14'h3e76 	:	val_out <= 16'hffd1;
             14'h3e77 	:	val_out <= 16'hffd1;
             14'h3e78 	:	val_out <= 16'hffd1;
             14'h3e79 	:	val_out <= 16'hffd2;
             14'h3e7a 	:	val_out <= 16'hffd2;
             14'h3e7b 	:	val_out <= 16'hffd2;
             14'h3e7c 	:	val_out <= 16'hffd2;
             14'h3e7d 	:	val_out <= 16'hffd3;
             14'h3e7e 	:	val_out <= 16'hffd3;
             14'h3e7f 	:	val_out <= 16'hffd3;
             14'h3e80 	:	val_out <= 16'hffd3;
             14'h3e81 	:	val_out <= 16'hffd3;
             14'h3e82 	:	val_out <= 16'hffd4;
             14'h3e83 	:	val_out <= 16'hffd4;
             14'h3e84 	:	val_out <= 16'hffd4;
             14'h3e85 	:	val_out <= 16'hffd4;
             14'h3e86 	:	val_out <= 16'hffd5;
             14'h3e87 	:	val_out <= 16'hffd5;
             14'h3e88 	:	val_out <= 16'hffd5;
             14'h3e89 	:	val_out <= 16'hffd5;
             14'h3e8a 	:	val_out <= 16'hffd5;
             14'h3e8b 	:	val_out <= 16'hffd6;
             14'h3e8c 	:	val_out <= 16'hffd6;
             14'h3e8d 	:	val_out <= 16'hffd6;
             14'h3e8e 	:	val_out <= 16'hffd6;
             14'h3e8f 	:	val_out <= 16'hffd7;
             14'h3e90 	:	val_out <= 16'hffd7;
             14'h3e91 	:	val_out <= 16'hffd7;
             14'h3e92 	:	val_out <= 16'hffd7;
             14'h3e93 	:	val_out <= 16'hffd7;
             14'h3e94 	:	val_out <= 16'hffd8;
             14'h3e95 	:	val_out <= 16'hffd8;
             14'h3e96 	:	val_out <= 16'hffd8;
             14'h3e97 	:	val_out <= 16'hffd8;
             14'h3e98 	:	val_out <= 16'hffd9;
             14'h3e99 	:	val_out <= 16'hffd9;
             14'h3e9a 	:	val_out <= 16'hffd9;
             14'h3e9b 	:	val_out <= 16'hffd9;
             14'h3e9c 	:	val_out <= 16'hffd9;
             14'h3e9d 	:	val_out <= 16'hffda;
             14'h3e9e 	:	val_out <= 16'hffda;
             14'h3e9f 	:	val_out <= 16'hffda;
             14'h3ea0 	:	val_out <= 16'hffda;
             14'h3ea1 	:	val_out <= 16'hffdb;
             14'h3ea2 	:	val_out <= 16'hffdb;
             14'h3ea3 	:	val_out <= 16'hffdb;
             14'h3ea4 	:	val_out <= 16'hffdb;
             14'h3ea5 	:	val_out <= 16'hffdb;
             14'h3ea6 	:	val_out <= 16'hffdc;
             14'h3ea7 	:	val_out <= 16'hffdc;
             14'h3ea8 	:	val_out <= 16'hffdc;
             14'h3ea9 	:	val_out <= 16'hffdc;
             14'h3eaa 	:	val_out <= 16'hffdc;
             14'h3eab 	:	val_out <= 16'hffdd;
             14'h3eac 	:	val_out <= 16'hffdd;
             14'h3ead 	:	val_out <= 16'hffdd;
             14'h3eae 	:	val_out <= 16'hffdd;
             14'h3eaf 	:	val_out <= 16'hffdd;
             14'h3eb0 	:	val_out <= 16'hffde;
             14'h3eb1 	:	val_out <= 16'hffde;
             14'h3eb2 	:	val_out <= 16'hffde;
             14'h3eb3 	:	val_out <= 16'hffde;
             14'h3eb4 	:	val_out <= 16'hffde;
             14'h3eb5 	:	val_out <= 16'hffdf;
             14'h3eb6 	:	val_out <= 16'hffdf;
             14'h3eb7 	:	val_out <= 16'hffdf;
             14'h3eb8 	:	val_out <= 16'hffdf;
             14'h3eb9 	:	val_out <= 16'hffdf;
             14'h3eba 	:	val_out <= 16'hffe0;
             14'h3ebb 	:	val_out <= 16'hffe0;
             14'h3ebc 	:	val_out <= 16'hffe0;
             14'h3ebd 	:	val_out <= 16'hffe0;
             14'h3ebe 	:	val_out <= 16'hffe0;
             14'h3ebf 	:	val_out <= 16'hffe1;
             14'h3ec0 	:	val_out <= 16'hffe1;
             14'h3ec1 	:	val_out <= 16'hffe1;
             14'h3ec2 	:	val_out <= 16'hffe1;
             14'h3ec3 	:	val_out <= 16'hffe1;
             14'h3ec4 	:	val_out <= 16'hffe2;
             14'h3ec5 	:	val_out <= 16'hffe2;
             14'h3ec6 	:	val_out <= 16'hffe2;
             14'h3ec7 	:	val_out <= 16'hffe2;
             14'h3ec8 	:	val_out <= 16'hffe2;
             14'h3ec9 	:	val_out <= 16'hffe2;
             14'h3eca 	:	val_out <= 16'hffe3;
             14'h3ecb 	:	val_out <= 16'hffe3;
             14'h3ecc 	:	val_out <= 16'hffe3;
             14'h3ecd 	:	val_out <= 16'hffe3;
             14'h3ece 	:	val_out <= 16'hffe3;
             14'h3ecf 	:	val_out <= 16'hffe4;
             14'h3ed0 	:	val_out <= 16'hffe4;
             14'h3ed1 	:	val_out <= 16'hffe4;
             14'h3ed2 	:	val_out <= 16'hffe4;
             14'h3ed3 	:	val_out <= 16'hffe4;
             14'h3ed4 	:	val_out <= 16'hffe4;
             14'h3ed5 	:	val_out <= 16'hffe5;
             14'h3ed6 	:	val_out <= 16'hffe5;
             14'h3ed7 	:	val_out <= 16'hffe5;
             14'h3ed8 	:	val_out <= 16'hffe5;
             14'h3ed9 	:	val_out <= 16'hffe5;
             14'h3eda 	:	val_out <= 16'hffe6;
             14'h3edb 	:	val_out <= 16'hffe6;
             14'h3edc 	:	val_out <= 16'hffe6;
             14'h3edd 	:	val_out <= 16'hffe6;
             14'h3ede 	:	val_out <= 16'hffe6;
             14'h3edf 	:	val_out <= 16'hffe6;
             14'h3ee0 	:	val_out <= 16'hffe7;
             14'h3ee1 	:	val_out <= 16'hffe7;
             14'h3ee2 	:	val_out <= 16'hffe7;
             14'h3ee3 	:	val_out <= 16'hffe7;
             14'h3ee4 	:	val_out <= 16'hffe7;
             14'h3ee5 	:	val_out <= 16'hffe7;
             14'h3ee6 	:	val_out <= 16'hffe8;
             14'h3ee7 	:	val_out <= 16'hffe8;
             14'h3ee8 	:	val_out <= 16'hffe8;
             14'h3ee9 	:	val_out <= 16'hffe8;
             14'h3eea 	:	val_out <= 16'hffe8;
             14'h3eeb 	:	val_out <= 16'hffe8;
             14'h3eec 	:	val_out <= 16'hffe9;
             14'h3eed 	:	val_out <= 16'hffe9;
             14'h3eee 	:	val_out <= 16'hffe9;
             14'h3eef 	:	val_out <= 16'hffe9;
             14'h3ef0 	:	val_out <= 16'hffe9;
             14'h3ef1 	:	val_out <= 16'hffe9;
             14'h3ef2 	:	val_out <= 16'hffea;
             14'h3ef3 	:	val_out <= 16'hffea;
             14'h3ef4 	:	val_out <= 16'hffea;
             14'h3ef5 	:	val_out <= 16'hffea;
             14'h3ef6 	:	val_out <= 16'hffea;
             14'h3ef7 	:	val_out <= 16'hffea;
             14'h3ef8 	:	val_out <= 16'hffeb;
             14'h3ef9 	:	val_out <= 16'hffeb;
             14'h3efa 	:	val_out <= 16'hffeb;
             14'h3efb 	:	val_out <= 16'hffeb;
             14'h3efc 	:	val_out <= 16'hffeb;
             14'h3efd 	:	val_out <= 16'hffeb;
             14'h3efe 	:	val_out <= 16'hffec;
             14'h3eff 	:	val_out <= 16'hffec;
             14'h3f00 	:	val_out <= 16'hffec;
             14'h3f01 	:	val_out <= 16'hffec;
             14'h3f02 	:	val_out <= 16'hffec;
             14'h3f03 	:	val_out <= 16'hffec;
             14'h3f04 	:	val_out <= 16'hffec;
             14'h3f05 	:	val_out <= 16'hffed;
             14'h3f06 	:	val_out <= 16'hffed;
             14'h3f07 	:	val_out <= 16'hffed;
             14'h3f08 	:	val_out <= 16'hffed;
             14'h3f09 	:	val_out <= 16'hffed;
             14'h3f0a 	:	val_out <= 16'hffed;
             14'h3f0b 	:	val_out <= 16'hffed;
             14'h3f0c 	:	val_out <= 16'hffee;
             14'h3f0d 	:	val_out <= 16'hffee;
             14'h3f0e 	:	val_out <= 16'hffee;
             14'h3f0f 	:	val_out <= 16'hffee;
             14'h3f10 	:	val_out <= 16'hffee;
             14'h3f11 	:	val_out <= 16'hffee;
             14'h3f12 	:	val_out <= 16'hffef;
             14'h3f13 	:	val_out <= 16'hffef;
             14'h3f14 	:	val_out <= 16'hffef;
             14'h3f15 	:	val_out <= 16'hffef;
             14'h3f16 	:	val_out <= 16'hffef;
             14'h3f17 	:	val_out <= 16'hffef;
             14'h3f18 	:	val_out <= 16'hffef;
             14'h3f19 	:	val_out <= 16'hffef;
             14'h3f1a 	:	val_out <= 16'hfff0;
             14'h3f1b 	:	val_out <= 16'hfff0;
             14'h3f1c 	:	val_out <= 16'hfff0;
             14'h3f1d 	:	val_out <= 16'hfff0;
             14'h3f1e 	:	val_out <= 16'hfff0;
             14'h3f1f 	:	val_out <= 16'hfff0;
             14'h3f20 	:	val_out <= 16'hfff0;
             14'h3f21 	:	val_out <= 16'hfff1;
             14'h3f22 	:	val_out <= 16'hfff1;
             14'h3f23 	:	val_out <= 16'hfff1;
             14'h3f24 	:	val_out <= 16'hfff1;
             14'h3f25 	:	val_out <= 16'hfff1;
             14'h3f26 	:	val_out <= 16'hfff1;
             14'h3f27 	:	val_out <= 16'hfff1;
             14'h3f28 	:	val_out <= 16'hfff2;
             14'h3f29 	:	val_out <= 16'hfff2;
             14'h3f2a 	:	val_out <= 16'hfff2;
             14'h3f2b 	:	val_out <= 16'hfff2;
             14'h3f2c 	:	val_out <= 16'hfff2;
             14'h3f2d 	:	val_out <= 16'hfff2;
             14'h3f2e 	:	val_out <= 16'hfff2;
             14'h3f2f 	:	val_out <= 16'hfff2;
             14'h3f30 	:	val_out <= 16'hfff3;
             14'h3f31 	:	val_out <= 16'hfff3;
             14'h3f32 	:	val_out <= 16'hfff3;
             14'h3f33 	:	val_out <= 16'hfff3;
             14'h3f34 	:	val_out <= 16'hfff3;
             14'h3f35 	:	val_out <= 16'hfff3;
             14'h3f36 	:	val_out <= 16'hfff3;
             14'h3f37 	:	val_out <= 16'hfff3;
             14'h3f38 	:	val_out <= 16'hfff4;
             14'h3f39 	:	val_out <= 16'hfff4;
             14'h3f3a 	:	val_out <= 16'hfff4;
             14'h3f3b 	:	val_out <= 16'hfff4;
             14'h3f3c 	:	val_out <= 16'hfff4;
             14'h3f3d 	:	val_out <= 16'hfff4;
             14'h3f3e 	:	val_out <= 16'hfff4;
             14'h3f3f 	:	val_out <= 16'hfff4;
             14'h3f40 	:	val_out <= 16'hfff4;
             14'h3f41 	:	val_out <= 16'hfff5;
             14'h3f42 	:	val_out <= 16'hfff5;
             14'h3f43 	:	val_out <= 16'hfff5;
             14'h3f44 	:	val_out <= 16'hfff5;
             14'h3f45 	:	val_out <= 16'hfff5;
             14'h3f46 	:	val_out <= 16'hfff5;
             14'h3f47 	:	val_out <= 16'hfff5;
             14'h3f48 	:	val_out <= 16'hfff5;
             14'h3f49 	:	val_out <= 16'hfff5;
             14'h3f4a 	:	val_out <= 16'hfff6;
             14'h3f4b 	:	val_out <= 16'hfff6;
             14'h3f4c 	:	val_out <= 16'hfff6;
             14'h3f4d 	:	val_out <= 16'hfff6;
             14'h3f4e 	:	val_out <= 16'hfff6;
             14'h3f4f 	:	val_out <= 16'hfff6;
             14'h3f50 	:	val_out <= 16'hfff6;
             14'h3f51 	:	val_out <= 16'hfff6;
             14'h3f52 	:	val_out <= 16'hfff6;
             14'h3f53 	:	val_out <= 16'hfff7;
             14'h3f54 	:	val_out <= 16'hfff7;
             14'h3f55 	:	val_out <= 16'hfff7;
             14'h3f56 	:	val_out <= 16'hfff7;
             14'h3f57 	:	val_out <= 16'hfff7;
             14'h3f58 	:	val_out <= 16'hfff7;
             14'h3f59 	:	val_out <= 16'hfff7;
             14'h3f5a 	:	val_out <= 16'hfff7;
             14'h3f5b 	:	val_out <= 16'hfff7;
             14'h3f5c 	:	val_out <= 16'hfff7;
             14'h3f5d 	:	val_out <= 16'hfff8;
             14'h3f5e 	:	val_out <= 16'hfff8;
             14'h3f5f 	:	val_out <= 16'hfff8;
             14'h3f60 	:	val_out <= 16'hfff8;
             14'h3f61 	:	val_out <= 16'hfff8;
             14'h3f62 	:	val_out <= 16'hfff8;
             14'h3f63 	:	val_out <= 16'hfff8;
             14'h3f64 	:	val_out <= 16'hfff8;
             14'h3f65 	:	val_out <= 16'hfff8;
             14'h3f66 	:	val_out <= 16'hfff8;
             14'h3f67 	:	val_out <= 16'hfff8;
             14'h3f68 	:	val_out <= 16'hfff9;
             14'h3f69 	:	val_out <= 16'hfff9;
             14'h3f6a 	:	val_out <= 16'hfff9;
             14'h3f6b 	:	val_out <= 16'hfff9;
             14'h3f6c 	:	val_out <= 16'hfff9;
             14'h3f6d 	:	val_out <= 16'hfff9;
             14'h3f6e 	:	val_out <= 16'hfff9;
             14'h3f6f 	:	val_out <= 16'hfff9;
             14'h3f70 	:	val_out <= 16'hfff9;
             14'h3f71 	:	val_out <= 16'hfff9;
             14'h3f72 	:	val_out <= 16'hfff9;
             14'h3f73 	:	val_out <= 16'hfffa;
             14'h3f74 	:	val_out <= 16'hfffa;
             14'h3f75 	:	val_out <= 16'hfffa;
             14'h3f76 	:	val_out <= 16'hfffa;
             14'h3f77 	:	val_out <= 16'hfffa;
             14'h3f78 	:	val_out <= 16'hfffa;
             14'h3f79 	:	val_out <= 16'hfffa;
             14'h3f7a 	:	val_out <= 16'hfffa;
             14'h3f7b 	:	val_out <= 16'hfffa;
             14'h3f7c 	:	val_out <= 16'hfffa;
             14'h3f7d 	:	val_out <= 16'hfffa;
             14'h3f7e 	:	val_out <= 16'hfffa;
             14'h3f7f 	:	val_out <= 16'hfffb;
             14'h3f80 	:	val_out <= 16'hfffb;
             14'h3f81 	:	val_out <= 16'hfffb;
             14'h3f82 	:	val_out <= 16'hfffb;
             14'h3f83 	:	val_out <= 16'hfffb;
             14'h3f84 	:	val_out <= 16'hfffb;
             14'h3f85 	:	val_out <= 16'hfffb;
             14'h3f86 	:	val_out <= 16'hfffb;
             14'h3f87 	:	val_out <= 16'hfffb;
             14'h3f88 	:	val_out <= 16'hfffb;
             14'h3f89 	:	val_out <= 16'hfffb;
             14'h3f8a 	:	val_out <= 16'hfffb;
             14'h3f8b 	:	val_out <= 16'hfffb;
             14'h3f8c 	:	val_out <= 16'hfffb;
             14'h3f8d 	:	val_out <= 16'hfffc;
             14'h3f8e 	:	val_out <= 16'hfffc;
             14'h3f8f 	:	val_out <= 16'hfffc;
             14'h3f90 	:	val_out <= 16'hfffc;
             14'h3f91 	:	val_out <= 16'hfffc;
             14'h3f92 	:	val_out <= 16'hfffc;
             14'h3f93 	:	val_out <= 16'hfffc;
             14'h3f94 	:	val_out <= 16'hfffc;
             14'h3f95 	:	val_out <= 16'hfffc;
             14'h3f96 	:	val_out <= 16'hfffc;
             14'h3f97 	:	val_out <= 16'hfffc;
             14'h3f98 	:	val_out <= 16'hfffc;
             14'h3f99 	:	val_out <= 16'hfffc;
             14'h3f9a 	:	val_out <= 16'hfffc;
             14'h3f9b 	:	val_out <= 16'hfffc;
             14'h3f9c 	:	val_out <= 16'hfffd;
             14'h3f9d 	:	val_out <= 16'hfffd;
             14'h3f9e 	:	val_out <= 16'hfffd;
             14'h3f9f 	:	val_out <= 16'hfffd;
             14'h3fa0 	:	val_out <= 16'hfffd;
             14'h3fa1 	:	val_out <= 16'hfffd;
             14'h3fa2 	:	val_out <= 16'hfffd;
             14'h3fa3 	:	val_out <= 16'hfffd;
             14'h3fa4 	:	val_out <= 16'hfffd;
             14'h3fa5 	:	val_out <= 16'hfffd;
             14'h3fa6 	:	val_out <= 16'hfffd;
             14'h3fa7 	:	val_out <= 16'hfffd;
             14'h3fa8 	:	val_out <= 16'hfffd;
             14'h3fa9 	:	val_out <= 16'hfffd;
             14'h3faa 	:	val_out <= 16'hfffd;
             14'h3fab 	:	val_out <= 16'hfffd;
             14'h3fac 	:	val_out <= 16'hfffd;
             14'h3fad 	:	val_out <= 16'hfffd;
             14'h3fae 	:	val_out <= 16'hfffd;
             14'h3faf 	:	val_out <= 16'hfffe;
             14'h3fb0 	:	val_out <= 16'hfffe;
             14'h3fb1 	:	val_out <= 16'hfffe;
             14'h3fb2 	:	val_out <= 16'hfffe;
             14'h3fb3 	:	val_out <= 16'hfffe;
             14'h3fb4 	:	val_out <= 16'hfffe;
             14'h3fb5 	:	val_out <= 16'hfffe;
             14'h3fb6 	:	val_out <= 16'hfffe;
             14'h3fb7 	:	val_out <= 16'hfffe;
             14'h3fb8 	:	val_out <= 16'hfffe;
             14'h3fb9 	:	val_out <= 16'hfffe;
             14'h3fba 	:	val_out <= 16'hfffe;
             14'h3fbb 	:	val_out <= 16'hfffe;
             14'h3fbc 	:	val_out <= 16'hfffe;
             14'h3fbd 	:	val_out <= 16'hfffe;
             14'h3fbe 	:	val_out <= 16'hfffe;
             14'h3fbf 	:	val_out <= 16'hfffe;
             14'h3fc0 	:	val_out <= 16'hfffe;
             14'h3fc1 	:	val_out <= 16'hfffe;
             14'h3fc2 	:	val_out <= 16'hfffe;
             14'h3fc3 	:	val_out <= 16'hfffe;
             14'h3fc4 	:	val_out <= 16'hfffe;
             14'h3fc5 	:	val_out <= 16'hfffe;
             14'h3fc6 	:	val_out <= 16'hffff;
             14'h3fc7 	:	val_out <= 16'hffff;
             14'h3fc8 	:	val_out <= 16'hffff;
             14'h3fc9 	:	val_out <= 16'hffff;
             14'h3fca 	:	val_out <= 16'hffff;
             14'h3fcb 	:	val_out <= 16'hffff;
             14'h3fcc 	:	val_out <= 16'hffff;
             14'h3fcd 	:	val_out <= 16'hffff;
             14'h3fce 	:	val_out <= 16'hffff;
             14'h3fcf 	:	val_out <= 16'hffff;
             14'h3fd0 	:	val_out <= 16'hffff;
             14'h3fd1 	:	val_out <= 16'hffff;
             14'h3fd2 	:	val_out <= 16'hffff;
             14'h3fd3 	:	val_out <= 16'hffff;
             14'h3fd4 	:	val_out <= 16'hffff;
             14'h3fd5 	:	val_out <= 16'hffff;
             14'h3fd6 	:	val_out <= 16'hffff;
             14'h3fd7 	:	val_out <= 16'hffff;
             14'h3fd8 	:	val_out <= 16'hffff;
             14'h3fd9 	:	val_out <= 16'hffff;
             14'h3fda 	:	val_out <= 16'hffff;
             14'h3fdb 	:	val_out <= 16'hffff;
             14'h3fdc 	:	val_out <= 16'hffff;
             14'h3fdd 	:	val_out <= 16'hffff;
             14'h3fde 	:	val_out <= 16'hffff;
             14'h3fdf 	:	val_out <= 16'hffff;
             14'h3fe0 	:	val_out <= 16'hffff;
             14'h3fe1 	:	val_out <= 16'hffff;
             14'h3fe2 	:	val_out <= 16'hffff;
             14'h3fe3 	:	val_out <= 16'hffff;
             14'h3fe4 	:	val_out <= 16'hffff;
             14'h3fe5 	:	val_out <= 16'hffff;
             14'h3fe6 	:	val_out <= 16'hffff;
             14'h3fe7 	:	val_out <= 16'hffff;
             14'h3fe8 	:	val_out <= 16'hffff;
             14'h3fe9 	:	val_out <= 16'hffff;
             14'h3fea 	:	val_out <= 16'hffff;
             14'h3feb 	:	val_out <= 16'hffff;
             14'h3fec 	:	val_out <= 16'hffff;
             14'h3fed 	:	val_out <= 16'hffff;
             14'h3fee 	:	val_out <= 16'hffff;
             14'h3fef 	:	val_out <= 16'hffff;
             14'h3ff0 	:	val_out <= 16'hffff;
             14'h3ff1 	:	val_out <= 16'hffff;
             14'h3ff2 	:	val_out <= 16'hffff;
             14'h3ff3 	:	val_out <= 16'hffff;
             14'h3ff4 	:	val_out <= 16'hffff;
             14'h3ff5 	:	val_out <= 16'hffff;
             14'h3ff6 	:	val_out <= 16'hffff;
             14'h3ff7 	:	val_out <= 16'hffff;
             14'h3ff8 	:	val_out <= 16'hffff;
             14'h3ff9 	:	val_out <= 16'hffff;
             14'h3ffa 	:	val_out <= 16'hffff;
             14'h3ffb 	:	val_out <= 16'hffff;
             14'h3ffc 	:	val_out <= 16'hffff;
             14'h3ffd 	:	val_out <= 16'hffff;
             14'h3ffe 	:	val_out <= 16'hffff;
             14'h3fff 	:	val_out <= 16'hffff;
				 default		:	val_out <= 16'h0000;
			endcase
		end
endmodule
								
