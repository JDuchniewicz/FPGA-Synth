// Pipelined phase bank module

module phase_bank_p(input clk,
						input clk_en,
						input rst,
						input[6:0] i_midi,
						output reg[6:0] o_midi,
						output reg o_valid, 
						output reg[23:0] o_phase);
		parameter NBANKS = 10;
		
		// for now holding 24 bits, feeding LUT with only 16 upper bits of bank -> losing precision but frequency should be right
		// if want make phase interpolation then need to output both integer and fractional part then interpolate in sine
		reg[23:0] phase_banks[NBANKS-1:0];
		wire[23:0] w_tw;
		
		tuning_word_lut tw_lut(.i_midi(i_midi), .o_tw(w_tw));
		
		integer v_idx;
		integer i;
		
		initial begin
			o_phase = 16'b0;
			v_idx = 9;
			for (i = 0; i < NBANKS; i = i + 1) begin
				phase_banks[i] = 24'b0;
			end
			o_midi = 7'b0;
		end
		
		always @(posedge clk or posedge rst) begin
			if (rst) begin
				o_phase = 16'b0;
				v_idx = 9;
				for (i = 0; i < NBANKS; i = i + 1) begin
					phase_banks[i] <= 24'b0;
				end
				o_midi <= 7'b0;
			end else if (clk_en) begin
				if (i_midi !== 7'h0) begin
					phase_banks[v_idx] <= phase_banks[v_idx] + w_tw;
					o_phase <= phase_banks[v_idx]; // output a delayed value (one whole loop)
				end else begin
					o_phase <= 16'b0;
				end
					
				o_valid <= (i_midi == 7'h0) ? 1'b0 : 1'b1;
				o_midi <= i_midi;
				
				if (v_idx == NBANKS - 1)
					v_idx <= 0;
				else
					v_idx <= v_idx + 1;
			end
		end
						
endmodule

// right now increasing tw to 24 bits
module tuning_word_lut(input[6:0] i_midi,
								output reg[23:0] o_tw);
		initial o_tw = 24'b0;
		
		always @(i_midi) begin
			case(i_midi)
            7'h00 	:	o_tw <= 24'b000000000000000000001101;
            7'h01 	:	o_tw <= 24'b000000000000000000001110;
            7'h02 	:	o_tw <= 24'b000000000000000000001111;
            7'h03 	:	o_tw <= 24'b000000000000000000010000;
            7'h04 	:	o_tw <= 24'b000000000000000000010001;
            7'h05 	:	o_tw <= 24'b000000000000000000010010;
            7'h06 	:	o_tw <= 24'b000000000000000000010011;
            7'h07 	:	o_tw <= 24'b000000000000000000010100;
            7'h08 	:	o_tw <= 24'b000000000000000000010101;
            7'h09 	:	o_tw <= 24'b000000000000000000010111;
            7'h0a 	:	o_tw <= 24'b000000000000000000011000;
            7'h0b 	:	o_tw <= 24'b000000000000000000011001;
            7'h0c 	:	o_tw <= 24'b000000000000000000011011;
            7'h0d 	:	o_tw <= 24'b000000000000000000011101;
            7'h0e 	:	o_tw <= 24'b000000000000000000011110;
            7'h0f 	:	o_tw <= 24'b000000000000000000100000;
            7'h10 	:	o_tw <= 24'b000000000000000000100010;
            7'h11 	:	o_tw <= 24'b000000000000000000100100;
            7'h12 	:	o_tw <= 24'b000000000000000000100110;
            7'h13 	:	o_tw <= 24'b000000000000000000101001;
            7'h14 	:	o_tw <= 24'b000000000000000000101011;
            7'h15 	:	o_tw <= 24'b000000000000000000101110;
            7'h16 	:	o_tw <= 24'b000000000000000000110000;
            7'h17 	:	o_tw <= 24'b000000000000000000110011;
            7'h18 	:	o_tw <= 24'b000000000000000000110110;
            7'h19 	:	o_tw <= 24'b000000000000000000111010;
            7'h1a 	:	o_tw <= 24'b000000000000000000111101;
            7'h1b 	:	o_tw <= 24'b000000000000000001000001;
            7'h1c 	:	o_tw <= 24'b000000000000000001000101;
            7'h1d 	:	o_tw <= 24'b000000000000000001001001;
            7'h1e 	:	o_tw <= 24'b000000000000000001001101;
            7'h1f 	:	o_tw <= 24'b000000000000000001010010;
            7'h20 	:	o_tw <= 24'b000000000000000001010111;
            7'h21 	:	o_tw <= 24'b000000000000000001011100;
            7'h22 	:	o_tw <= 24'b000000000000000001100001;
            7'h23 	:	o_tw <= 24'b000000000000000001100111;
            7'h24 	:	o_tw <= 24'b000000000000000001101101;
            7'h25 	:	o_tw <= 24'b000000000000000001110100;
            7'h26 	:	o_tw <= 24'b000000000000000001111011;
            7'h27 	:	o_tw <= 24'b000000000000000010000010;
            7'h28 	:	o_tw <= 24'b000000000000000010001010;
            7'h29 	:	o_tw <= 24'b000000000000000010010010;
            7'h2a 	:	o_tw <= 24'b000000000000000010011011;
            7'h2b 	:	o_tw <= 24'b000000000000000010100100;
            7'h2c 	:	o_tw <= 24'b000000000000000010101110;
            7'h2d 	:	o_tw <= 24'b000000000000000010111000;
            7'h2e 	:	o_tw <= 24'b000000000000000011000011;
            7'h2f 	:	o_tw <= 24'b000000000000000011001111;
            7'h30 	:	o_tw <= 24'b000000000000000011011011;
            7'h31 	:	o_tw <= 24'b000000000000000011101000;
            7'h32 	:	o_tw <= 24'b000000000000000011110110;
            7'h33 	:	o_tw <= 24'b000000000000000100000100;
            7'h34 	:	o_tw <= 24'b000000000000000100010100;
            7'h35 	:	o_tw <= 24'b000000000000000100100100;
            7'h36 	:	o_tw <= 24'b000000000000000100110110;
            7'h37 	:	o_tw <= 24'b000000000000000101001000;
            7'h38 	:	o_tw <= 24'b000000000000000101011100;
            7'h39 	:	o_tw <= 24'b000000000000000101110001;
            7'h3a 	:	o_tw <= 24'b000000000000000110000111;
            7'h3b 	:	o_tw <= 24'b000000000000000110011110;
            7'h3c 	:	o_tw <= 24'b000000000000000110110110;
            7'h3d 	:	o_tw <= 24'b000000000000000111010001;
            7'h3e 	:	o_tw <= 24'b000000000000000111101100;
            7'h3f 	:	o_tw <= 24'b000000000000001000001001;
            7'h40 	:	o_tw <= 24'b000000000000001000101001;
            7'h41 	:	o_tw <= 24'b000000000000001001001001;
            7'h42 	:	o_tw <= 24'b000000000000001001101100;
            7'h43 	:	o_tw <= 24'b000000000000001010010001;
            7'h44 	:	o_tw <= 24'b000000000000001010111000;
            7'h45 	:	o_tw <= 24'b000000000000001011100010;
            7'h46 	:	o_tw <= 24'b000000000000001100001110;
            7'h47 	:	o_tw <= 24'b000000000000001100111100;
            7'h48 	:	o_tw <= 24'b000000000000001101101101;
            7'h49 	:	o_tw <= 24'b000000000000001110100010;
            7'h4a 	:	o_tw <= 24'b000000000000001111011001;
            7'h4b 	:	o_tw <= 24'b000000000000010000010011;
            7'h4c 	:	o_tw <= 24'b000000000000010001010010;
            7'h4d 	:	o_tw <= 24'b000000000000010010010011;
            7'h4e 	:	o_tw <= 24'b000000000000010011011001;
            7'h4f 	:	o_tw <= 24'b000000000000010100100011;
            7'h50 	:	o_tw <= 24'b000000000000010101110001;
            7'h51 	:	o_tw <= 24'b000000000000010111000100;
            7'h52 	:	o_tw <= 24'b000000000000011000011100;
            7'h53 	:	o_tw <= 24'b000000000000011001111001;
            7'h54 	:	o_tw <= 24'b000000000000011011011011;
            7'h55 	:	o_tw <= 24'b000000000000011101000100;
            7'h56 	:	o_tw <= 24'b000000000000011110110010;
            7'h57 	:	o_tw <= 24'b000000000000100000100111;
            7'h58 	:	o_tw <= 24'b000000000000100010100100;
            7'h59 	:	o_tw <= 24'b000000000000100100100111;
            7'h5a 	:	o_tw <= 24'b000000000000100110110010;
            7'h5b 	:	o_tw <= 24'b000000000000101001000110;
            7'h5c 	:	o_tw <= 24'b000000000000101011100011;
            7'h5d 	:	o_tw <= 24'b000000000000101110001000;
            7'h5e 	:	o_tw <= 24'b000000000000110000111000;
            7'h5f 	:	o_tw <= 24'b000000000000110011110010;
            7'h60 	:	o_tw <= 24'b000000000000110110110111;
            7'h61 	:	o_tw <= 24'b000000000000111010001000;
            7'h62 	:	o_tw <= 24'b000000000000111101100101;
            7'h63 	:	o_tw <= 24'b000000000001000001001111;
            7'h64 	:	o_tw <= 24'b000000000001000101001000;
            7'h65 	:	o_tw <= 24'b000000000001001001001111;
            7'h66 	:	o_tw <= 24'b000000000001001101100101;
            7'h67 	:	o_tw <= 24'b000000000001010010001101;
            7'h68 	:	o_tw <= 24'b000000000001010111000110;
            7'h69 	:	o_tw <= 24'b000000000001011100010001;
            7'h6a 	:	o_tw <= 24'b000000000001100001110000;
            7'h6b 	:	o_tw <= 24'b000000000001100111100100;
            7'h6c 	:	o_tw <= 24'b000000000001101101101110;
            7'h6d 	:	o_tw <= 24'b000000000001110100010000;
            7'h6e 	:	o_tw <= 24'b000000000001111011001011;
            7'h6f 	:	o_tw <= 24'b000000000010000010011111;
            7'h70 	:	o_tw <= 24'b000000000010001010010000;
            7'h71 	:	o_tw <= 24'b000000000010010010011110;
            7'h72 	:	o_tw <= 24'b000000000010011011001011;
            7'h73 	:	o_tw <= 24'b000000000010100100011010;
            7'h74 	:	o_tw <= 24'b000000000010101110001100;
            7'h75 	:	o_tw <= 24'b000000000010111000100011;
            7'h76 	:	o_tw <= 24'b000000000011000011100001;
            7'h77 	:	o_tw <= 24'b000000000011001111001001;
            7'h78 	:	o_tw <= 24'b000000000011011011011101;
            7'h79 	:	o_tw <= 24'b000000000011101000100001;
            7'h7a 	:	o_tw <= 24'b000000000011110110010110;
            7'h7b 	:	o_tw <= 24'b000000000100000100111111;
            7'h7c 	:	o_tw <= 24'b000000000100010100100000;
            7'h7d 	:	o_tw <= 24'b000000000100100100111101;
            7'h7e 	:	o_tw <= 24'b000000000100110110010111;
            7'h7f 	:	o_tw <= 24'b000000000101001000110101;
				default 	:	o_tw <= 24'h0000; // h00 is MIDI 0 value
			endcase
		end	
endmodule
